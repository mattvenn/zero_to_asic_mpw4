magic
tech sky130A
magscale 1 2
timestamp 1640263499
<< metal1 >>
rect 75822 703604 75828 703656
rect 75880 703644 75886 703656
rect 202598 703644 202604 703656
rect 75880 703616 202604 703644
rect 75880 703604 75886 703616
rect 202598 703604 202604 703616
rect 202656 703604 202662 703656
rect 86770 703536 86776 703588
rect 86828 703576 86834 703588
rect 234982 703576 234988 703588
rect 86828 703548 234988 703576
rect 86828 703536 86834 703548
rect 234982 703536 234988 703548
rect 235040 703536 235046 703588
rect 67634 703468 67640 703520
rect 67692 703508 67698 703520
rect 267458 703508 267464 703520
rect 67692 703480 267464 703508
rect 67692 703468 67698 703480
rect 267458 703468 267464 703480
rect 267516 703468 267522 703520
rect 93762 703400 93768 703452
rect 93820 703440 93826 703452
rect 300118 703440 300124 703452
rect 93820 703412 300124 703440
rect 93820 703400 93826 703412
rect 300118 703400 300124 703412
rect 300176 703400 300182 703452
rect 59262 703332 59268 703384
rect 59320 703372 59326 703384
rect 283834 703372 283840 703384
rect 59320 703344 283840 703372
rect 59320 703332 59326 703344
rect 283834 703332 283840 703344
rect 283892 703332 283898 703384
rect 73062 703264 73068 703316
rect 73120 703304 73126 703316
rect 332502 703304 332508 703316
rect 73120 703276 332508 703304
rect 73120 703264 73126 703276
rect 332502 703264 332508 703276
rect 332560 703264 332566 703316
rect 130378 703196 130384 703248
rect 130436 703236 130442 703248
rect 413646 703236 413652 703248
rect 130436 703208 413652 703236
rect 130436 703196 130442 703208
rect 413646 703196 413652 703208
rect 413704 703196 413710 703248
rect 61838 703128 61844 703180
rect 61896 703168 61902 703180
rect 348786 703168 348792 703180
rect 61896 703140 348792 703168
rect 61896 703128 61902 703140
rect 348786 703128 348792 703140
rect 348844 703128 348850 703180
rect 101398 703060 101404 703112
rect 101456 703100 101462 703112
rect 397454 703100 397460 703112
rect 101456 703072 397460 703100
rect 101456 703060 101462 703072
rect 397454 703060 397460 703072
rect 397512 703060 397518 703112
rect 124858 702992 124864 703044
rect 124916 703032 124922 703044
rect 429838 703032 429844 703044
rect 124916 703004 429844 703032
rect 124916 702992 124922 703004
rect 429838 702992 429844 703004
rect 429896 702992 429902 703044
rect 57698 702924 57704 702976
rect 57756 702964 57762 702976
rect 364978 702964 364984 702976
rect 57756 702936 364984 702964
rect 57756 702924 57762 702936
rect 364978 702924 364984 702936
rect 365036 702924 365042 702976
rect 126238 702856 126244 702908
rect 126296 702896 126302 702908
rect 462314 702896 462320 702908
rect 126296 702868 462320 702896
rect 126296 702856 126302 702868
rect 462314 702856 462320 702868
rect 462372 702856 462378 702908
rect 71038 702788 71044 702840
rect 71096 702828 71102 702840
rect 494790 702828 494796 702840
rect 71096 702800 494796 702828
rect 71096 702788 71102 702800
rect 494790 702788 494796 702800
rect 494848 702788 494854 702840
rect 97902 702720 97908 702772
rect 97960 702760 97966 702772
rect 478506 702760 478512 702772
rect 97960 702732 478512 702760
rect 97960 702720 97966 702732
rect 478506 702720 478512 702732
rect 478564 702720 478570 702772
rect 128998 702652 129004 702704
rect 129056 702692 129062 702704
rect 543458 702692 543464 702704
rect 129056 702664 543464 702692
rect 129056 702652 129062 702664
rect 543458 702652 543464 702664
rect 543516 702652 543522 702704
rect 8110 702584 8116 702636
rect 8168 702624 8174 702636
rect 89806 702624 89812 702636
rect 8168 702596 89812 702624
rect 8168 702584 8174 702596
rect 89806 702584 89812 702596
rect 89864 702584 89870 702636
rect 94498 702584 94504 702636
rect 94556 702624 94562 702636
rect 527174 702624 527180 702636
rect 94556 702596 527180 702624
rect 94556 702584 94562 702596
rect 527174 702584 527180 702596
rect 527232 702584 527238 702636
rect 53742 702516 53748 702568
rect 53800 702556 53806 702568
rect 580258 702556 580264 702568
rect 53800 702528 580264 702556
rect 53800 702516 53806 702528
rect 580258 702516 580264 702528
rect 580316 702516 580322 702568
rect 66162 702448 66168 702500
rect 66220 702488 66226 702500
rect 559650 702488 559656 702500
rect 66220 702460 559656 702488
rect 66220 702448 66226 702460
rect 559650 702448 559656 702460
rect 559708 702448 559714 702500
rect 84102 700272 84108 700324
rect 84160 700312 84166 700324
rect 89162 700312 89168 700324
rect 84160 700284 89168 700312
rect 84160 700272 84166 700284
rect 89162 700272 89168 700284
rect 89220 700272 89226 700324
rect 105446 700312 105452 700324
rect 93826 700284 105452 700312
rect 88978 700204 88984 700256
rect 89036 700244 89042 700256
rect 93826 700244 93854 700284
rect 105446 700272 105452 700284
rect 105504 700272 105510 700324
rect 133138 700272 133144 700324
rect 133196 700312 133202 700324
rect 218974 700312 218980 700324
rect 133196 700284 218980 700312
rect 133196 700272 133202 700284
rect 218974 700272 218980 700284
rect 219032 700272 219038 700324
rect 89036 700216 93854 700244
rect 89036 700204 89042 700216
rect 24302 698912 24308 698964
rect 24360 698952 24366 698964
rect 79318 698952 79324 698964
rect 24360 698924 79324 698952
rect 24360 698912 24366 698924
rect 79318 698912 79324 698924
rect 79376 698912 79382 698964
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 18598 683176 18604 683188
rect 3476 683148 18604 683176
rect 3476 683136 3482 683148
rect 18598 683136 18604 683148
rect 18656 683136 18662 683188
rect 3510 656888 3516 656940
rect 3568 656928 3574 656940
rect 22738 656928 22744 656940
rect 3568 656900 22744 656928
rect 3568 656888 3574 656900
rect 22738 656888 22744 656900
rect 22796 656888 22802 656940
rect 3418 639548 3424 639600
rect 3476 639588 3482 639600
rect 39298 639588 39304 639600
rect 3476 639560 39304 639588
rect 3476 639548 3482 639560
rect 39298 639548 39304 639560
rect 39356 639548 39362 639600
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 11698 632108 11704 632120
rect 3476 632080 11704 632108
rect 3476 632068 3482 632080
rect 11698 632068 11704 632080
rect 11756 632068 11762 632120
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 15838 618304 15844 618316
rect 3200 618276 15844 618304
rect 3200 618264 3206 618276
rect 15838 618264 15844 618276
rect 15896 618264 15902 618316
rect 3234 600924 3240 600976
rect 3292 600964 3298 600976
rect 88794 600964 88800 600976
rect 3292 600936 88800 600964
rect 3292 600924 3298 600936
rect 88794 600924 88800 600936
rect 88852 600924 88858 600976
rect 67450 599564 67456 599616
rect 67508 599604 67514 599616
rect 88978 599604 88984 599616
rect 67508 599576 88984 599604
rect 67508 599564 67514 599576
rect 88978 599564 88984 599576
rect 89036 599564 89042 599616
rect 79318 598884 79324 598936
rect 79376 598924 79382 598936
rect 80054 598924 80060 598936
rect 79376 598896 80060 598924
rect 79376 598884 79382 598896
rect 80054 598884 80060 598896
rect 80112 598884 80118 598936
rect 40034 598204 40040 598256
rect 40092 598244 40098 598256
rect 91094 598244 91100 598256
rect 40092 598216 91100 598244
rect 40092 598204 40098 598216
rect 91094 598204 91100 598216
rect 91152 598204 91158 598256
rect 80054 597524 80060 597576
rect 80112 597564 80118 597576
rect 106918 597564 106924 597576
rect 80112 597536 106924 597564
rect 80112 597524 80118 597536
rect 106918 597524 106924 597536
rect 106976 597524 106982 597576
rect 67542 596776 67548 596828
rect 67600 596816 67606 596828
rect 169754 596816 169760 596828
rect 67600 596788 169760 596816
rect 67600 596776 67606 596788
rect 169754 596776 169760 596788
rect 169812 596776 169818 596828
rect 72418 595416 72424 595468
rect 72476 595456 72482 595468
rect 84102 595456 84108 595468
rect 72476 595428 84108 595456
rect 72476 595416 72482 595428
rect 84102 595416 84108 595428
rect 84160 595456 84166 595468
rect 92474 595456 92480 595468
rect 84160 595428 92480 595456
rect 84160 595416 84166 595428
rect 92474 595416 92480 595428
rect 92532 595416 92538 595468
rect 74166 594804 74172 594856
rect 74224 594844 74230 594856
rect 95878 594844 95884 594856
rect 74224 594816 95884 594844
rect 74224 594804 74230 594816
rect 95878 594804 95884 594816
rect 95936 594804 95942 594856
rect 83458 593444 83464 593496
rect 83516 593484 83522 593496
rect 110414 593484 110420 593496
rect 83516 593456 110420 593484
rect 83516 593444 83522 593456
rect 110414 593444 110420 593456
rect 110472 593444 110478 593496
rect 90358 593376 90364 593428
rect 90416 593416 90422 593428
rect 582742 593416 582748 593428
rect 90416 593388 582748 593416
rect 90416 593376 90422 593388
rect 582742 593376 582748 593388
rect 582800 593376 582806 593428
rect 22738 592628 22744 592680
rect 22796 592668 22802 592680
rect 69014 592668 69020 592680
rect 22796 592640 69020 592668
rect 22796 592628 22802 592640
rect 69014 592628 69020 592640
rect 69072 592628 69078 592680
rect 75822 592084 75828 592136
rect 75880 592124 75886 592136
rect 96614 592124 96620 592136
rect 75880 592096 96620 592124
rect 75880 592084 75886 592096
rect 96614 592084 96620 592096
rect 96672 592084 96678 592136
rect 84102 592016 84108 592068
rect 84160 592056 84166 592068
rect 112438 592056 112444 592068
rect 84160 592028 112444 592056
rect 84160 592016 84166 592028
rect 112438 592016 112444 592028
rect 112496 592016 112502 592068
rect 78398 590792 78404 590844
rect 78456 590832 78462 590844
rect 89070 590832 89076 590844
rect 78456 590804 89076 590832
rect 78456 590792 78462 590804
rect 89070 590792 89076 590804
rect 89128 590792 89134 590844
rect 71682 590724 71688 590776
rect 71740 590764 71746 590776
rect 71740 590736 75040 590764
rect 71740 590724 71746 590736
rect 75012 590708 75040 590736
rect 86218 590724 86224 590776
rect 86276 590764 86282 590776
rect 90358 590764 90364 590776
rect 86276 590736 90364 590764
rect 86276 590724 86282 590736
rect 90358 590724 90364 590736
rect 90416 590724 90422 590776
rect 70302 590656 70308 590708
rect 70360 590696 70366 590708
rect 74442 590696 74448 590708
rect 70360 590668 74448 590696
rect 70360 590656 70366 590668
rect 74442 590656 74448 590668
rect 74500 590656 74506 590708
rect 74994 590656 75000 590708
rect 75052 590696 75058 590708
rect 75822 590696 75828 590708
rect 75052 590668 75828 590696
rect 75052 590656 75058 590668
rect 75822 590656 75828 590668
rect 75880 590656 75886 590708
rect 88794 590656 88800 590708
rect 88852 590696 88858 590708
rect 132494 590696 132500 590708
rect 88852 590668 132500 590696
rect 88852 590656 88858 590668
rect 132494 590656 132500 590668
rect 132552 590656 132558 590708
rect 3418 589976 3424 590028
rect 3476 590016 3482 590028
rect 71682 590016 71688 590028
rect 3476 589988 71688 590016
rect 3476 589976 3482 589988
rect 71682 589976 71688 589988
rect 71740 589976 71746 590028
rect 74442 589976 74448 590028
rect 74500 590016 74506 590028
rect 89714 590016 89720 590028
rect 74500 589988 89720 590016
rect 74500 589976 74506 589988
rect 89714 589976 89720 589988
rect 89772 589976 89778 590028
rect 67726 589908 67732 589960
rect 67784 589948 67790 589960
rect 580166 589948 580172 589960
rect 67784 589920 580172 589948
rect 67784 589908 67790 589920
rect 580166 589908 580172 589920
rect 580224 589908 580230 589960
rect 81434 589228 81440 589280
rect 81492 589268 81498 589280
rect 88242 589268 88248 589280
rect 81492 589240 88248 589268
rect 81492 589228 81498 589240
rect 88242 589228 88248 589240
rect 88300 589228 88306 589280
rect 69474 588616 69480 588668
rect 69532 588656 69538 588668
rect 88978 588656 88984 588668
rect 69532 588628 88984 588656
rect 69532 588616 69538 588628
rect 88978 588616 88984 588628
rect 89036 588616 89042 588668
rect 85298 588548 85304 588600
rect 85356 588588 85362 588600
rect 86954 588588 86960 588600
rect 85356 588560 86960 588588
rect 85356 588548 85362 588560
rect 86954 588548 86960 588560
rect 87012 588588 87018 588600
rect 113174 588588 113180 588600
rect 87012 588560 113180 588588
rect 87012 588548 87018 588560
rect 113174 588548 113180 588560
rect 113232 588548 113238 588600
rect 79778 588412 79784 588464
rect 79836 588412 79842 588464
rect 63310 587868 63316 587920
rect 63368 587908 63374 587920
rect 66806 587908 66812 587920
rect 63368 587880 66812 587908
rect 63368 587868 63374 587880
rect 66806 587868 66812 587880
rect 66864 587868 66870 587920
rect 79796 587160 79824 588412
rect 105538 587160 105544 587172
rect 79796 587132 105544 587160
rect 105538 587120 105544 587132
rect 105596 587120 105602 587172
rect 59170 586508 59176 586560
rect 59228 586548 59234 586560
rect 66254 586548 66260 586560
rect 59228 586520 66260 586548
rect 59228 586508 59234 586520
rect 66254 586508 66260 586520
rect 66312 586508 66318 586560
rect 91186 586508 91192 586560
rect 91244 586548 91250 586560
rect 141418 586548 141424 586560
rect 91244 586520 141424 586548
rect 91244 586508 91250 586520
rect 141418 586508 141424 586520
rect 141476 586508 141482 586560
rect 89070 585760 89076 585812
rect 89128 585800 89134 585812
rect 103514 585800 103520 585812
rect 89128 585772 103520 585800
rect 89128 585760 89134 585772
rect 103514 585760 103520 585772
rect 103572 585760 103578 585812
rect 50982 585148 50988 585200
rect 51040 585188 51046 585200
rect 67726 585188 67732 585200
rect 51040 585160 67732 585188
rect 51040 585148 51046 585160
rect 67726 585148 67732 585160
rect 67784 585148 67790 585200
rect 92106 584400 92112 584452
rect 92164 584440 92170 584452
rect 93762 584440 93768 584452
rect 92164 584412 93768 584440
rect 92164 584400 92170 584412
rect 93762 584400 93768 584412
rect 93820 584440 93826 584452
rect 115198 584440 115204 584452
rect 93820 584412 115204 584440
rect 93820 584400 93826 584412
rect 115198 584400 115204 584412
rect 115256 584400 115262 584452
rect 91922 583652 91928 583704
rect 91980 583692 91986 583704
rect 93762 583692 93768 583704
rect 91980 583664 93768 583692
rect 91980 583652 91986 583664
rect 93762 583652 93768 583664
rect 93820 583692 93826 583704
rect 94498 583692 94504 583704
rect 93820 583664 94504 583692
rect 93820 583652 93826 583664
rect 94498 583652 94504 583664
rect 94556 583652 94562 583704
rect 48130 582360 48136 582412
rect 48188 582400 48194 582412
rect 66806 582400 66812 582412
rect 48188 582372 66812 582400
rect 48188 582360 48194 582372
rect 66806 582360 66812 582372
rect 66864 582360 66870 582412
rect 64690 581000 64696 581052
rect 64748 581040 64754 581052
rect 66990 581040 66996 581052
rect 64748 581012 66996 581040
rect 64748 581000 64754 581012
rect 66990 581000 66996 581012
rect 67048 581000 67054 581052
rect 91186 581000 91192 581052
rect 91244 581040 91250 581052
rect 102778 581040 102784 581052
rect 91244 581012 102784 581040
rect 91244 581000 91250 581012
rect 102778 581000 102784 581012
rect 102836 581000 102842 581052
rect 91186 578212 91192 578264
rect 91244 578252 91250 578264
rect 121546 578252 121552 578264
rect 91244 578224 121552 578252
rect 91244 578212 91250 578224
rect 121546 578212 121552 578224
rect 121604 578212 121610 578264
rect 104802 577464 104808 577516
rect 104860 577504 104866 577516
rect 582466 577504 582472 577516
rect 104860 577476 582472 577504
rect 104860 577464 104866 577476
rect 582466 577464 582472 577476
rect 582524 577464 582530 577516
rect 91186 576852 91192 576904
rect 91244 576892 91250 576904
rect 104802 576892 104808 576904
rect 91244 576864 104808 576892
rect 91244 576852 91250 576864
rect 104802 576852 104808 576864
rect 104860 576852 104866 576904
rect 11698 576104 11704 576156
rect 11756 576144 11762 576156
rect 51074 576144 51080 576156
rect 11756 576116 51080 576144
rect 11756 576104 11762 576116
rect 51074 576104 51080 576116
rect 51132 576104 51138 576156
rect 51074 575492 51080 575544
rect 51132 575532 51138 575544
rect 52270 575532 52276 575544
rect 51132 575504 52276 575532
rect 51132 575492 51138 575504
rect 52270 575492 52276 575504
rect 52328 575532 52334 575544
rect 66898 575532 66904 575544
rect 52328 575504 66904 575532
rect 52328 575492 52334 575504
rect 66898 575492 66904 575504
rect 66956 575492 66962 575544
rect 88886 575492 88892 575544
rect 88944 575532 88950 575544
rect 105630 575532 105636 575544
rect 88944 575504 105636 575532
rect 88944 575492 88950 575504
rect 105630 575492 105636 575504
rect 105688 575492 105694 575544
rect 55030 574744 55036 574796
rect 55088 574784 55094 574796
rect 67450 574784 67456 574796
rect 55088 574756 67456 574784
rect 55088 574744 55094 574756
rect 67450 574744 67456 574756
rect 67508 574744 67514 574796
rect 91922 574744 91928 574796
rect 91980 574784 91986 574796
rect 93762 574784 93768 574796
rect 91980 574756 93768 574784
rect 91980 574744 91986 574756
rect 93762 574744 93768 574756
rect 93820 574784 93826 574796
rect 101398 574784 101404 574796
rect 93820 574756 101404 574784
rect 93820 574744 93826 574756
rect 101398 574744 101404 574756
rect 101456 574744 101462 574796
rect 41322 572704 41328 572756
rect 41380 572744 41386 572756
rect 66438 572744 66444 572756
rect 41380 572716 66444 572744
rect 41380 572704 41386 572716
rect 66438 572704 66444 572716
rect 66496 572704 66502 572756
rect 91094 572704 91100 572756
rect 91152 572744 91158 572756
rect 120810 572744 120816 572756
rect 91152 572716 120816 572744
rect 91152 572704 91158 572716
rect 120810 572704 120816 572716
rect 120868 572704 120874 572756
rect 91094 571412 91100 571464
rect 91152 571452 91158 571464
rect 97258 571452 97264 571464
rect 91152 571424 97264 571452
rect 91152 571412 91158 571424
rect 97258 571412 97264 571424
rect 97316 571412 97322 571464
rect 49602 571344 49608 571396
rect 49660 571384 49666 571396
rect 66438 571384 66444 571396
rect 49660 571356 66444 571384
rect 49660 571344 49666 571356
rect 66438 571344 66444 571356
rect 66496 571344 66502 571396
rect 91186 571344 91192 571396
rect 91244 571384 91250 571396
rect 126974 571384 126980 571396
rect 91244 571356 126980 571384
rect 91244 571344 91250 571356
rect 126974 571344 126980 571356
rect 127032 571344 127038 571396
rect 91094 569916 91100 569968
rect 91152 569956 91158 569968
rect 125594 569956 125600 569968
rect 91152 569928 125600 569956
rect 91152 569916 91158 569928
rect 125594 569916 125600 569928
rect 125652 569916 125658 569968
rect 93762 569168 93768 569220
rect 93820 569208 93826 569220
rect 123386 569208 123392 569220
rect 93820 569180 123392 569208
rect 93820 569168 93826 569180
rect 123386 569168 123392 569180
rect 123444 569168 123450 569220
rect 64782 568556 64788 568608
rect 64840 568596 64846 568608
rect 66806 568596 66812 568608
rect 64840 568568 66812 568596
rect 64840 568556 64846 568568
rect 66806 568556 66812 568568
rect 66864 568556 66870 568608
rect 91094 567808 91100 567860
rect 91152 567848 91158 567860
rect 91278 567848 91284 567860
rect 91152 567820 91284 567848
rect 91152 567808 91158 567820
rect 91278 567808 91284 567820
rect 91336 567848 91342 567860
rect 128354 567848 128360 567860
rect 91336 567820 128360 567848
rect 91336 567808 91342 567820
rect 128354 567808 128360 567820
rect 128412 567808 128418 567860
rect 57790 567196 57796 567248
rect 57848 567236 57854 567248
rect 66898 567236 66904 567248
rect 57848 567208 66904 567236
rect 57848 567196 57854 567208
rect 66898 567196 66904 567208
rect 66956 567196 66962 567248
rect 53650 566448 53656 566500
rect 53708 566488 53714 566500
rect 67542 566488 67548 566500
rect 53708 566460 67548 566488
rect 53708 566448 53714 566460
rect 67542 566448 67548 566460
rect 67600 566448 67606 566500
rect 91094 565836 91100 565888
rect 91152 565876 91158 565888
rect 101398 565876 101404 565888
rect 91152 565848 101404 565876
rect 91152 565836 91158 565848
rect 101398 565836 101404 565848
rect 101456 565836 101462 565888
rect 59998 564408 60004 564460
rect 60056 564448 60062 564460
rect 66622 564448 66628 564460
rect 60056 564420 66628 564448
rect 60056 564408 60062 564420
rect 66622 564408 66628 564420
rect 66680 564408 66686 564460
rect 91094 564408 91100 564460
rect 91152 564448 91158 564460
rect 120626 564448 120632 564460
rect 91152 564420 120632 564448
rect 91152 564408 91158 564420
rect 120626 564408 120632 564420
rect 120684 564408 120690 564460
rect 50890 564340 50896 564392
rect 50948 564380 50954 564392
rect 53742 564380 53748 564392
rect 50948 564352 53748 564380
rect 50948 564340 50954 564352
rect 53742 564340 53748 564352
rect 53800 564380 53806 564392
rect 66438 564380 66444 564392
rect 53800 564352 66444 564380
rect 53800 564340 53806 564352
rect 66438 564340 66444 564352
rect 66496 564340 66502 564392
rect 91094 563048 91100 563100
rect 91152 563088 91158 563100
rect 133874 563088 133880 563100
rect 91152 563060 133880 563088
rect 91152 563048 91158 563060
rect 133874 563048 133880 563060
rect 133932 563048 133938 563100
rect 45462 561688 45468 561740
rect 45520 561728 45526 561740
rect 66438 561728 66444 561740
rect 45520 561700 66444 561728
rect 45520 561688 45526 561700
rect 66438 561688 66444 561700
rect 66496 561688 66502 561740
rect 43990 560260 43996 560312
rect 44048 560300 44054 560312
rect 66622 560300 66628 560312
rect 44048 560272 66628 560300
rect 44048 560260 44054 560272
rect 66622 560260 66628 560272
rect 66680 560260 66686 560312
rect 56502 558900 56508 558952
rect 56560 558940 56566 558952
rect 66622 558940 66628 558952
rect 56560 558912 66628 558940
rect 56560 558900 56566 558912
rect 66622 558900 66628 558912
rect 66680 558900 66686 558952
rect 48222 557540 48228 557592
rect 48280 557580 48286 557592
rect 67634 557580 67640 557592
rect 48280 557552 67640 557580
rect 48280 557540 48286 557552
rect 67634 557540 67640 557552
rect 67692 557540 67698 557592
rect 91186 557540 91192 557592
rect 91244 557580 91250 557592
rect 124214 557580 124220 557592
rect 91244 557552 124220 557580
rect 91244 557540 91250 557552
rect 124214 557540 124220 557552
rect 124272 557540 124278 557592
rect 91186 556180 91192 556232
rect 91244 556220 91250 556232
rect 122098 556220 122104 556232
rect 91244 556192 122104 556220
rect 91244 556180 91250 556192
rect 122098 556180 122104 556192
rect 122156 556180 122162 556232
rect 58894 554752 58900 554804
rect 58952 554792 58958 554804
rect 66346 554792 66352 554804
rect 58952 554764 66352 554792
rect 58952 554752 58958 554764
rect 66346 554752 66352 554764
rect 66404 554752 66410 554804
rect 91186 554752 91192 554804
rect 91244 554792 91250 554804
rect 108942 554792 108948 554804
rect 91244 554764 108948 554792
rect 91244 554752 91250 554764
rect 108942 554752 108948 554764
rect 109000 554792 109006 554804
rect 582466 554792 582472 554804
rect 109000 554764 582472 554792
rect 109000 554752 109006 554764
rect 582466 554752 582472 554764
rect 582524 554752 582530 554804
rect 59262 554684 59268 554736
rect 59320 554724 59326 554736
rect 65518 554724 65524 554736
rect 59320 554696 65524 554724
rect 59320 554684 59326 554696
rect 65518 554684 65524 554696
rect 65576 554724 65582 554736
rect 66254 554724 66260 554736
rect 65576 554696 66260 554724
rect 65576 554684 65582 554696
rect 66254 554684 66260 554696
rect 66312 554684 66318 554736
rect 2774 553800 2780 553852
rect 2832 553840 2838 553852
rect 4798 553840 4804 553852
rect 2832 553812 4804 553840
rect 2832 553800 2838 553812
rect 4798 553800 4804 553812
rect 4856 553800 4862 553852
rect 107102 553052 107108 553104
rect 107160 553092 107166 553104
rect 109034 553092 109040 553104
rect 107160 553064 109040 553092
rect 107160 553052 107166 553064
rect 109034 553052 109040 553064
rect 109092 553052 109098 553104
rect 91186 552100 91192 552152
rect 91244 552140 91250 552152
rect 107010 552140 107016 552152
rect 91244 552112 107016 552140
rect 91244 552100 91250 552112
rect 107010 552100 107016 552112
rect 107068 552100 107074 552152
rect 91278 552032 91284 552084
rect 91336 552072 91342 552084
rect 130470 552072 130476 552084
rect 91336 552044 130476 552072
rect 91336 552032 91342 552044
rect 130470 552032 130476 552044
rect 130528 552032 130534 552084
rect 100018 551284 100024 551336
rect 100076 551324 100082 551336
rect 117314 551324 117320 551336
rect 100076 551296 117320 551324
rect 100076 551284 100082 551296
rect 117314 551284 117320 551296
rect 117372 551284 117378 551336
rect 63402 549244 63408 549296
rect 63460 549284 63466 549296
rect 66530 549284 66536 549296
rect 63460 549256 66536 549284
rect 63460 549244 63466 549256
rect 66530 549244 66536 549256
rect 66588 549244 66594 549296
rect 91186 549244 91192 549296
rect 91244 549284 91250 549296
rect 111058 549284 111064 549296
rect 91244 549256 111064 549284
rect 91244 549244 91250 549256
rect 111058 549244 111064 549256
rect 111116 549244 111122 549296
rect 91830 548496 91836 548548
rect 91888 548536 91894 548548
rect 121454 548536 121460 548548
rect 91888 548508 121460 548536
rect 91888 548496 91894 548508
rect 121454 548496 121460 548508
rect 121512 548496 121518 548548
rect 62022 547884 62028 547936
rect 62080 547924 62086 547936
rect 66530 547924 66536 547936
rect 62080 547896 66536 547924
rect 62080 547884 62086 547896
rect 66530 547884 66536 547896
rect 66588 547884 66594 547936
rect 61838 547748 61844 547800
rect 61896 547788 61902 547800
rect 66806 547788 66812 547800
rect 61896 547760 66812 547788
rect 61896 547748 61902 547760
rect 66806 547748 66812 547760
rect 66864 547748 66870 547800
rect 53742 547136 53748 547188
rect 53800 547176 53806 547188
rect 61838 547176 61844 547188
rect 53800 547148 61844 547176
rect 53800 547136 53806 547148
rect 61838 547136 61844 547148
rect 61896 547136 61902 547188
rect 91278 546456 91284 546508
rect 91336 546496 91342 546508
rect 104158 546496 104164 546508
rect 91336 546468 104164 546496
rect 91336 546456 91342 546468
rect 104158 546456 104164 546468
rect 104216 546456 104222 546508
rect 57882 545708 57888 545760
rect 57940 545748 57946 545760
rect 66162 545748 66168 545760
rect 57940 545720 66168 545748
rect 57940 545708 57946 545720
rect 66162 545708 66168 545720
rect 66220 545708 66226 545760
rect 108114 545708 108120 545760
rect 108172 545748 108178 545760
rect 126238 545748 126244 545760
rect 108172 545720 126244 545748
rect 108172 545708 108178 545720
rect 126238 545708 126244 545720
rect 126296 545708 126302 545760
rect 52362 545028 52368 545080
rect 52420 545068 52426 545080
rect 57698 545068 57704 545080
rect 52420 545040 57704 545068
rect 52420 545028 52426 545040
rect 57698 545028 57704 545040
rect 57756 545068 57762 545080
rect 66806 545068 66812 545080
rect 57756 545040 66812 545068
rect 57756 545028 57762 545040
rect 66806 545028 66812 545040
rect 66864 545028 66870 545080
rect 91278 544348 91284 544400
rect 91336 544388 91342 544400
rect 96522 544388 96528 544400
rect 91336 544360 96528 544388
rect 91336 544348 91342 544360
rect 96522 544348 96528 544360
rect 96580 544388 96586 544400
rect 128998 544388 129004 544400
rect 96580 544360 129004 544388
rect 96580 544348 96586 544360
rect 128998 544348 129004 544360
rect 129056 544348 129062 544400
rect 18598 542988 18604 543040
rect 18656 543028 18662 543040
rect 39942 543028 39948 543040
rect 18656 543000 39948 543028
rect 18656 542988 18662 543000
rect 39942 542988 39948 543000
rect 40000 542988 40006 543040
rect 39942 542376 39948 542428
rect 40000 542416 40006 542428
rect 66806 542416 66812 542428
rect 40000 542388 66812 542416
rect 40000 542376 40006 542388
rect 66806 542376 66812 542388
rect 66864 542376 66870 542428
rect 91278 542376 91284 542428
rect 91336 542416 91342 542428
rect 94498 542416 94504 542428
rect 91336 542388 94504 542416
rect 91336 542376 91342 542388
rect 94498 542376 94504 542388
rect 94556 542376 94562 542428
rect 39298 541628 39304 541680
rect 39356 541668 39362 541680
rect 67082 541668 67088 541680
rect 39356 541640 67088 541668
rect 39356 541628 39362 541640
rect 67082 541628 67088 541640
rect 67140 541628 67146 541680
rect 91278 541628 91284 541680
rect 91336 541668 91342 541680
rect 136634 541668 136640 541680
rect 91336 541640 136640 541668
rect 91336 541628 91342 541640
rect 136634 541628 136640 541640
rect 136692 541628 136698 541680
rect 67542 540880 67548 540932
rect 67600 540920 67606 540932
rect 68646 540920 68652 540932
rect 67600 540892 68652 540920
rect 67600 540880 67606 540892
rect 68646 540880 68652 540892
rect 68704 540920 68710 540932
rect 582650 540920 582656 540932
rect 68704 540892 582656 540920
rect 68704 540880 68710 540892
rect 582650 540880 582656 540892
rect 582708 540880 582714 540932
rect 3418 540200 3424 540252
rect 3476 540240 3482 540252
rect 3476 540212 64874 540240
rect 3476 540200 3482 540212
rect 64846 539696 64874 540212
rect 64846 539668 69888 539696
rect 69860 539640 69888 539668
rect 91278 539656 91284 539708
rect 91336 539696 91342 539708
rect 93118 539696 93124 539708
rect 91336 539668 93124 539696
rect 91336 539656 91342 539668
rect 93118 539656 93124 539668
rect 93176 539656 93182 539708
rect 55122 539588 55128 539640
rect 55180 539628 55186 539640
rect 67542 539628 67548 539640
rect 55180 539600 67548 539628
rect 55180 539588 55186 539600
rect 67542 539588 67548 539600
rect 67600 539588 67606 539640
rect 69842 539588 69848 539640
rect 69900 539588 69906 539640
rect 115382 539520 115388 539572
rect 115440 539560 115446 539572
rect 582558 539560 582564 539572
rect 115440 539532 582564 539560
rect 115440 539520 115446 539532
rect 582558 539520 582564 539532
rect 582616 539520 582622 539572
rect 67082 539452 67088 539504
rect 67140 539492 67146 539504
rect 67542 539492 67548 539504
rect 67140 539464 67548 539492
rect 67140 539452 67146 539464
rect 67542 539452 67548 539464
rect 67600 539452 67606 539504
rect 67818 538976 67824 539028
rect 67876 539016 67882 539028
rect 74626 539016 74632 539028
rect 67876 538988 74632 539016
rect 67876 538976 67882 538988
rect 74626 538976 74632 538988
rect 74684 538976 74690 539028
rect 3418 538840 3424 538892
rect 3476 538880 3482 538892
rect 89898 538880 89904 538892
rect 3476 538852 89904 538880
rect 3476 538840 3482 538852
rect 89898 538840 89904 538852
rect 89956 538840 89962 538892
rect 81066 538228 81072 538280
rect 81124 538268 81130 538280
rect 115382 538268 115388 538280
rect 81124 538240 115388 538268
rect 81124 538228 81130 538240
rect 115382 538228 115388 538240
rect 115440 538228 115446 538280
rect 4798 538160 4804 538212
rect 4856 538200 4862 538212
rect 70670 538200 70676 538212
rect 4856 538172 70676 538200
rect 4856 538160 4862 538172
rect 70670 538160 70676 538172
rect 70728 538160 70734 538212
rect 86862 538160 86868 538212
rect 86920 538200 86926 538212
rect 133138 538200 133144 538212
rect 86920 538172 133144 538200
rect 86920 538160 86926 538172
rect 133138 538160 133144 538172
rect 133196 538160 133202 538212
rect 72418 537480 72424 537532
rect 72476 537520 72482 537532
rect 579798 537520 579804 537532
rect 72476 537492 579804 537520
rect 72476 537480 72482 537492
rect 579798 537480 579804 537492
rect 579856 537480 579862 537532
rect 82722 536732 82728 536784
rect 82780 536772 82786 536784
rect 130378 536772 130384 536784
rect 82780 536744 130384 536772
rect 82780 536732 82786 536744
rect 130378 536732 130384 536744
rect 130436 536732 130442 536784
rect 85482 536188 85488 536240
rect 85540 536228 85546 536240
rect 86218 536228 86224 536240
rect 85540 536200 86224 536228
rect 85540 536188 85546 536200
rect 86218 536188 86224 536200
rect 86276 536188 86282 536240
rect 66162 536120 66168 536172
rect 66220 536160 66226 536172
rect 76190 536160 76196 536172
rect 66220 536132 76196 536160
rect 66220 536120 66226 536132
rect 76190 536120 76196 536132
rect 76248 536120 76254 536172
rect 15838 536052 15844 536104
rect 15896 536092 15902 536104
rect 44082 536092 44088 536104
rect 15896 536064 44088 536092
rect 15896 536052 15902 536064
rect 44082 536052 44088 536064
rect 44140 536092 44146 536104
rect 73154 536092 73160 536104
rect 44140 536064 73160 536092
rect 44140 536052 44146 536064
rect 73154 536052 73160 536064
rect 73212 536052 73218 536104
rect 73154 535440 73160 535492
rect 73212 535480 73218 535492
rect 73982 535480 73988 535492
rect 73212 535452 73988 535480
rect 73212 535440 73218 535452
rect 73982 535440 73988 535452
rect 74040 535440 74046 535492
rect 78766 535440 78772 535492
rect 78824 535480 78830 535492
rect 79502 535480 79508 535492
rect 78824 535452 79508 535480
rect 78824 535440 78830 535452
rect 79502 535440 79508 535452
rect 79560 535440 79566 535492
rect 7558 534692 7564 534744
rect 7616 534732 7622 534744
rect 91370 534732 91376 534744
rect 7616 534704 91376 534732
rect 7616 534692 7622 534704
rect 91370 534692 91376 534704
rect 91428 534692 91434 534744
rect 56502 534012 56508 534064
rect 56560 534052 56566 534064
rect 580258 534052 580264 534064
rect 56560 534024 580264 534052
rect 56560 534012 56566 534024
rect 580258 534012 580264 534024
rect 580316 534012 580322 534064
rect 5442 533332 5448 533384
rect 5500 533372 5506 533384
rect 91186 533372 91192 533384
rect 5500 533344 91192 533372
rect 5500 533332 5506 533344
rect 91186 533332 91192 533344
rect 91244 533332 91250 533384
rect 66070 531972 66076 532024
rect 66128 532012 66134 532024
rect 77938 532012 77944 532024
rect 66128 531984 77944 532012
rect 66128 531972 66134 531984
rect 77938 531972 77944 531984
rect 77996 531972 78002 532024
rect 15838 530544 15844 530596
rect 15896 530584 15902 530596
rect 91094 530584 91100 530596
rect 15896 530556 91100 530584
rect 15896 530544 15902 530556
rect 91094 530544 91100 530556
rect 91152 530544 91158 530596
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 14458 514808 14464 514820
rect 3568 514780 14464 514808
rect 3568 514768 3574 514780
rect 14458 514768 14464 514780
rect 14516 514768 14522 514820
rect 43990 511232 43996 511284
rect 44048 511272 44054 511284
rect 580166 511272 580172 511284
rect 44048 511244 580172 511272
rect 44048 511232 44054 511244
rect 580166 511232 580172 511244
rect 580224 511232 580230 511284
rect 3326 502052 3332 502104
rect 3384 502092 3390 502104
rect 7558 502092 7564 502104
rect 3384 502064 7564 502092
rect 3384 502052 3390 502064
rect 7558 502052 7564 502064
rect 7616 502052 7622 502104
rect 4062 475328 4068 475380
rect 4120 475368 4126 475380
rect 5442 475368 5448 475380
rect 4120 475340 5448 475368
rect 4120 475328 4126 475340
rect 5442 475328 5448 475340
rect 5500 475368 5506 475380
rect 11698 475368 11704 475380
rect 5500 475340 11704 475368
rect 5500 475328 5506 475340
rect 11698 475328 11704 475340
rect 11756 475328 11762 475380
rect 67726 467780 67732 467832
rect 67784 467820 67790 467832
rect 76558 467820 76564 467832
rect 67784 467792 76564 467820
rect 67784 467780 67790 467792
rect 76558 467780 76564 467792
rect 76616 467780 76622 467832
rect 63310 465060 63316 465112
rect 63368 465100 63374 465112
rect 87046 465100 87052 465112
rect 63368 465072 87052 465100
rect 63368 465060 63374 465072
rect 87046 465060 87052 465072
rect 87104 465060 87110 465112
rect 56410 464312 56416 464364
rect 56468 464352 56474 464364
rect 78766 464352 78772 464364
rect 56468 464324 78772 464352
rect 56468 464312 56474 464324
rect 78766 464312 78772 464324
rect 78824 464312 78830 464364
rect 2774 462544 2780 462596
rect 2832 462584 2838 462596
rect 4798 462584 4804 462596
rect 2832 462556 4804 462584
rect 2832 462544 2838 462556
rect 4798 462544 4804 462556
rect 4856 462544 4862 462596
rect 59170 461592 59176 461644
rect 59228 461632 59234 461644
rect 85574 461632 85580 461644
rect 59228 461604 85580 461632
rect 59228 461592 59234 461604
rect 85574 461592 85580 461604
rect 85632 461592 85638 461644
rect 64690 460164 64696 460216
rect 64748 460204 64754 460216
rect 78674 460204 78680 460216
rect 64748 460176 78680 460204
rect 64748 460164 64754 460176
rect 78674 460164 78680 460176
rect 78732 460164 78738 460216
rect 64690 458872 64696 458924
rect 64748 458912 64754 458924
rect 70486 458912 70492 458924
rect 64748 458884 70492 458912
rect 64748 458872 64754 458884
rect 70486 458872 70492 458884
rect 70544 458872 70550 458924
rect 53466 458804 53472 458856
rect 53524 458844 53530 458856
rect 77294 458844 77300 458856
rect 53524 458816 77300 458844
rect 53524 458804 53530 458816
rect 77294 458804 77300 458816
rect 77352 458804 77358 458856
rect 102778 458804 102784 458856
rect 102836 458844 102842 458856
rect 123110 458844 123116 458856
rect 102836 458816 123116 458844
rect 102836 458804 102842 458816
rect 123110 458804 123116 458816
rect 123168 458804 123174 458856
rect 50982 457444 50988 457496
rect 51040 457484 51046 457496
rect 83458 457484 83464 457496
rect 51040 457456 83464 457484
rect 51040 457444 51046 457456
rect 83458 457444 83464 457456
rect 83516 457444 83522 457496
rect 105630 457444 105636 457496
rect 105688 457484 105694 457496
rect 122926 457484 122932 457496
rect 105688 457456 122932 457484
rect 105688 457444 105694 457456
rect 122926 457444 122932 457456
rect 122984 457444 122990 457496
rect 60550 456084 60556 456136
rect 60608 456124 60614 456136
rect 76098 456124 76104 456136
rect 60608 456096 76104 456124
rect 60608 456084 60614 456096
rect 76098 456084 76104 456096
rect 76156 456084 76162 456136
rect 101398 456084 101404 456136
rect 101456 456124 101462 456136
rect 123570 456124 123576 456136
rect 101456 456096 123576 456124
rect 101456 456084 101462 456096
rect 123570 456084 123576 456096
rect 123628 456084 123634 456136
rect 61930 456016 61936 456068
rect 61988 456056 61994 456068
rect 91094 456056 91100 456068
rect 61988 456028 91100 456056
rect 61988 456016 61994 456028
rect 91094 456016 91100 456028
rect 91152 456016 91158 456068
rect 97258 456016 97264 456068
rect 97316 456056 97322 456068
rect 124398 456056 124404 456068
rect 97316 456028 124404 456056
rect 97316 456016 97322 456028
rect 124398 456016 124404 456028
rect 124456 456016 124462 456068
rect 59078 454724 59084 454776
rect 59136 454764 59142 454776
rect 73154 454764 73160 454776
rect 59136 454736 73160 454764
rect 59136 454724 59142 454736
rect 73154 454724 73160 454736
rect 73212 454724 73218 454776
rect 55030 454656 55036 454708
rect 55088 454696 55094 454708
rect 72050 454696 72056 454708
rect 55088 454668 72056 454696
rect 55088 454656 55094 454668
rect 72050 454656 72056 454668
rect 72108 454656 72114 454708
rect 91094 454044 91100 454096
rect 91152 454084 91158 454096
rect 161474 454084 161480 454096
rect 91152 454056 161480 454084
rect 91152 454044 91158 454056
rect 161474 454044 161480 454056
rect 161532 454044 161538 454096
rect 49602 453296 49608 453348
rect 49660 453336 49666 453348
rect 67634 453336 67640 453348
rect 49660 453308 67640 453336
rect 49660 453296 49666 453308
rect 67634 453296 67640 453308
rect 67692 453296 67698 453348
rect 72050 452684 72056 452736
rect 72108 452724 72114 452736
rect 126330 452724 126336 452736
rect 72108 452696 126336 452724
rect 72108 452684 72114 452696
rect 126330 452684 126336 452696
rect 126388 452684 126394 452736
rect 112438 452616 112444 452668
rect 112496 452656 112502 452668
rect 179414 452656 179420 452668
rect 112496 452628 179420 452656
rect 112496 452616 112502 452628
rect 179414 452616 179420 452628
rect 179472 452616 179478 452668
rect 61930 451936 61936 451988
rect 61988 451976 61994 451988
rect 78858 451976 78864 451988
rect 61988 451948 78864 451976
rect 61988 451936 61994 451948
rect 78858 451936 78864 451948
rect 78916 451936 78922 451988
rect 3418 451868 3424 451920
rect 3476 451908 3482 451920
rect 120718 451908 120724 451920
rect 3476 451880 120724 451908
rect 3476 451868 3482 451880
rect 120718 451868 120724 451880
rect 120776 451868 120782 451920
rect 14458 451188 14464 451240
rect 14516 451228 14522 451240
rect 112438 451228 112444 451240
rect 14516 451200 112444 451228
rect 14516 451188 14522 451200
rect 112438 451188 112444 451200
rect 112496 451188 112502 451240
rect 116578 449964 116584 450016
rect 116636 450004 116642 450016
rect 160094 450004 160100 450016
rect 116636 449976 160100 450004
rect 116636 449964 116642 449976
rect 160094 449964 160100 449976
rect 160152 449964 160158 450016
rect 49510 449896 49516 449948
rect 49568 449936 49574 449948
rect 74626 449936 74632 449948
rect 49568 449908 74632 449936
rect 49568 449896 49574 449908
rect 74626 449896 74632 449908
rect 74684 449896 74690 449948
rect 95878 449896 95884 449948
rect 95936 449936 95942 449948
rect 178034 449936 178040 449948
rect 95936 449908 178040 449936
rect 95936 449896 95942 449908
rect 178034 449896 178040 449908
rect 178092 449896 178098 449948
rect 41322 449828 41328 449880
rect 41380 449868 41386 449880
rect 69658 449868 69664 449880
rect 41380 449840 69664 449868
rect 41380 449828 41386 449840
rect 69658 449828 69664 449840
rect 69716 449828 69722 449880
rect 48130 449148 48136 449200
rect 48188 449188 48194 449200
rect 80054 449188 80060 449200
rect 48188 449160 80060 449188
rect 48188 449148 48194 449160
rect 80054 449148 80060 449160
rect 80112 449148 80118 449200
rect 173802 449148 173808 449200
rect 173860 449188 173866 449200
rect 582466 449188 582472 449200
rect 173860 449160 582472 449188
rect 173860 449148 173866 449160
rect 582466 449148 582472 449160
rect 582524 449148 582530 449200
rect 77938 448604 77944 448656
rect 77996 448644 78002 448656
rect 124306 448644 124312 448656
rect 77996 448616 124312 448644
rect 77996 448604 78002 448616
rect 124306 448604 124312 448616
rect 124364 448604 124370 448656
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 14458 448576 14464 448588
rect 3200 448548 14464 448576
rect 3200 448536 3206 448548
rect 14458 448536 14464 448548
rect 14516 448536 14522 448588
rect 80054 448536 80060 448588
rect 80112 448576 80118 448588
rect 80882 448576 80888 448588
rect 80112 448548 80888 448576
rect 80112 448536 80118 448548
rect 80882 448536 80888 448548
rect 80940 448576 80946 448588
rect 173802 448576 173808 448588
rect 80940 448548 173808 448576
rect 80940 448536 80946 448548
rect 173802 448536 173808 448548
rect 173860 448536 173866 448588
rect 52270 447856 52276 447908
rect 52328 447896 52334 447908
rect 73338 447896 73344 447908
rect 52328 447868 73344 447896
rect 52328 447856 52334 447868
rect 73338 447856 73344 447868
rect 73396 447856 73402 447908
rect 4798 447788 4804 447840
rect 4856 447828 4862 447840
rect 68278 447828 68284 447840
rect 4856 447800 68284 447828
rect 4856 447788 4862 447800
rect 68278 447788 68284 447800
rect 68336 447788 68342 447840
rect 115198 447788 115204 447840
rect 115256 447828 115262 447840
rect 125686 447828 125692 447840
rect 115256 447800 125692 447828
rect 115256 447788 115262 447800
rect 125686 447788 125692 447800
rect 125744 447788 125750 447840
rect 68278 447176 68284 447228
rect 68336 447216 68342 447228
rect 68554 447216 68560 447228
rect 68336 447188 68560 447216
rect 68336 447176 68342 447188
rect 68554 447176 68560 447188
rect 68612 447216 68618 447228
rect 103514 447216 103520 447228
rect 68612 447188 103520 447216
rect 68612 447176 68618 447188
rect 103514 447176 103520 447188
rect 103572 447176 103578 447228
rect 98638 447108 98644 447160
rect 98696 447148 98702 447160
rect 170398 447148 170404 447160
rect 98696 447120 170404 447148
rect 98696 447108 98702 447120
rect 170398 447108 170404 447120
rect 170456 447108 170462 447160
rect 78674 446904 78680 446956
rect 78732 446944 78738 446956
rect 79134 446944 79140 446956
rect 78732 446916 79140 446944
rect 78732 446904 78738 446916
rect 79134 446904 79140 446916
rect 79192 446904 79198 446956
rect 64506 446360 64512 446412
rect 64564 446400 64570 446412
rect 74534 446400 74540 446412
rect 64564 446372 74540 446400
rect 64564 446360 64570 446372
rect 74534 446360 74540 446372
rect 74592 446360 74598 446412
rect 106918 445816 106924 445868
rect 106976 445856 106982 445868
rect 124858 445856 124864 445868
rect 106976 445828 124864 445856
rect 106976 445816 106982 445828
rect 124858 445816 124864 445828
rect 124916 445816 124922 445868
rect 50982 445748 50988 445800
rect 51040 445788 51046 445800
rect 79134 445788 79140 445800
rect 51040 445760 79140 445788
rect 51040 445748 51046 445760
rect 79134 445748 79140 445760
rect 79192 445748 79198 445800
rect 97994 445748 98000 445800
rect 98052 445788 98058 445800
rect 102134 445788 102140 445800
rect 98052 445760 102140 445788
rect 98052 445748 98058 445760
rect 102134 445748 102140 445760
rect 102192 445748 102198 445800
rect 105538 445748 105544 445800
rect 105596 445788 105602 445800
rect 201494 445788 201500 445800
rect 105596 445760 201500 445788
rect 105596 445748 105602 445760
rect 201494 445748 201500 445760
rect 201552 445748 201558 445800
rect 66070 445000 66076 445052
rect 66128 445040 66134 445052
rect 72418 445040 72424 445052
rect 66128 445012 72424 445040
rect 66128 445000 66134 445012
rect 72418 445000 72424 445012
rect 72476 445000 72482 445052
rect 67634 444592 67640 444644
rect 67692 444632 67698 444644
rect 67818 444632 67824 444644
rect 67692 444604 67824 444632
rect 67692 444592 67698 444604
rect 67818 444592 67824 444604
rect 67876 444632 67882 444644
rect 68784 444632 68790 444644
rect 67876 444604 68790 444632
rect 67876 444592 67882 444604
rect 68784 444592 68790 444604
rect 68842 444592 68848 444644
rect 73338 444456 73344 444508
rect 73396 444496 73402 444508
rect 144178 444496 144184 444508
rect 73396 444468 144184 444496
rect 73396 444456 73402 444468
rect 144178 444456 144184 444468
rect 144236 444456 144242 444508
rect 4798 444388 4804 444440
rect 4856 444428 4862 444440
rect 119154 444428 119160 444440
rect 4856 444400 119160 444428
rect 4856 444388 4862 444400
rect 119154 444388 119160 444400
rect 119212 444428 119218 444440
rect 120902 444428 120908 444440
rect 119212 444400 120908 444428
rect 119212 444388 119218 444400
rect 120902 444388 120908 444400
rect 120960 444388 120966 444440
rect 124122 444320 124128 444372
rect 124180 444360 124186 444372
rect 132494 444360 132500 444372
rect 124180 444332 132500 444360
rect 124180 444320 124186 444332
rect 132494 444320 132500 444332
rect 132552 444360 132558 444372
rect 133782 444360 133788 444372
rect 132552 444332 133788 444360
rect 132552 444320 132558 444332
rect 133782 444320 133788 444332
rect 133840 444320 133846 444372
rect 133782 443640 133788 443692
rect 133840 443680 133846 443692
rect 166258 443680 166264 443692
rect 133840 443652 166264 443680
rect 133840 443640 133846 443652
rect 166258 443640 166264 443652
rect 166316 443640 166322 443692
rect 67266 442892 67272 442944
rect 67324 442932 67330 442944
rect 67726 442932 67732 442944
rect 67324 442904 67732 442932
rect 67324 442892 67330 442904
rect 67726 442892 67732 442904
rect 67784 442892 67790 442944
rect 124122 441600 124128 441652
rect 124180 441640 124186 441652
rect 133138 441640 133144 441652
rect 124180 441612 133144 441640
rect 124180 441600 124186 441612
rect 133138 441600 133144 441612
rect 133196 441600 133202 441652
rect 64782 439084 64788 439136
rect 64840 439124 64846 439136
rect 66990 439124 66996 439136
rect 64840 439096 66996 439124
rect 64840 439084 64846 439096
rect 66990 439084 66996 439096
rect 67048 439124 67054 439136
rect 67266 439124 67272 439136
rect 67048 439096 67272 439124
rect 67048 439084 67054 439096
rect 67266 439084 67272 439096
rect 67324 439084 67330 439136
rect 121178 438880 121184 438932
rect 121236 438920 121242 438932
rect 169754 438920 169760 438932
rect 121236 438892 169760 438920
rect 121236 438880 121242 438892
rect 169754 438880 169760 438892
rect 169812 438880 169818 438932
rect 123846 438132 123852 438184
rect 123904 438172 123910 438184
rect 125686 438172 125692 438184
rect 123904 438144 125692 438172
rect 123904 438132 123910 438144
rect 125686 438132 125692 438144
rect 125744 438172 125750 438184
rect 157978 438172 157984 438184
rect 125744 438144 157984 438172
rect 125744 438132 125750 438144
rect 157978 438132 157984 438144
rect 158036 438132 158042 438184
rect 57790 437452 57796 437504
rect 57848 437492 57854 437504
rect 60642 437492 60648 437504
rect 57848 437464 60648 437492
rect 57848 437452 57854 437464
rect 60642 437452 60648 437464
rect 60700 437492 60706 437504
rect 66806 437492 66812 437504
rect 60700 437464 66812 437492
rect 60700 437452 60706 437464
rect 66806 437452 66812 437464
rect 66864 437452 66870 437504
rect 53650 436024 53656 436076
rect 53708 436064 53714 436076
rect 57698 436064 57704 436076
rect 53708 436036 57704 436064
rect 53708 436024 53714 436036
rect 57698 436024 57704 436036
rect 57756 436024 57762 436076
rect 57698 434732 57704 434784
rect 57756 434772 57762 434784
rect 66806 434772 66812 434784
rect 57756 434744 66812 434772
rect 57756 434732 57762 434744
rect 66806 434732 66812 434744
rect 66864 434732 66870 434784
rect 58986 433848 58992 433900
rect 59044 433888 59050 433900
rect 59998 433888 60004 433900
rect 59044 433860 60004 433888
rect 59044 433848 59050 433860
rect 59998 433848 60004 433860
rect 60056 433848 60062 433900
rect 124122 432556 124128 432608
rect 124180 432596 124186 432608
rect 135162 432596 135168 432608
rect 124180 432568 135168 432596
rect 124180 432556 124186 432568
rect 135162 432556 135168 432568
rect 135220 432596 135226 432608
rect 582374 432596 582380 432608
rect 135220 432568 582380 432596
rect 135220 432556 135226 432568
rect 582374 432556 582380 432568
rect 582432 432556 582438 432608
rect 58986 432012 58992 432064
rect 59044 432052 59050 432064
rect 66898 432052 66904 432064
rect 59044 432024 66904 432052
rect 59044 432012 59050 432024
rect 66898 432012 66904 432024
rect 66956 432012 66962 432064
rect 50890 431876 50896 431928
rect 50948 431916 50954 431928
rect 66898 431916 66904 431928
rect 50948 431888 66904 431916
rect 50948 431876 50954 431888
rect 66898 431876 66904 431888
rect 66956 431876 66962 431928
rect 48130 430584 48136 430636
rect 48188 430624 48194 430636
rect 50890 430624 50896 430636
rect 48188 430596 50896 430624
rect 48188 430584 48194 430596
rect 50890 430584 50896 430596
rect 50948 430584 50954 430636
rect 40678 429088 40684 429140
rect 40736 429128 40742 429140
rect 45462 429128 45468 429140
rect 40736 429100 45468 429128
rect 40736 429088 40742 429100
rect 45462 429088 45468 429100
rect 45520 429128 45526 429140
rect 66806 429128 66812 429140
rect 45520 429100 66812 429128
rect 45520 429088 45526 429100
rect 66806 429088 66812 429100
rect 66864 429088 66870 429140
rect 61838 426368 61844 426420
rect 61896 426408 61902 426420
rect 66254 426408 66260 426420
rect 61896 426380 66260 426408
rect 61896 426368 61902 426380
rect 66254 426368 66260 426380
rect 66312 426368 66318 426420
rect 56502 425008 56508 425060
rect 56560 425048 56566 425060
rect 66254 425048 66260 425060
rect 56560 425020 66260 425048
rect 56560 425008 56566 425020
rect 66254 425008 66260 425020
rect 66312 425008 66318 425060
rect 3142 422900 3148 422952
rect 3200 422940 3206 422952
rect 15838 422940 15844 422952
rect 3200 422912 15844 422940
rect 3200 422900 3206 422912
rect 15838 422900 15844 422912
rect 15896 422900 15902 422952
rect 48222 421540 48228 421592
rect 48280 421580 48286 421592
rect 61838 421580 61844 421592
rect 48280 421552 61844 421580
rect 48280 421540 48286 421552
rect 61838 421540 61844 421552
rect 61896 421580 61902 421592
rect 66254 421580 66260 421592
rect 61896 421552 66260 421580
rect 61896 421540 61902 421552
rect 66254 421540 66260 421552
rect 66312 421540 66318 421592
rect 123386 421540 123392 421592
rect 123444 421580 123450 421592
rect 148318 421580 148324 421592
rect 123444 421552 148324 421580
rect 123444 421540 123450 421552
rect 148318 421540 148324 421552
rect 148376 421540 148382 421592
rect 121546 418072 121552 418124
rect 121604 418112 121610 418124
rect 126974 418112 126980 418124
rect 121604 418084 126980 418112
rect 121604 418072 121610 418084
rect 126974 418072 126980 418084
rect 127032 418072 127038 418124
rect 58894 416780 58900 416832
rect 58952 416820 58958 416832
rect 63310 416820 63316 416832
rect 58952 416792 63316 416820
rect 58952 416780 58958 416792
rect 63310 416780 63316 416792
rect 63368 416820 63374 416832
rect 66898 416820 66904 416832
rect 63368 416792 66904 416820
rect 63368 416780 63374 416792
rect 66898 416780 66904 416792
rect 66956 416780 66962 416832
rect 65518 415148 65524 415200
rect 65576 415188 65582 415200
rect 66438 415188 66444 415200
rect 65576 415160 66444 415188
rect 65576 415148 65582 415160
rect 66438 415148 66444 415160
rect 66496 415148 66502 415200
rect 123110 415080 123116 415132
rect 123168 415120 123174 415132
rect 124398 415120 124404 415132
rect 123168 415092 124404 415120
rect 123168 415080 123174 415092
rect 124398 415080 124404 415092
rect 124456 415120 124462 415132
rect 126974 415120 126980 415132
rect 124456 415092 126980 415120
rect 124456 415080 124462 415092
rect 126974 415080 126980 415092
rect 127032 415080 127038 415132
rect 57790 414672 57796 414724
rect 57848 414712 57854 414724
rect 65518 414712 65524 414724
rect 57848 414684 65524 414712
rect 57848 414672 57854 414684
rect 65518 414672 65524 414684
rect 65576 414672 65582 414724
rect 123110 413924 123116 413976
rect 123168 413964 123174 413976
rect 125594 413964 125600 413976
rect 123168 413936 125600 413964
rect 123168 413924 123174 413936
rect 125594 413924 125600 413936
rect 125652 413924 125658 413976
rect 121638 409844 121644 409896
rect 121696 409884 121702 409896
rect 162854 409884 162860 409896
rect 121696 409856 162860 409884
rect 121696 409844 121702 409856
rect 162854 409844 162860 409856
rect 162912 409844 162918 409896
rect 63402 408416 63408 408468
rect 63460 408456 63466 408468
rect 65978 408456 65984 408468
rect 63460 408428 65984 408456
rect 63460 408416 63466 408428
rect 65978 408416 65984 408428
rect 66036 408456 66042 408468
rect 66530 408456 66536 408468
rect 66036 408428 66536 408456
rect 66036 408416 66042 408428
rect 66530 408416 66536 408428
rect 66588 408416 66594 408468
rect 124122 408348 124128 408400
rect 124180 408388 124186 408400
rect 128354 408388 128360 408400
rect 124180 408360 128360 408388
rect 124180 408348 124186 408360
rect 128354 408348 128360 408360
rect 128412 408348 128418 408400
rect 128354 407736 128360 407788
rect 128412 407776 128418 407788
rect 135898 407776 135904 407788
rect 128412 407748 135904 407776
rect 128412 407736 128418 407748
rect 135898 407736 135904 407748
rect 135956 407736 135962 407788
rect 122098 407056 122104 407108
rect 122156 407096 122162 407108
rect 123018 407096 123024 407108
rect 122156 407068 123024 407096
rect 122156 407056 122162 407068
rect 123018 407056 123024 407068
rect 123076 407056 123082 407108
rect 123570 405832 123576 405884
rect 123628 405872 123634 405884
rect 124858 405872 124864 405884
rect 123628 405844 124864 405872
rect 123628 405832 123634 405844
rect 124858 405832 124864 405844
rect 124916 405832 124922 405884
rect 62022 405764 62028 405816
rect 62080 405804 62086 405816
rect 64598 405804 64604 405816
rect 62080 405776 64604 405804
rect 62080 405764 62086 405776
rect 64598 405764 64604 405776
rect 64656 405804 64662 405816
rect 66622 405804 66628 405816
rect 64656 405776 66628 405804
rect 64656 405764 64662 405776
rect 66622 405764 66628 405776
rect 66680 405764 66686 405816
rect 57606 404812 57612 404864
rect 57664 404852 57670 404864
rect 57882 404852 57888 404864
rect 57664 404824 57888 404852
rect 57664 404812 57670 404824
rect 57882 404812 57888 404824
rect 57940 404812 57946 404864
rect 57974 403588 57980 403640
rect 58032 403628 58038 403640
rect 66346 403628 66352 403640
rect 58032 403600 66352 403628
rect 58032 403588 58038 403600
rect 66346 403588 66352 403600
rect 66404 403588 66410 403640
rect 162762 403588 162768 403640
rect 162820 403628 162826 403640
rect 582374 403628 582380 403640
rect 162820 403600 582380 403628
rect 162820 403588 162826 403600
rect 582374 403588 582380 403600
rect 582432 403588 582438 403640
rect 120626 402976 120632 403028
rect 120684 403016 120690 403028
rect 161566 403016 161572 403028
rect 120684 402988 161572 403016
rect 120684 402976 120690 402988
rect 161566 402976 161572 402988
rect 161624 403016 161630 403028
rect 162762 403016 162768 403028
rect 161624 402988 162768 403016
rect 161624 402976 161630 402988
rect 162762 402976 162768 402988
rect 162820 402976 162826 403028
rect 53558 402228 53564 402280
rect 53616 402268 53622 402280
rect 57974 402268 57980 402280
rect 53616 402240 57980 402268
rect 53616 402228 53622 402240
rect 57974 402228 57980 402240
rect 58032 402228 58038 402280
rect 50890 401548 50896 401600
rect 50948 401588 50954 401600
rect 57606 401588 57612 401600
rect 50948 401560 57612 401588
rect 50948 401548 50954 401560
rect 57606 401548 57612 401560
rect 57664 401588 57670 401600
rect 66806 401588 66812 401600
rect 57664 401560 66812 401588
rect 57664 401548 57670 401560
rect 66806 401548 66812 401560
rect 66864 401548 66870 401600
rect 124122 401548 124128 401600
rect 124180 401588 124186 401600
rect 133874 401588 133880 401600
rect 124180 401560 133880 401588
rect 124180 401548 124186 401560
rect 133874 401548 133880 401560
rect 133932 401588 133938 401600
rect 135070 401588 135076 401600
rect 133932 401560 135076 401588
rect 133932 401548 133938 401560
rect 135070 401548 135076 401560
rect 135128 401548 135134 401600
rect 135070 400868 135076 400920
rect 135128 400908 135134 400920
rect 158070 400908 158076 400920
rect 135128 400880 158076 400908
rect 135128 400868 135134 400880
rect 158070 400868 158076 400880
rect 158128 400868 158134 400920
rect 52362 398828 52368 398880
rect 52420 398868 52426 398880
rect 53650 398868 53656 398880
rect 52420 398840 53656 398868
rect 52420 398828 52426 398840
rect 53650 398828 53656 398840
rect 53708 398868 53714 398880
rect 66898 398868 66904 398880
rect 53708 398840 66904 398868
rect 53708 398828 53714 398840
rect 66898 398828 66904 398840
rect 66956 398828 66962 398880
rect 123662 398828 123668 398880
rect 123720 398868 123726 398880
rect 124950 398868 124956 398880
rect 123720 398840 124956 398868
rect 123720 398828 123726 398840
rect 124950 398828 124956 398840
rect 125008 398828 125014 398880
rect 2774 398692 2780 398744
rect 2832 398732 2838 398744
rect 4798 398732 4804 398744
rect 2832 398704 4804 398732
rect 2832 398692 2838 398704
rect 4798 398692 4804 398704
rect 4856 398692 4862 398744
rect 39942 396720 39948 396772
rect 40000 396760 40006 396772
rect 66254 396760 66260 396772
rect 40000 396732 66260 396760
rect 40000 396720 40006 396732
rect 66254 396720 66260 396732
rect 66312 396720 66318 396772
rect 121454 396040 121460 396092
rect 121512 396080 121518 396092
rect 177390 396080 177396 396092
rect 121512 396052 177396 396080
rect 121512 396040 121518 396052
rect 177390 396040 177396 396052
rect 177448 396040 177454 396092
rect 55122 392572 55128 392624
rect 55180 392612 55186 392624
rect 65518 392612 65524 392624
rect 55180 392584 65524 392612
rect 55180 392572 55186 392584
rect 65518 392572 65524 392584
rect 65576 392572 65582 392624
rect 124950 391960 124956 392012
rect 125008 392000 125014 392012
rect 166350 392000 166356 392012
rect 125008 391972 166356 392000
rect 125008 391960 125014 391972
rect 166350 391960 166356 391972
rect 166408 391960 166414 392012
rect 15838 391348 15844 391400
rect 15896 391388 15902 391400
rect 124950 391388 124956 391400
rect 15896 391360 124956 391388
rect 15896 391348 15902 391360
rect 124950 391348 124956 391360
rect 125008 391348 125014 391400
rect 111702 389784 111708 389836
rect 111760 389824 111766 389836
rect 121546 389824 121552 389836
rect 111760 389796 121552 389824
rect 111760 389784 111766 389796
rect 121546 389784 121552 389796
rect 121604 389784 121610 389836
rect 59078 389240 59084 389292
rect 59136 389280 59142 389292
rect 77386 389280 77392 389292
rect 59136 389252 77392 389280
rect 59136 389240 59142 389252
rect 77386 389240 77392 389252
rect 77444 389240 77450 389292
rect 11698 389172 11704 389224
rect 11756 389212 11762 389224
rect 111610 389212 111616 389224
rect 11756 389184 111616 389212
rect 11756 389172 11762 389184
rect 111610 389172 111616 389184
rect 111668 389172 111674 389224
rect 130470 389212 130476 389224
rect 129752 389184 130476 389212
rect 64690 389104 64696 389156
rect 64748 389144 64754 389156
rect 73154 389144 73160 389156
rect 64748 389116 73160 389144
rect 64748 389104 64754 389116
rect 73154 389104 73160 389116
rect 73212 389144 73218 389156
rect 73338 389144 73344 389156
rect 73212 389116 73344 389144
rect 73212 389104 73218 389116
rect 73338 389104 73344 389116
rect 73396 389104 73402 389156
rect 91922 389104 91928 389156
rect 91980 389144 91986 389156
rect 93210 389144 93216 389156
rect 91980 389116 93216 389144
rect 91980 389104 91986 389116
rect 93210 389104 93216 389116
rect 93268 389104 93274 389156
rect 102594 389104 102600 389156
rect 102652 389144 102658 389156
rect 105538 389144 105544 389156
rect 102652 389116 105544 389144
rect 102652 389104 102658 389116
rect 105538 389104 105544 389116
rect 105596 389104 105602 389156
rect 117866 389104 117872 389156
rect 117924 389144 117930 389156
rect 129752 389144 129780 389184
rect 130470 389172 130476 389184
rect 130528 389212 130534 389224
rect 168374 389212 168380 389224
rect 130528 389184 168380 389212
rect 130528 389172 130534 389184
rect 168374 389172 168380 389184
rect 168432 389172 168438 389224
rect 117924 389116 129780 389144
rect 117924 389104 117930 389116
rect 66070 389036 66076 389088
rect 66128 389076 66134 389088
rect 74534 389076 74540 389088
rect 66128 389048 74540 389076
rect 66128 389036 66134 389048
rect 74534 389036 74540 389048
rect 74592 389036 74598 389088
rect 111610 388628 111616 388680
rect 111668 388668 111674 388680
rect 112438 388668 112444 388680
rect 111668 388640 112444 388668
rect 111668 388628 111674 388640
rect 112438 388628 112444 388640
rect 112496 388628 112502 388680
rect 93394 388424 93400 388476
rect 93452 388464 93458 388476
rect 100110 388464 100116 388476
rect 93452 388436 100116 388464
rect 93452 388424 93458 388436
rect 100110 388424 100116 388436
rect 100168 388424 100174 388476
rect 101398 388424 101404 388476
rect 101456 388464 101462 388476
rect 120166 388464 120172 388476
rect 101456 388436 120172 388464
rect 101456 388424 101462 388436
rect 120166 388424 120172 388436
rect 120224 388424 120230 388476
rect 94682 387812 94688 387864
rect 94740 387812 94746 387864
rect 64506 387744 64512 387796
rect 64564 387784 64570 387796
rect 79134 387784 79140 387796
rect 64564 387756 79140 387784
rect 64564 387744 64570 387756
rect 79134 387744 79140 387756
rect 79192 387744 79198 387796
rect 93118 387744 93124 387796
rect 93176 387784 93182 387796
rect 94700 387784 94728 387812
rect 128446 387784 128452 387796
rect 93176 387756 128452 387784
rect 93176 387744 93182 387756
rect 128446 387744 128452 387756
rect 128504 387744 128510 387796
rect 78674 387268 78680 387320
rect 78732 387308 78738 387320
rect 79134 387308 79140 387320
rect 78732 387280 79140 387308
rect 78732 387268 78738 387280
rect 79134 387268 79140 387280
rect 79192 387268 79198 387320
rect 60550 386316 60556 386368
rect 60608 386356 60614 386368
rect 82078 386356 82084 386368
rect 60608 386328 82084 386356
rect 60608 386316 60614 386328
rect 82078 386316 82084 386328
rect 82136 386316 82142 386368
rect 110138 385636 110144 385688
rect 110196 385676 110202 385688
rect 155218 385676 155224 385688
rect 110196 385648 155224 385676
rect 110196 385636 110202 385648
rect 155218 385636 155224 385648
rect 155276 385636 155282 385688
rect 56410 384956 56416 385008
rect 56468 384996 56474 385008
rect 87046 384996 87052 385008
rect 56468 384968 87052 384996
rect 56468 384956 56474 384968
rect 87046 384956 87052 384968
rect 87104 384956 87110 385008
rect 104066 384956 104072 385008
rect 104124 384996 104130 385008
rect 136634 384996 136640 385008
rect 104124 384968 136640 384996
rect 104124 384956 104130 384968
rect 136634 384956 136640 384968
rect 136692 384996 136698 385008
rect 137094 384996 137100 385008
rect 136692 384968 137100 384996
rect 136692 384956 136698 384968
rect 137094 384956 137100 384968
rect 137152 384956 137158 385008
rect 87046 384344 87052 384396
rect 87104 384384 87110 384396
rect 88242 384384 88248 384396
rect 87104 384356 88248 384384
rect 87104 384344 87110 384356
rect 88242 384344 88248 384356
rect 88300 384344 88306 384396
rect 5442 384276 5448 384328
rect 5500 384316 5506 384328
rect 123110 384316 123116 384328
rect 5500 384288 123116 384316
rect 5500 384276 5506 384288
rect 123110 384276 123116 384288
rect 123168 384276 123174 384328
rect 137094 384276 137100 384328
rect 137152 384316 137158 384328
rect 169110 384316 169116 384328
rect 137152 384288 169116 384316
rect 137152 384276 137158 384288
rect 169110 384276 169116 384288
rect 169168 384276 169174 384328
rect 36538 382236 36544 382288
rect 36596 382276 36602 382288
rect 118694 382276 118700 382288
rect 36596 382248 118700 382276
rect 36596 382236 36602 382248
rect 118694 382236 118700 382248
rect 118752 382276 118758 382288
rect 119430 382276 119436 382288
rect 118752 382248 119436 382276
rect 118752 382236 118758 382248
rect 119430 382236 119436 382248
rect 119488 382236 119494 382288
rect 88334 382168 88340 382220
rect 88392 382208 88398 382220
rect 115106 382208 115112 382220
rect 88392 382180 115112 382208
rect 88392 382168 88398 382180
rect 115106 382168 115112 382180
rect 115164 382208 115170 382220
rect 115750 382208 115756 382220
rect 115164 382180 115756 382208
rect 115164 382168 115170 382180
rect 115750 382168 115756 382180
rect 115808 382168 115814 382220
rect 115750 380876 115756 380928
rect 115808 380916 115814 380928
rect 130470 380916 130476 380928
rect 115808 380888 130476 380916
rect 115808 380876 115814 380888
rect 130470 380876 130476 380888
rect 130528 380876 130534 380928
rect 67634 380196 67640 380248
rect 67692 380236 67698 380248
rect 123202 380236 123208 380248
rect 67692 380208 123208 380236
rect 67692 380196 67698 380208
rect 123202 380196 123208 380208
rect 123260 380196 123266 380248
rect 61746 380128 61752 380180
rect 61804 380168 61810 380180
rect 158714 380168 158720 380180
rect 61804 380140 158720 380168
rect 61804 380128 61810 380140
rect 158714 380128 158720 380140
rect 158772 380128 158778 380180
rect 44082 379448 44088 379500
rect 44140 379488 44146 379500
rect 75914 379488 75920 379500
rect 44140 379460 75920 379488
rect 44140 379448 44146 379460
rect 75914 379448 75920 379460
rect 75972 379488 75978 379500
rect 76558 379488 76564 379500
rect 75972 379460 76564 379488
rect 75972 379448 75978 379460
rect 76558 379448 76564 379460
rect 76616 379448 76622 379500
rect 63218 378768 63224 378820
rect 63276 378808 63282 378820
rect 87598 378808 87604 378820
rect 63276 378780 87604 378808
rect 63276 378768 63282 378780
rect 87598 378768 87604 378780
rect 87656 378768 87662 378820
rect 67818 375980 67824 376032
rect 67876 376020 67882 376032
rect 145558 376020 145564 376032
rect 67876 375992 145564 376020
rect 67876 375980 67882 375992
rect 145558 375980 145564 375992
rect 145616 375980 145622 376032
rect 67726 374620 67732 374672
rect 67784 374660 67790 374672
rect 124950 374660 124956 374672
rect 67784 374632 124956 374660
rect 67784 374620 67790 374632
rect 124950 374620 124956 374632
rect 125008 374620 125014 374672
rect 150250 374076 150256 374128
rect 150308 374116 150314 374128
rect 242158 374116 242164 374128
rect 150308 374088 242164 374116
rect 150308 374076 150314 374088
rect 242158 374076 242164 374088
rect 242216 374076 242222 374128
rect 57698 374008 57704 374060
rect 57756 374048 57762 374060
rect 193858 374048 193864 374060
rect 57756 374020 193864 374048
rect 57756 374008 57762 374020
rect 193858 374008 193864 374020
rect 193916 374008 193922 374060
rect 107470 373260 107476 373312
rect 107528 373300 107534 373312
rect 164234 373300 164240 373312
rect 107528 373272 164240 373300
rect 107528 373260 107534 373272
rect 164234 373260 164240 373272
rect 164292 373260 164298 373312
rect 150342 372580 150348 372632
rect 150400 372620 150406 372632
rect 248506 372620 248512 372632
rect 150400 372592 248512 372620
rect 150400 372580 150406 372592
rect 248506 372580 248512 372592
rect 248564 372580 248570 372632
rect 137278 372172 137284 372224
rect 137336 372212 137342 372224
rect 137922 372212 137928 372224
rect 137336 372184 137928 372212
rect 137336 372172 137342 372184
rect 137922 372172 137928 372184
rect 137980 372172 137986 372224
rect 70302 371832 70308 371884
rect 70360 371872 70366 371884
rect 155954 371872 155960 371884
rect 70360 371844 155960 371872
rect 70360 371832 70366 371844
rect 155954 371832 155960 371844
rect 156012 371832 156018 371884
rect 137922 371220 137928 371272
rect 137980 371260 137986 371272
rect 180794 371260 180800 371272
rect 137980 371232 180800 371260
rect 137980 371220 137986 371232
rect 180794 371220 180800 371232
rect 180852 371220 180858 371272
rect 133138 370540 133144 370592
rect 133196 370580 133202 370592
rect 164878 370580 164884 370592
rect 133196 370552 164884 370580
rect 133196 370540 133202 370552
rect 164878 370540 164884 370552
rect 164936 370540 164942 370592
rect 64598 370472 64604 370524
rect 64656 370512 64662 370524
rect 108298 370512 108304 370524
rect 64656 370484 108304 370512
rect 64656 370472 64662 370484
rect 108298 370472 108304 370484
rect 108356 370472 108362 370524
rect 108850 370472 108856 370524
rect 108908 370512 108914 370524
rect 160738 370512 160744 370524
rect 108908 370484 160744 370512
rect 108908 370472 108914 370484
rect 160738 370472 160744 370484
rect 160796 370472 160802 370524
rect 121454 368908 121460 368960
rect 121512 368948 121518 368960
rect 122098 368948 122104 368960
rect 121512 368920 122104 368948
rect 121512 368908 121518 368920
rect 122098 368908 122104 368920
rect 122156 368908 122162 368960
rect 85574 368568 85580 368620
rect 85632 368608 85638 368620
rect 215386 368608 215392 368620
rect 85632 368580 215392 368608
rect 85632 368568 85638 368580
rect 215386 368568 215392 368580
rect 215444 368568 215450 368620
rect 62022 368500 62028 368552
rect 62080 368540 62086 368552
rect 121454 368540 121460 368552
rect 62080 368512 121460 368540
rect 62080 368500 62086 368512
rect 121454 368500 121460 368512
rect 121512 368500 121518 368552
rect 144822 368500 144828 368552
rect 144880 368540 144886 368552
rect 306742 368540 306748 368552
rect 144880 368512 306748 368540
rect 144880 368500 144886 368512
rect 306742 368500 306748 368512
rect 306800 368500 306806 368552
rect 119430 367752 119436 367804
rect 119488 367792 119494 367804
rect 166994 367792 167000 367804
rect 119488 367764 167000 367792
rect 119488 367752 119494 367764
rect 166994 367752 167000 367764
rect 167052 367752 167058 367804
rect 126330 367072 126336 367124
rect 126388 367112 126394 367124
rect 209038 367112 209044 367124
rect 126388 367084 209044 367112
rect 126388 367072 126394 367084
rect 209038 367072 209044 367084
rect 209096 367072 209102 367124
rect 86954 366324 86960 366376
rect 87012 366364 87018 366376
rect 95234 366364 95240 366376
rect 87012 366336 95240 366364
rect 87012 366324 87018 366336
rect 95234 366324 95240 366336
rect 95292 366324 95298 366376
rect 99282 366324 99288 366376
rect 99340 366364 99346 366376
rect 173250 366364 173256 366376
rect 99340 366336 173256 366364
rect 99340 366324 99346 366336
rect 173250 366324 173256 366336
rect 173308 366324 173314 366376
rect 102778 365712 102784 365764
rect 102836 365752 102842 365764
rect 304994 365752 305000 365764
rect 102836 365724 305000 365752
rect 102836 365712 102842 365724
rect 304994 365712 305000 365724
rect 305052 365712 305058 365764
rect 81434 365644 81440 365696
rect 81492 365684 81498 365696
rect 82078 365684 82084 365696
rect 81492 365656 82084 365684
rect 81492 365644 81498 365656
rect 82078 365644 82084 365656
rect 82136 365644 82142 365696
rect 71682 365236 71688 365288
rect 71740 365276 71746 365288
rect 73154 365276 73160 365288
rect 71740 365248 73160 365276
rect 71740 365236 71746 365248
rect 73154 365236 73160 365248
rect 73212 365236 73218 365288
rect 136634 364420 136640 364472
rect 136692 364460 136698 364472
rect 204898 364460 204904 364472
rect 136692 364432 204904 364460
rect 136692 364420 136698 364432
rect 204898 364420 204904 364432
rect 204956 364420 204962 364472
rect 81434 364352 81440 364404
rect 81492 364392 81498 364404
rect 240502 364392 240508 364404
rect 81492 364364 240508 364392
rect 81492 364352 81498 364364
rect 240502 364352 240508 364364
rect 240560 364352 240566 364404
rect 122098 363604 122104 363656
rect 122156 363644 122162 363656
rect 208118 363644 208124 363656
rect 122156 363616 208124 363644
rect 122156 363604 122162 363616
rect 208118 363604 208124 363616
rect 208176 363604 208182 363656
rect 100018 362924 100024 362976
rect 100076 362964 100082 362976
rect 196618 362964 196624 362976
rect 100076 362936 196624 362964
rect 100076 362924 100082 362936
rect 196618 362924 196624 362936
rect 196676 362924 196682 362976
rect 147674 361632 147680 361684
rect 147732 361672 147738 361684
rect 155586 361672 155592 361684
rect 147732 361644 155592 361672
rect 147732 361632 147738 361644
rect 155586 361632 155592 361644
rect 155644 361632 155650 361684
rect 107562 361564 107568 361616
rect 107620 361604 107626 361616
rect 186958 361604 186964 361616
rect 107620 361576 186964 361604
rect 107620 361564 107626 361576
rect 186958 361564 186964 361576
rect 187016 361564 187022 361616
rect 124858 360272 124864 360324
rect 124916 360312 124922 360324
rect 125594 360312 125600 360324
rect 124916 360284 125600 360312
rect 124916 360272 124922 360284
rect 125594 360272 125600 360284
rect 125652 360272 125658 360324
rect 128354 360272 128360 360324
rect 128412 360312 128418 360324
rect 166442 360312 166448 360324
rect 128412 360284 166448 360312
rect 128412 360272 128418 360284
rect 166442 360272 166448 360284
rect 166500 360272 166506 360324
rect 120074 360204 120080 360256
rect 120132 360244 120138 360256
rect 214558 360244 214564 360256
rect 120132 360216 214564 360244
rect 120132 360204 120138 360216
rect 214558 360204 214564 360216
rect 214616 360204 214622 360256
rect 132494 358844 132500 358896
rect 132552 358884 132558 358896
rect 174722 358884 174728 358896
rect 132552 358856 174728 358884
rect 132552 358844 132558 358856
rect 174722 358844 174728 358856
rect 174780 358844 174786 358896
rect 88978 358776 88984 358828
rect 89036 358816 89042 358828
rect 91186 358816 91192 358828
rect 89036 358788 91192 358816
rect 89036 358776 89042 358788
rect 91186 358776 91192 358788
rect 91244 358816 91250 358828
rect 213178 358816 213184 358828
rect 91244 358788 213184 358816
rect 91244 358776 91250 358788
rect 213178 358776 213184 358788
rect 213236 358776 213242 358828
rect 3326 358708 3332 358760
rect 3384 358748 3390 358760
rect 36538 358748 36544 358760
rect 3384 358720 36544 358748
rect 3384 358708 3390 358720
rect 36538 358708 36544 358720
rect 36596 358708 36602 358760
rect 107838 358708 107844 358760
rect 107896 358748 107902 358760
rect 108298 358748 108304 358760
rect 107896 358720 108304 358748
rect 107896 358708 107902 358720
rect 108298 358708 108304 358720
rect 108356 358708 108362 358760
rect 135898 357484 135904 357536
rect 135956 357524 135962 357536
rect 192570 357524 192576 357536
rect 135956 357496 192576 357524
rect 135956 357484 135962 357496
rect 192570 357484 192576 357496
rect 192628 357484 192634 357536
rect 107838 357416 107844 357468
rect 107896 357456 107902 357468
rect 241514 357456 241520 357468
rect 107896 357428 241520 357456
rect 107896 357416 107902 357428
rect 241514 357416 241520 357428
rect 241572 357416 241578 357468
rect 92382 356668 92388 356720
rect 92440 356708 92446 356720
rect 121454 356708 121460 356720
rect 92440 356680 121460 356708
rect 92440 356668 92446 356680
rect 121454 356668 121460 356680
rect 121512 356668 121518 356720
rect 132402 356124 132408 356176
rect 132460 356164 132466 356176
rect 176102 356164 176108 356176
rect 132460 356136 176108 356164
rect 132460 356124 132466 356136
rect 176102 356124 176108 356136
rect 176160 356124 176166 356176
rect 122834 356056 122840 356108
rect 122892 356096 122898 356108
rect 225598 356096 225604 356108
rect 122892 356068 225604 356096
rect 122892 356056 122898 356068
rect 225598 356056 225604 356068
rect 225656 356056 225662 356108
rect 155586 355988 155592 356040
rect 155644 356028 155650 356040
rect 159358 356028 159364 356040
rect 155644 356000 159364 356028
rect 155644 355988 155650 356000
rect 159358 355988 159364 356000
rect 159416 355988 159422 356040
rect 52270 355308 52276 355360
rect 52328 355348 52334 355360
rect 93854 355348 93860 355360
rect 52328 355320 93860 355348
rect 52328 355308 52334 355320
rect 93854 355308 93860 355320
rect 93912 355348 93918 355360
rect 95142 355348 95148 355360
rect 93912 355320 95148 355348
rect 93912 355308 93918 355320
rect 95142 355308 95148 355320
rect 95200 355308 95206 355360
rect 97810 355308 97816 355360
rect 97868 355348 97874 355360
rect 154666 355348 154672 355360
rect 97868 355320 154672 355348
rect 97868 355308 97874 355320
rect 154666 355308 154672 355320
rect 154724 355308 154730 355360
rect 51718 355036 51724 355088
rect 51776 355076 51782 355088
rect 52270 355076 52276 355088
rect 51776 355048 52276 355076
rect 51776 355036 51782 355048
rect 52270 355036 52276 355048
rect 52328 355036 52334 355088
rect 123478 354696 123484 354748
rect 123536 354736 123542 354748
rect 184290 354736 184296 354748
rect 123536 354708 184296 354736
rect 123536 354696 123542 354708
rect 184290 354696 184296 354708
rect 184348 354696 184354 354748
rect 93210 353948 93216 354000
rect 93268 353988 93274 354000
rect 118786 353988 118792 354000
rect 93268 353960 118792 353988
rect 93268 353948 93274 353960
rect 118786 353948 118792 353960
rect 118844 353948 118850 354000
rect 122742 353948 122748 354000
rect 122800 353988 122806 354000
rect 126330 353988 126336 354000
rect 122800 353960 126336 353988
rect 122800 353948 122806 353960
rect 126330 353948 126336 353960
rect 126388 353948 126394 354000
rect 132586 353336 132592 353388
rect 132644 353376 132650 353388
rect 222930 353376 222936 353388
rect 132644 353348 222936 353376
rect 132644 353336 132650 353348
rect 222930 353336 222936 353348
rect 222988 353336 222994 353388
rect 61930 353268 61936 353320
rect 61988 353308 61994 353320
rect 218698 353308 218704 353320
rect 61988 353280 218704 353308
rect 61988 353268 61994 353280
rect 218698 353268 218704 353280
rect 218756 353268 218762 353320
rect 104802 352588 104808 352640
rect 104860 352628 104866 352640
rect 120718 352628 120724 352640
rect 104860 352600 120724 352628
rect 104860 352588 104866 352600
rect 120718 352588 120724 352600
rect 120776 352588 120782 352640
rect 83458 352520 83464 352572
rect 83516 352560 83522 352572
rect 101398 352560 101404 352572
rect 83516 352532 101404 352560
rect 83516 352520 83522 352532
rect 101398 352520 101404 352532
rect 101456 352520 101462 352572
rect 105630 352520 105636 352572
rect 105688 352560 105694 352572
rect 155310 352560 155316 352572
rect 105688 352532 155316 352560
rect 105688 352520 105694 352532
rect 155310 352520 155316 352532
rect 155368 352520 155374 352572
rect 144178 352248 144184 352300
rect 144236 352288 144242 352300
rect 144730 352288 144736 352300
rect 144236 352260 144736 352288
rect 144236 352248 144242 352260
rect 144730 352248 144736 352260
rect 144788 352248 144794 352300
rect 144730 351908 144736 351960
rect 144788 351948 144794 351960
rect 184382 351948 184388 351960
rect 144788 351920 184388 351948
rect 144788 351908 144794 351920
rect 184382 351908 184388 351920
rect 184440 351908 184446 351960
rect 79962 351228 79968 351280
rect 80020 351268 80026 351280
rect 111058 351268 111064 351280
rect 80020 351240 111064 351268
rect 80020 351228 80026 351240
rect 111058 351228 111064 351240
rect 111116 351228 111122 351280
rect 67818 351160 67824 351212
rect 67876 351200 67882 351212
rect 122834 351200 122840 351212
rect 67876 351172 122840 351200
rect 67876 351160 67882 351172
rect 122834 351160 122840 351172
rect 122892 351160 122898 351212
rect 118786 350548 118792 350600
rect 118844 350588 118850 350600
rect 178770 350588 178776 350600
rect 118844 350560 178776 350588
rect 118844 350548 118850 350560
rect 178770 350548 178776 350560
rect 178828 350548 178834 350600
rect 112438 349800 112444 349852
rect 112496 349840 112502 349852
rect 156046 349840 156052 349852
rect 112496 349812 156052 349840
rect 112496 349800 112502 349812
rect 156046 349800 156052 349812
rect 156104 349800 156110 349852
rect 128998 349120 129004 349172
rect 129056 349160 129062 349172
rect 180058 349160 180064 349172
rect 129056 349132 180064 349160
rect 129056 349120 129062 349132
rect 180058 349120 180064 349132
rect 180116 349120 180122 349172
rect 117222 347828 117228 347880
rect 117280 347868 117286 347880
rect 235258 347868 235264 347880
rect 117280 347840 235264 347868
rect 117280 347828 117286 347840
rect 235258 347828 235264 347840
rect 235316 347828 235322 347880
rect 89714 347760 89720 347812
rect 89772 347800 89778 347812
rect 91002 347800 91008 347812
rect 89772 347772 91008 347800
rect 89772 347760 89778 347772
rect 91002 347760 91008 347772
rect 91060 347800 91066 347812
rect 255406 347800 255412 347812
rect 91060 347772 255412 347800
rect 91060 347760 91066 347772
rect 255406 347760 255412 347772
rect 255464 347760 255470 347812
rect 3418 347012 3424 347064
rect 3476 347052 3482 347064
rect 78674 347052 78680 347064
rect 3476 347024 78680 347052
rect 3476 347012 3482 347024
rect 78674 347012 78680 347024
rect 78732 347052 78738 347064
rect 78732 347024 103514 347052
rect 78732 347012 78738 347024
rect 103486 346984 103514 347024
rect 124122 347012 124128 347064
rect 124180 347052 124186 347064
rect 140774 347052 140780 347064
rect 124180 347024 140780 347052
rect 124180 347012 124186 347024
rect 140774 347012 140780 347024
rect 140832 347012 140838 347064
rect 122926 346984 122932 346996
rect 103486 346956 122932 346984
rect 122926 346944 122932 346956
rect 122984 346944 122990 346996
rect 142798 346468 142804 346520
rect 142856 346508 142862 346520
rect 162118 346508 162124 346520
rect 142856 346480 162124 346508
rect 142856 346468 142862 346480
rect 162118 346468 162124 346480
rect 162176 346468 162182 346520
rect 101950 346400 101956 346452
rect 102008 346440 102014 346452
rect 221458 346440 221464 346452
rect 102008 346412 221464 346440
rect 102008 346400 102014 346412
rect 221458 346400 221464 346412
rect 221516 346400 221522 346452
rect 3142 346332 3148 346384
rect 3200 346372 3206 346384
rect 7558 346372 7564 346384
rect 3200 346344 7564 346372
rect 3200 346332 3206 346344
rect 7558 346332 7564 346344
rect 7616 346332 7622 346384
rect 74442 345652 74448 345704
rect 74500 345692 74506 345704
rect 89714 345692 89720 345704
rect 74500 345664 89720 345692
rect 74500 345652 74506 345664
rect 89714 345652 89720 345664
rect 89772 345652 89778 345704
rect 129826 345108 129832 345160
rect 129884 345148 129890 345160
rect 231118 345148 231124 345160
rect 129884 345120 231124 345148
rect 129884 345108 129890 345120
rect 231118 345108 231124 345120
rect 231176 345108 231182 345160
rect 84194 345040 84200 345092
rect 84252 345080 84258 345092
rect 85482 345080 85488 345092
rect 84252 345052 85488 345080
rect 84252 345040 84258 345052
rect 85482 345040 85488 345052
rect 85540 345080 85546 345092
rect 195238 345080 195244 345092
rect 85540 345052 195244 345080
rect 85540 345040 85546 345052
rect 195238 345040 195244 345052
rect 195296 345040 195302 345092
rect 90910 343680 90916 343732
rect 90968 343720 90974 343732
rect 211798 343720 211804 343732
rect 90968 343692 211804 343720
rect 90968 343680 90974 343692
rect 211798 343680 211804 343692
rect 211856 343680 211862 343732
rect 77202 343612 77208 343664
rect 77260 343652 77266 343664
rect 204346 343652 204352 343664
rect 77260 343624 204352 343652
rect 77260 343612 77266 343624
rect 204346 343612 204352 343624
rect 204404 343612 204410 343664
rect 79870 342864 79876 342916
rect 79928 342904 79934 342916
rect 88978 342904 88984 342916
rect 79928 342876 88984 342904
rect 79928 342864 79934 342876
rect 88978 342864 88984 342876
rect 89036 342864 89042 342916
rect 105538 342320 105544 342372
rect 105596 342360 105602 342372
rect 220078 342360 220084 342372
rect 105596 342332 220084 342360
rect 105596 342320 105602 342332
rect 220078 342320 220084 342332
rect 220136 342320 220142 342372
rect 93670 342252 93676 342304
rect 93728 342292 93734 342304
rect 251174 342292 251180 342304
rect 93728 342264 251180 342292
rect 93728 342252 93734 342264
rect 251174 342252 251180 342264
rect 251232 342252 251238 342304
rect 75822 341504 75828 341556
rect 75880 341544 75886 341556
rect 101490 341544 101496 341556
rect 75880 341516 101496 341544
rect 75880 341504 75886 341516
rect 101490 341504 101496 341516
rect 101548 341504 101554 341556
rect 142890 340960 142896 341012
rect 142948 341000 142954 341012
rect 160922 341000 160928 341012
rect 142948 340972 160928 341000
rect 142948 340960 142954 340972
rect 160922 340960 160928 340972
rect 160980 340960 160986 341012
rect 102686 340892 102692 340944
rect 102744 340932 102750 340944
rect 258166 340932 258172 340944
rect 102744 340904 258172 340932
rect 102744 340892 102750 340904
rect 258166 340892 258172 340904
rect 258224 340892 258230 340944
rect 77294 340212 77300 340264
rect 77352 340252 77358 340264
rect 93118 340252 93124 340264
rect 77352 340224 93124 340252
rect 77352 340212 77358 340224
rect 93118 340212 93124 340224
rect 93176 340212 93182 340264
rect 64598 340144 64604 340196
rect 64656 340184 64662 340196
rect 72418 340184 72424 340196
rect 64656 340156 72424 340184
rect 64656 340144 64662 340156
rect 72418 340144 72424 340156
rect 72476 340184 72482 340196
rect 134518 340184 134524 340196
rect 72476 340156 134524 340184
rect 72476 340144 72482 340156
rect 134518 340144 134524 340156
rect 134576 340144 134582 340196
rect 114462 339532 114468 339584
rect 114520 339572 114526 339584
rect 177482 339572 177488 339584
rect 114520 339544 177488 339572
rect 114520 339532 114526 339544
rect 177482 339532 177488 339544
rect 177540 339532 177546 339584
rect 134242 339464 134248 339516
rect 134300 339504 134306 339516
rect 236638 339504 236644 339516
rect 134300 339476 236644 339504
rect 134300 339464 134306 339476
rect 236638 339464 236644 339476
rect 236696 339464 236702 339516
rect 77110 338716 77116 338768
rect 77168 338756 77174 338768
rect 87598 338756 87604 338768
rect 77168 338728 87604 338756
rect 77168 338716 77174 338728
rect 87598 338716 87604 338728
rect 87656 338716 87662 338768
rect 106458 338172 106464 338224
rect 106516 338212 106522 338224
rect 191190 338212 191196 338224
rect 106516 338184 191196 338212
rect 106516 338172 106522 338184
rect 191190 338172 191196 338184
rect 191248 338172 191254 338224
rect 85666 338104 85672 338156
rect 85724 338144 85730 338156
rect 249978 338144 249984 338156
rect 85724 338116 249984 338144
rect 85724 338104 85730 338116
rect 249978 338104 249984 338116
rect 250036 338104 250042 338156
rect 63402 336812 63408 336864
rect 63460 336852 63466 336864
rect 163590 336852 163596 336864
rect 63460 336824 163596 336852
rect 63460 336812 63466 336824
rect 163590 336812 163596 336824
rect 163648 336812 163654 336864
rect 115934 336744 115940 336796
rect 115992 336784 115998 336796
rect 247310 336784 247316 336796
rect 115992 336756 247316 336784
rect 115992 336744 115998 336756
rect 247310 336744 247316 336756
rect 247368 336744 247374 336796
rect 66070 335996 66076 336048
rect 66128 336036 66134 336048
rect 74534 336036 74540 336048
rect 66128 336008 74540 336036
rect 66128 335996 66134 336008
rect 74534 335996 74540 336008
rect 74592 335996 74598 336048
rect 104894 335384 104900 335436
rect 104952 335424 104958 335436
rect 228450 335424 228456 335436
rect 104952 335396 228456 335424
rect 104952 335384 104958 335396
rect 228450 335384 228456 335396
rect 228508 335384 228514 335436
rect 67174 335316 67180 335368
rect 67232 335356 67238 335368
rect 206370 335356 206376 335368
rect 67232 335328 206376 335356
rect 67232 335316 67238 335328
rect 206370 335316 206376 335328
rect 206428 335316 206434 335368
rect 65978 334568 65984 334620
rect 66036 334608 66042 334620
rect 142890 334608 142896 334620
rect 66036 334580 142896 334608
rect 66036 334568 66042 334580
rect 142890 334568 142896 334580
rect 142948 334568 142954 334620
rect 144454 334024 144460 334076
rect 144512 334064 144518 334076
rect 160830 334064 160836 334076
rect 144512 334036 160836 334064
rect 144512 334024 144518 334036
rect 160830 334024 160836 334036
rect 160888 334024 160894 334076
rect 146202 333956 146208 334008
rect 146260 333996 146266 334008
rect 171778 333996 171784 334008
rect 146260 333968 171784 333996
rect 146260 333956 146266 333968
rect 171778 333956 171784 333968
rect 171836 333956 171842 334008
rect 115014 332704 115020 332716
rect 103486 332676 115020 332704
rect 67358 332596 67364 332648
rect 67416 332636 67422 332648
rect 67542 332636 67548 332648
rect 67416 332608 67548 332636
rect 67416 332596 67422 332608
rect 67542 332596 67548 332608
rect 67600 332636 67606 332648
rect 103486 332636 103514 332676
rect 115014 332664 115020 332676
rect 115072 332664 115078 332716
rect 141418 332664 141424 332716
rect 141476 332704 141482 332716
rect 158806 332704 158812 332716
rect 141476 332676 158812 332704
rect 141476 332664 141482 332676
rect 158806 332664 158812 332676
rect 158864 332664 158870 332716
rect 67600 332608 103514 332636
rect 67600 332596 67606 332608
rect 115658 332596 115664 332648
rect 115716 332636 115722 332648
rect 169202 332636 169208 332648
rect 115716 332608 169208 332636
rect 115716 332596 115722 332608
rect 169202 332596 169208 332608
rect 169260 332596 169266 332648
rect 86310 331848 86316 331900
rect 86368 331888 86374 331900
rect 97258 331888 97264 331900
rect 86368 331860 97264 331888
rect 86368 331848 86374 331860
rect 97258 331848 97264 331860
rect 97316 331848 97322 331900
rect 102502 331304 102508 331356
rect 102560 331344 102566 331356
rect 164970 331344 164976 331356
rect 102560 331316 164976 331344
rect 102560 331304 102566 331316
rect 164970 331304 164976 331316
rect 165028 331304 165034 331356
rect 49602 331236 49608 331288
rect 49660 331276 49666 331288
rect 83734 331276 83740 331288
rect 49660 331248 83740 331276
rect 49660 331236 49666 331248
rect 83734 331236 83740 331248
rect 83792 331236 83798 331288
rect 97902 331236 97908 331288
rect 97960 331276 97966 331288
rect 215938 331276 215944 331288
rect 97960 331248 215944 331276
rect 97960 331236 97966 331248
rect 215938 331236 215944 331248
rect 215996 331236 216002 331288
rect 159358 331168 159364 331220
rect 159416 331208 159422 331220
rect 161750 331208 161756 331220
rect 159416 331180 161756 331208
rect 159416 331168 159422 331180
rect 161750 331168 161756 331180
rect 161808 331168 161814 331220
rect 76466 331100 76472 331152
rect 76524 331140 76530 331152
rect 77110 331140 77116 331152
rect 76524 331112 77116 331140
rect 76524 331100 76530 331112
rect 77110 331100 77116 331112
rect 77168 331100 77174 331152
rect 95326 331100 95332 331152
rect 95384 331140 95390 331152
rect 95878 331140 95884 331152
rect 95384 331112 95884 331140
rect 95384 331100 95390 331112
rect 95878 331100 95884 331112
rect 95936 331100 95942 331152
rect 101490 331100 101496 331152
rect 101548 331140 101554 331152
rect 101950 331140 101956 331152
rect 101548 331112 101956 331140
rect 101548 331100 101554 331112
rect 101950 331100 101956 331112
rect 102008 331100 102014 331152
rect 107562 331100 107568 331152
rect 107620 331140 107626 331152
rect 108022 331140 108028 331152
rect 107620 331112 108028 331140
rect 107620 331100 107626 331112
rect 108022 331100 108028 331112
rect 108080 331100 108086 331152
rect 114370 331100 114376 331152
rect 114428 331140 114434 331152
rect 116578 331140 116584 331152
rect 114428 331112 116584 331140
rect 114428 331100 114434 331112
rect 116578 331100 116584 331112
rect 116636 331100 116642 331152
rect 117774 331100 117780 331152
rect 117832 331140 117838 331152
rect 118602 331140 118608 331152
rect 117832 331112 118608 331140
rect 117832 331100 117838 331112
rect 118602 331100 118608 331112
rect 118660 331100 118666 331152
rect 118694 331100 118700 331152
rect 118752 331140 118758 331152
rect 119430 331140 119436 331152
rect 118752 331112 119436 331140
rect 118752 331100 118758 331112
rect 119430 331100 119436 331112
rect 119488 331100 119494 331152
rect 122834 331100 122840 331152
rect 122892 331140 122898 331152
rect 123662 331140 123668 331152
rect 122892 331112 123668 331140
rect 122892 331100 122898 331112
rect 123662 331100 123668 331112
rect 123720 331100 123726 331152
rect 125594 331100 125600 331152
rect 125652 331140 125658 331152
rect 126422 331140 126428 331152
rect 125652 331112 126428 331140
rect 125652 331100 125658 331112
rect 126422 331100 126428 331112
rect 126480 331100 126486 331152
rect 137922 331100 137928 331152
rect 137980 331140 137986 331152
rect 139394 331140 139400 331152
rect 137980 331112 139400 331140
rect 137980 331100 137986 331112
rect 139394 331100 139400 331112
rect 139452 331100 139458 331152
rect 144178 331100 144184 331152
rect 144236 331140 144242 331152
rect 144822 331140 144828 331152
rect 144236 331112 144828 331140
rect 144236 331100 144242 331112
rect 144822 331100 144828 331112
rect 144880 331100 144886 331152
rect 95786 331032 95792 331084
rect 95844 331072 95850 331084
rect 96522 331072 96528 331084
rect 95844 331044 96528 331072
rect 95844 331032 95850 331044
rect 96522 331032 96528 331044
rect 96580 331032 96586 331084
rect 140682 331032 140688 331084
rect 140740 331072 140746 331084
rect 142798 331072 142804 331084
rect 140740 331044 142804 331072
rect 140740 331032 140746 331044
rect 142798 331032 142804 331044
rect 142856 331032 142862 331084
rect 144730 331032 144736 331084
rect 144788 331072 144794 331084
rect 146478 331072 146484 331084
rect 144788 331044 146484 331072
rect 144788 331032 144794 331044
rect 146478 331032 146484 331044
rect 146536 331032 146542 331084
rect 108298 330828 108304 330880
rect 108356 330868 108362 330880
rect 115198 330868 115204 330880
rect 108356 330840 115204 330868
rect 108356 330828 108362 330840
rect 115198 330828 115204 330840
rect 115256 330828 115262 330880
rect 196710 330556 196716 330608
rect 196768 330596 196774 330608
rect 251358 330596 251364 330608
rect 196768 330568 251364 330596
rect 196768 330556 196774 330568
rect 251358 330556 251364 330568
rect 251416 330556 251422 330608
rect 72234 330488 72240 330540
rect 72292 330528 72298 330540
rect 97902 330528 97908 330540
rect 72292 330500 97908 330528
rect 72292 330488 72298 330500
rect 97902 330488 97908 330500
rect 97960 330488 97966 330540
rect 115014 330488 115020 330540
rect 115072 330528 115078 330540
rect 140774 330528 140780 330540
rect 115072 330500 140780 330528
rect 115072 330488 115078 330500
rect 140774 330488 140780 330500
rect 140832 330488 140838 330540
rect 162118 330488 162124 330540
rect 162176 330528 162182 330540
rect 239490 330528 239496 330540
rect 162176 330500 239496 330528
rect 162176 330488 162182 330500
rect 239490 330488 239496 330500
rect 239548 330488 239554 330540
rect 110598 330352 110604 330404
rect 110656 330392 110662 330404
rect 111702 330392 111708 330404
rect 110656 330364 111708 330392
rect 110656 330352 110662 330364
rect 111702 330352 111708 330364
rect 111760 330352 111766 330404
rect 104250 330080 104256 330132
rect 104308 330120 104314 330132
rect 105538 330120 105544 330132
rect 104308 330092 105544 330120
rect 104308 330080 104314 330092
rect 105538 330080 105544 330092
rect 105596 330080 105602 330132
rect 127710 330080 127716 330132
rect 127768 330120 127774 330132
rect 128998 330120 129004 330132
rect 127768 330092 129004 330120
rect 127768 330080 127774 330092
rect 128998 330080 129004 330092
rect 129056 330080 129062 330132
rect 100018 330012 100024 330064
rect 100076 330052 100082 330064
rect 102778 330052 102784 330064
rect 100076 330024 102784 330052
rect 100076 330012 100082 330024
rect 102778 330012 102784 330024
rect 102836 330012 102842 330064
rect 79410 329944 79416 329996
rect 79468 329984 79474 329996
rect 79962 329984 79968 329996
rect 79468 329956 79968 329984
rect 79468 329944 79474 329956
rect 79962 329944 79968 329956
rect 80020 329944 80026 329996
rect 113634 329944 113640 329996
rect 113692 329984 113698 329996
rect 114462 329984 114468 329996
rect 113692 329956 114468 329984
rect 113692 329944 113698 329956
rect 114462 329944 114468 329956
rect 114520 329944 114526 329996
rect 153654 329876 153660 329928
rect 153712 329916 153718 329928
rect 159450 329916 159456 329928
rect 153712 329888 159456 329916
rect 153712 329876 153718 329888
rect 159450 329876 159456 329888
rect 159508 329876 159514 329928
rect 44082 329808 44088 329860
rect 44140 329848 44146 329860
rect 69106 329848 69112 329860
rect 44140 329820 69112 329848
rect 44140 329808 44146 329820
rect 69106 329808 69112 329820
rect 69164 329808 69170 329860
rect 91094 329808 91100 329860
rect 91152 329848 91158 329860
rect 111886 329848 111892 329860
rect 91152 329820 111892 329848
rect 91152 329808 91158 329820
rect 111886 329808 111892 329820
rect 111944 329808 111950 329860
rect 134150 329808 134156 329860
rect 134208 329848 134214 329860
rect 135070 329848 135076 329860
rect 134208 329820 135076 329848
rect 134208 329808 134214 329820
rect 135070 329808 135076 329820
rect 135128 329808 135134 329860
rect 135254 329808 135260 329860
rect 135312 329848 135318 329860
rect 135806 329848 135812 329860
rect 135312 329820 135812 329848
rect 135312 329808 135318 329820
rect 135806 329808 135812 329820
rect 135864 329808 135870 329860
rect 151630 329808 151636 329860
rect 151688 329848 151694 329860
rect 195422 329848 195428 329860
rect 151688 329820 195428 329848
rect 151688 329808 151694 329820
rect 195422 329808 195428 329820
rect 195480 329808 195486 329860
rect 134518 329128 134524 329180
rect 134576 329168 134582 329180
rect 196710 329168 196716 329180
rect 134576 329140 196716 329168
rect 134576 329128 134582 329140
rect 196710 329128 196716 329140
rect 196768 329128 196774 329180
rect 43438 329060 43444 329112
rect 43496 329100 43502 329112
rect 49510 329100 49516 329112
rect 43496 329072 49516 329100
rect 43496 329060 43502 329072
rect 49510 329060 49516 329072
rect 49568 329100 49574 329112
rect 135254 329100 135260 329112
rect 49568 329072 135260 329100
rect 49568 329060 49574 329072
rect 135254 329060 135260 329072
rect 135312 329060 135318 329112
rect 160922 329060 160928 329112
rect 160980 329100 160986 329112
rect 224218 329100 224224 329112
rect 160980 329072 224224 329100
rect 160980 329060 160986 329072
rect 224218 329060 224224 329072
rect 224276 329060 224282 329112
rect 36538 328448 36544 328500
rect 36596 328488 36602 328500
rect 124858 328488 124864 328500
rect 36596 328460 124864 328488
rect 36596 328448 36602 328460
rect 124858 328448 124864 328460
rect 124916 328448 124922 328500
rect 152090 328448 152096 328500
rect 152148 328488 152154 328500
rect 161014 328488 161020 328500
rect 152148 328460 161020 328488
rect 152148 328448 152154 328460
rect 161014 328448 161020 328460
rect 161072 328448 161078 328500
rect 213178 327768 213184 327820
rect 213236 327808 213242 327820
rect 248598 327808 248604 327820
rect 213236 327780 248604 327808
rect 213236 327768 213242 327780
rect 248598 327768 248604 327780
rect 248656 327768 248662 327820
rect 60550 327700 60556 327752
rect 60608 327740 60614 327752
rect 91094 327740 91100 327752
rect 60608 327712 91100 327740
rect 60608 327700 60614 327712
rect 91094 327700 91100 327712
rect 91152 327700 91158 327752
rect 158806 327700 158812 327752
rect 158864 327740 158870 327752
rect 185670 327740 185676 327752
rect 158864 327712 185676 327740
rect 158864 327700 158870 327712
rect 185670 327700 185676 327712
rect 185728 327700 185734 327752
rect 187050 327700 187056 327752
rect 187108 327740 187114 327752
rect 331214 327740 331220 327752
rect 187108 327712 331220 327740
rect 187108 327700 187114 327712
rect 331214 327700 331220 327712
rect 331272 327700 331278 327752
rect 33778 327156 33784 327208
rect 33836 327196 33842 327208
rect 114738 327196 114744 327208
rect 33836 327168 114744 327196
rect 33836 327156 33842 327168
rect 114738 327156 114744 327168
rect 114796 327156 114802 327208
rect 149882 327156 149888 327208
rect 149940 327196 149946 327208
rect 153654 327196 153660 327208
rect 149940 327168 153660 327196
rect 149940 327156 149946 327168
rect 153654 327156 153660 327168
rect 153712 327156 153718 327208
rect 154298 327156 154304 327208
rect 154356 327196 154362 327208
rect 158162 327196 158168 327208
rect 154356 327168 158168 327196
rect 154356 327156 154362 327168
rect 158162 327156 158168 327168
rect 158220 327156 158226 327208
rect 91554 327088 91560 327140
rect 91612 327128 91618 327140
rect 92382 327128 92388 327140
rect 91612 327100 92388 327128
rect 91612 327088 91618 327100
rect 92382 327088 92388 327100
rect 92440 327128 92446 327140
rect 180150 327128 180156 327140
rect 92440 327100 180156 327128
rect 92440 327088 92446 327100
rect 180150 327088 180156 327100
rect 180208 327088 180214 327140
rect 70026 327020 70032 327072
rect 70084 327060 70090 327072
rect 71038 327060 71044 327072
rect 70084 327032 71044 327060
rect 70084 327020 70090 327032
rect 71038 327020 71044 327032
rect 71096 327020 71102 327072
rect 139762 327020 139768 327072
rect 139820 327060 139826 327072
rect 151630 327060 151636 327072
rect 139820 327032 151636 327060
rect 139820 327020 139826 327032
rect 151630 327020 151636 327032
rect 151688 327020 151694 327072
rect 152826 326952 152832 327004
rect 152884 326992 152890 327004
rect 154206 326992 154212 327004
rect 152884 326964 154212 326992
rect 152884 326952 152890 326964
rect 154206 326952 154212 326964
rect 154264 326952 154270 327004
rect 68646 326884 68652 326936
rect 68704 326924 68710 326936
rect 71406 326924 71412 326936
rect 68704 326896 71412 326924
rect 68704 326884 68710 326896
rect 71406 326884 71412 326896
rect 71464 326884 71470 326936
rect 143442 326884 143448 326936
rect 143500 326884 143506 326936
rect 149146 326884 149152 326936
rect 149204 326924 149210 326936
rect 162210 326924 162216 326936
rect 149204 326896 162216 326924
rect 149204 326884 149210 326896
rect 162210 326884 162216 326896
rect 162268 326884 162274 326936
rect 66806 326816 66812 326868
rect 66864 326856 66870 326868
rect 68002 326856 68008 326868
rect 66864 326828 68008 326856
rect 66864 326816 66870 326828
rect 68002 326816 68008 326828
rect 68060 326816 68066 326868
rect 14 326340 20 326392
rect 72 326380 78 326392
rect 51718 326380 51724 326392
rect 72 326352 51724 326380
rect 72 326340 78 326352
rect 51718 326340 51724 326352
rect 51776 326340 51782 326392
rect 143460 325768 143488 326884
rect 161750 326340 161756 326392
rect 161808 326380 161814 326392
rect 177298 326380 177304 326392
rect 161808 326352 177304 326380
rect 161808 326340 161814 326352
rect 177298 326340 177304 326352
rect 177356 326340 177362 326392
rect 240778 325768 240784 325780
rect 143460 325740 240784 325768
rect 240778 325728 240784 325740
rect 240836 325728 240842 325780
rect 59170 325660 59176 325712
rect 59228 325700 59234 325712
rect 68094 325700 68100 325712
rect 59228 325672 68100 325700
rect 59228 325660 59234 325672
rect 68094 325660 68100 325672
rect 68152 325660 68158 325712
rect 161014 324980 161020 325032
rect 161072 325020 161078 325032
rect 258350 325020 258356 325032
rect 161072 324992 258356 325020
rect 161072 324980 161078 324992
rect 258350 324980 258356 324992
rect 258408 324980 258414 325032
rect 156046 324912 156052 324964
rect 156104 324952 156110 324964
rect 255498 324952 255504 324964
rect 156104 324924 255504 324952
rect 156104 324912 156110 324924
rect 255498 324912 255504 324924
rect 255556 324912 255562 324964
rect 56502 324300 56508 324352
rect 56560 324340 56566 324352
rect 66898 324340 66904 324352
rect 56560 324312 66904 324340
rect 56560 324300 56566 324312
rect 66898 324300 66904 324312
rect 66956 324300 66962 324352
rect 156138 324232 156144 324284
rect 156196 324272 156202 324284
rect 164234 324272 164240 324284
rect 156196 324244 164240 324272
rect 156196 324232 156202 324244
rect 164234 324232 164240 324244
rect 164292 324272 164298 324284
rect 172054 324272 172060 324284
rect 164292 324244 172060 324272
rect 164292 324232 164298 324244
rect 172054 324232 172060 324244
rect 172112 324232 172118 324284
rect 162302 323552 162308 323604
rect 162360 323592 162366 323604
rect 349154 323592 349160 323604
rect 162360 323564 349160 323592
rect 162360 323552 162366 323564
rect 349154 323552 349160 323564
rect 349212 323552 349218 323604
rect 156046 323416 156052 323468
rect 156104 323456 156110 323468
rect 162578 323456 162584 323468
rect 156104 323428 162584 323456
rect 156104 323416 156110 323428
rect 162578 323416 162584 323428
rect 162636 323416 162642 323468
rect 59262 322940 59268 322992
rect 59320 322980 59326 322992
rect 66714 322980 66720 322992
rect 59320 322952 66720 322980
rect 59320 322940 59326 322952
rect 66714 322940 66720 322952
rect 66772 322940 66778 322992
rect 154758 322532 154764 322584
rect 154816 322572 154822 322584
rect 155310 322572 155316 322584
rect 154816 322544 155316 322572
rect 154816 322532 154822 322544
rect 155310 322532 155316 322544
rect 155368 322532 155374 322584
rect 156046 321920 156052 321972
rect 156104 321960 156110 321972
rect 163498 321960 163504 321972
rect 156104 321932 163504 321960
rect 156104 321920 156110 321932
rect 163498 321920 163504 321932
rect 163556 321920 163562 321972
rect 54938 321580 54944 321632
rect 54996 321620 55002 321632
rect 64138 321620 64144 321632
rect 54996 321592 64144 321620
rect 54996 321580 55002 321592
rect 64138 321580 64144 321592
rect 64196 321620 64202 321632
rect 64196 321592 64874 321620
rect 64196 321580 64202 321592
rect 64846 321552 64874 321592
rect 154758 321580 154764 321632
rect 154816 321620 154822 321632
rect 243814 321620 243820 321632
rect 154816 321592 243820 321620
rect 154816 321580 154822 321592
rect 243814 321580 243820 321592
rect 243872 321580 243878 321632
rect 66622 321552 66628 321564
rect 64846 321524 66628 321552
rect 66622 321512 66628 321524
rect 66680 321512 66686 321564
rect 222930 320968 222936 321020
rect 222988 321008 222994 321020
rect 252646 321008 252652 321020
rect 222988 320980 252652 321008
rect 222988 320968 222994 320980
rect 252646 320968 252652 320980
rect 252704 320968 252710 321020
rect 204898 320900 204904 320952
rect 204956 320940 204962 320952
rect 238110 320940 238116 320952
rect 204956 320912 238116 320940
rect 204956 320900 204962 320912
rect 238110 320900 238116 320912
rect 238168 320900 238174 320952
rect 163590 320832 163596 320884
rect 163648 320872 163654 320884
rect 223022 320872 223028 320884
rect 163648 320844 223028 320872
rect 163648 320832 163654 320844
rect 223022 320832 223028 320844
rect 223080 320832 223086 320884
rect 156598 320152 156604 320204
rect 156656 320192 156662 320204
rect 195146 320192 195152 320204
rect 156656 320164 195152 320192
rect 156656 320152 156662 320164
rect 195146 320152 195152 320164
rect 195204 320152 195210 320204
rect 157242 319472 157248 319524
rect 157300 319512 157306 319524
rect 160094 319512 160100 319524
rect 157300 319484 160100 319512
rect 157300 319472 157306 319484
rect 160094 319472 160100 319484
rect 160152 319512 160158 319524
rect 199378 319512 199384 319524
rect 160152 319484 199384 319512
rect 160152 319472 160158 319484
rect 199378 319472 199384 319484
rect 199436 319472 199442 319524
rect 4062 319404 4068 319456
rect 4120 319444 4126 319456
rect 5442 319444 5448 319456
rect 4120 319416 5448 319444
rect 4120 319404 4126 319416
rect 5442 319404 5448 319416
rect 5500 319444 5506 319456
rect 29638 319444 29644 319456
rect 5500 319416 29644 319444
rect 5500 319404 5506 319416
rect 29638 319404 29644 319416
rect 29696 319404 29702 319456
rect 162578 319404 162584 319456
rect 162636 319444 162642 319456
rect 210418 319444 210424 319456
rect 162636 319416 210424 319444
rect 162636 319404 162642 319416
rect 210418 319404 210424 319416
rect 210476 319404 210482 319456
rect 64414 318792 64420 318844
rect 64472 318832 64478 318844
rect 66898 318832 66904 318844
rect 64472 318804 66904 318832
rect 64472 318792 64478 318804
rect 66898 318792 66904 318804
rect 66956 318792 66962 318844
rect 157242 318792 157248 318844
rect 157300 318832 157306 318844
rect 162118 318832 162124 318844
rect 157300 318804 162124 318832
rect 157300 318792 157306 318804
rect 162118 318792 162124 318804
rect 162176 318792 162182 318844
rect 210418 318792 210424 318844
rect 210476 318832 210482 318844
rect 258074 318832 258080 318844
rect 210476 318804 258080 318832
rect 210476 318792 210482 318804
rect 258074 318792 258080 318804
rect 258132 318792 258138 318844
rect 186958 318112 186964 318164
rect 187016 318152 187022 318164
rect 227622 318152 227628 318164
rect 187016 318124 227628 318152
rect 187016 318112 187022 318124
rect 227622 318112 227628 318124
rect 227680 318112 227686 318164
rect 3510 318044 3516 318096
rect 3568 318084 3574 318096
rect 46842 318084 46848 318096
rect 3568 318056 46848 318084
rect 3568 318044 3574 318056
rect 46842 318044 46848 318056
rect 46900 318044 46906 318096
rect 158162 318044 158168 318096
rect 158220 318084 158226 318096
rect 189902 318084 189908 318096
rect 158220 318056 189908 318084
rect 158220 318044 158226 318056
rect 189902 318044 189908 318056
rect 189960 318044 189966 318096
rect 195422 318044 195428 318096
rect 195480 318084 195486 318096
rect 242250 318084 242256 318096
rect 195480 318056 242256 318084
rect 195480 318044 195486 318056
rect 242250 318044 242256 318056
rect 242308 318044 242314 318096
rect 60642 317500 60648 317552
rect 60700 317540 60706 317552
rect 66898 317540 66904 317552
rect 60700 317512 66904 317540
rect 60700 317500 60706 317512
rect 66898 317500 66904 317512
rect 66956 317500 66962 317552
rect 46842 317432 46848 317484
rect 46900 317472 46906 317484
rect 66714 317472 66720 317484
rect 46900 317444 66720 317472
rect 46900 317432 46906 317444
rect 66714 317432 66720 317444
rect 66772 317432 66778 317484
rect 157242 316752 157248 316804
rect 157300 316792 157306 316804
rect 188430 316792 188436 316804
rect 157300 316764 188436 316792
rect 157300 316752 157306 316764
rect 188430 316752 188436 316764
rect 188488 316752 188494 316804
rect 166534 316684 166540 316736
rect 166592 316724 166598 316736
rect 305638 316724 305644 316736
rect 166592 316696 305644 316724
rect 166592 316684 166598 316696
rect 305638 316684 305644 316696
rect 305696 316684 305702 316736
rect 64782 315664 64788 315716
rect 64840 315704 64846 315716
rect 66990 315704 66996 315716
rect 64840 315676 66996 315704
rect 64840 315664 64846 315676
rect 66990 315664 66996 315676
rect 67048 315664 67054 315716
rect 155954 315324 155960 315376
rect 156012 315364 156018 315376
rect 171962 315364 171968 315376
rect 156012 315336 171968 315364
rect 156012 315324 156018 315336
rect 171962 315324 171968 315336
rect 172020 315324 172026 315376
rect 172054 315324 172060 315376
rect 172112 315364 172118 315376
rect 192478 315364 192484 315376
rect 172112 315336 192484 315364
rect 172112 315324 172118 315336
rect 192478 315324 192484 315336
rect 192536 315324 192542 315376
rect 163682 315256 163688 315308
rect 163740 315296 163746 315308
rect 244274 315296 244280 315308
rect 163740 315268 244280 315296
rect 163740 315256 163746 315268
rect 244274 315256 244280 315268
rect 244332 315256 244338 315308
rect 35158 314644 35164 314696
rect 35216 314684 35222 314696
rect 67542 314684 67548 314696
rect 35216 314656 67548 314684
rect 35216 314644 35222 314656
rect 67542 314644 67548 314656
rect 67600 314644 67606 314696
rect 217318 314644 217324 314696
rect 217376 314684 217382 314696
rect 217962 314684 217968 314696
rect 217376 314656 217968 314684
rect 217376 314644 217382 314656
rect 217962 314644 217968 314656
rect 218020 314684 218026 314696
rect 302234 314684 302240 314696
rect 218020 314656 302240 314684
rect 218020 314644 218026 314656
rect 302234 314644 302240 314656
rect 302292 314644 302298 314696
rect 178770 313964 178776 314016
rect 178828 314004 178834 314016
rect 235534 314004 235540 314016
rect 178828 313976 235540 314004
rect 178828 313964 178834 313976
rect 235534 313964 235540 313976
rect 235592 313964 235598 314016
rect 198090 313896 198096 313948
rect 198148 313936 198154 313948
rect 320174 313936 320180 313948
rect 198148 313908 320180 313936
rect 198148 313896 198154 313908
rect 320174 313896 320180 313908
rect 320232 313896 320238 313948
rect 61838 313284 61844 313336
rect 61896 313324 61902 313336
rect 65518 313324 65524 313336
rect 61896 313296 65524 313324
rect 61896 313284 61902 313296
rect 65518 313284 65524 313296
rect 65576 313284 65582 313336
rect 61930 313216 61936 313268
rect 61988 313256 61994 313268
rect 66898 313256 66904 313268
rect 61988 313228 66904 313256
rect 61988 313216 61994 313228
rect 66898 313216 66904 313228
rect 66956 313216 66962 313268
rect 166442 312604 166448 312656
rect 166500 312644 166506 312656
rect 230474 312644 230480 312656
rect 166500 312616 230480 312644
rect 166500 312604 166506 312616
rect 230474 312604 230480 312616
rect 230532 312604 230538 312656
rect 157334 312536 157340 312588
rect 157392 312576 157398 312588
rect 245654 312576 245660 312588
rect 157392 312548 245660 312576
rect 157392 312536 157398 312548
rect 245654 312536 245660 312548
rect 245712 312536 245718 312588
rect 157242 311856 157248 311908
rect 157300 311896 157306 311908
rect 166534 311896 166540 311908
rect 157300 311868 166540 311896
rect 157300 311856 157306 311868
rect 166534 311856 166540 311868
rect 166592 311856 166598 311908
rect 63402 311788 63408 311840
rect 63460 311828 63466 311840
rect 66898 311828 66904 311840
rect 63460 311800 66904 311828
rect 63460 311788 63466 311800
rect 66898 311788 66904 311800
rect 66956 311788 66962 311840
rect 214558 311176 214564 311228
rect 214616 311216 214622 311228
rect 227806 311216 227812 311228
rect 214616 311188 227812 311216
rect 214616 311176 214622 311188
rect 227806 311176 227812 311188
rect 227864 311176 227870 311228
rect 174722 311108 174728 311160
rect 174780 311148 174786 311160
rect 233970 311148 233976 311160
rect 174780 311120 233976 311148
rect 174780 311108 174786 311120
rect 233970 311108 233976 311120
rect 234028 311108 234034 311160
rect 157242 310496 157248 310548
rect 157300 310536 157306 310548
rect 166442 310536 166448 310548
rect 157300 310508 166448 310536
rect 157300 310496 157306 310508
rect 166442 310496 166448 310508
rect 166500 310496 166506 310548
rect 165062 309748 165068 309800
rect 165120 309788 165126 309800
rect 198090 309788 198096 309800
rect 165120 309760 198096 309788
rect 165120 309748 165126 309760
rect 198090 309748 198096 309760
rect 198148 309748 198154 309800
rect 197998 309204 198004 309256
rect 198056 309244 198062 309256
rect 198642 309244 198648 309256
rect 198056 309216 198648 309244
rect 198056 309204 198062 309216
rect 198642 309204 198648 309216
rect 198700 309244 198706 309256
rect 265618 309244 265624 309256
rect 198700 309216 265624 309244
rect 198700 309204 198706 309216
rect 265618 309204 265624 309216
rect 265676 309204 265682 309256
rect 63218 309136 63224 309188
rect 63276 309176 63282 309188
rect 66622 309176 66628 309188
rect 63276 309148 66628 309176
rect 63276 309136 63282 309148
rect 66622 309136 66628 309148
rect 66680 309136 66686 309188
rect 167730 309136 167736 309188
rect 167788 309176 167794 309188
rect 260834 309176 260840 309188
rect 167788 309148 260840 309176
rect 167788 309136 167794 309148
rect 260834 309136 260840 309148
rect 260892 309136 260898 309188
rect 50798 308388 50804 308440
rect 50856 308428 50862 308440
rect 67082 308428 67088 308440
rect 50856 308400 67088 308428
rect 50856 308388 50862 308400
rect 67082 308388 67088 308400
rect 67140 308388 67146 308440
rect 207658 307844 207664 307896
rect 207716 307884 207722 307896
rect 286318 307884 286324 307896
rect 207716 307856 286324 307884
rect 207716 307844 207722 307856
rect 286318 307844 286324 307856
rect 286376 307844 286382 307896
rect 11698 307776 11704 307828
rect 11756 307816 11762 307828
rect 50798 307816 50804 307828
rect 11756 307788 50804 307816
rect 11756 307776 11762 307788
rect 50798 307776 50804 307788
rect 50856 307776 50862 307828
rect 195330 307776 195336 307828
rect 195388 307816 195394 307828
rect 201678 307816 201684 307828
rect 195388 307788 201684 307816
rect 195388 307776 195394 307788
rect 201678 307776 201684 307788
rect 201736 307816 201742 307828
rect 583478 307816 583484 307828
rect 201736 307788 583484 307816
rect 201736 307776 201742 307788
rect 583478 307776 583484 307788
rect 583536 307776 583542 307828
rect 64598 307708 64604 307760
rect 64656 307748 64662 307760
rect 66530 307748 66536 307760
rect 64656 307720 66536 307748
rect 64656 307708 64662 307720
rect 66530 307708 66536 307720
rect 66588 307708 66594 307760
rect 22738 307028 22744 307080
rect 22796 307068 22802 307080
rect 67082 307068 67088 307080
rect 22796 307040 67088 307068
rect 22796 307028 22802 307040
rect 67082 307028 67088 307040
rect 67140 307028 67146 307080
rect 211798 306416 211804 306468
rect 211856 306456 211862 306468
rect 280890 306456 280896 306468
rect 211856 306428 280896 306456
rect 211856 306416 211862 306428
rect 280890 306416 280896 306428
rect 280948 306416 280954 306468
rect 156506 306348 156512 306400
rect 156564 306388 156570 306400
rect 318058 306388 318064 306400
rect 156564 306360 318064 306388
rect 156564 306348 156570 306360
rect 318058 306348 318064 306360
rect 318116 306348 318122 306400
rect 3510 306280 3516 306332
rect 3568 306320 3574 306332
rect 43438 306320 43444 306332
rect 3568 306292 43444 306320
rect 3568 306280 3574 306292
rect 43438 306280 43444 306292
rect 43496 306280 43502 306332
rect 64690 306280 64696 306332
rect 64748 306320 64754 306332
rect 66898 306320 66904 306332
rect 64748 306292 66904 306320
rect 64748 306280 64754 306292
rect 66898 306280 66904 306292
rect 66956 306280 66962 306332
rect 157242 306280 157248 306332
rect 157300 306320 157306 306332
rect 158714 306320 158720 306332
rect 157300 306292 158720 306320
rect 157300 306280 157306 306292
rect 158714 306280 158720 306292
rect 158772 306280 158778 306332
rect 162118 305600 162124 305652
rect 162176 305640 162182 305652
rect 245746 305640 245752 305652
rect 162176 305612 245752 305640
rect 162176 305600 162182 305612
rect 245746 305600 245752 305612
rect 245804 305600 245810 305652
rect 157242 305192 157248 305244
rect 157300 305232 157306 305244
rect 162302 305232 162308 305244
rect 157300 305204 162308 305232
rect 157300 305192 157306 305204
rect 162302 305192 162308 305204
rect 162360 305192 162366 305244
rect 198090 304988 198096 305040
rect 198148 305028 198154 305040
rect 198550 305028 198556 305040
rect 198148 305000 198556 305028
rect 198148 304988 198154 305000
rect 198550 304988 198556 305000
rect 198608 305028 198614 305040
rect 295334 305028 295340 305040
rect 198608 305000 295340 305028
rect 198608 304988 198614 305000
rect 295334 304988 295340 305000
rect 295392 304988 295398 305040
rect 221182 303696 221188 303748
rect 221240 303736 221246 303748
rect 271230 303736 271236 303748
rect 221240 303708 271236 303736
rect 221240 303696 221246 303708
rect 271230 303696 271236 303708
rect 271288 303696 271294 303748
rect 57882 303628 57888 303680
rect 57940 303668 57946 303680
rect 66898 303668 66904 303680
rect 57940 303640 66904 303668
rect 57940 303628 57946 303640
rect 66898 303628 66904 303640
rect 66956 303628 66962 303680
rect 156046 303628 156052 303680
rect 156104 303668 156110 303680
rect 213178 303668 213184 303680
rect 156104 303640 213184 303668
rect 156104 303628 156110 303640
rect 213178 303628 213184 303640
rect 213236 303628 213242 303680
rect 214742 303628 214748 303680
rect 214800 303668 214806 303680
rect 565078 303668 565084 303680
rect 214800 303640 565084 303668
rect 214800 303628 214806 303640
rect 565078 303628 565084 303640
rect 565136 303628 565142 303680
rect 60458 303560 60464 303612
rect 60516 303600 60522 303612
rect 66990 303600 66996 303612
rect 60516 303572 66996 303600
rect 60516 303560 60522 303572
rect 66990 303560 66996 303572
rect 67048 303560 67054 303612
rect 158714 302880 158720 302932
rect 158772 302920 158778 302932
rect 191190 302920 191196 302932
rect 158772 302892 191196 302920
rect 158772 302880 158778 302892
rect 191190 302880 191196 302892
rect 191248 302880 191254 302932
rect 220078 302268 220084 302320
rect 220136 302308 220142 302320
rect 220722 302308 220728 302320
rect 220136 302280 220728 302308
rect 220136 302268 220142 302280
rect 220722 302268 220728 302280
rect 220780 302308 220786 302320
rect 298186 302308 298192 302320
rect 220780 302280 298192 302308
rect 220780 302268 220786 302280
rect 298186 302268 298192 302280
rect 298244 302268 298250 302320
rect 157242 302200 157248 302252
rect 157300 302240 157306 302252
rect 243998 302240 244004 302252
rect 157300 302212 244004 302240
rect 157300 302200 157306 302212
rect 243998 302200 244004 302212
rect 244056 302200 244062 302252
rect 199470 302132 199476 302184
rect 199528 302172 199534 302184
rect 201402 302172 201408 302184
rect 199528 302144 201408 302172
rect 199528 302132 199534 302144
rect 201402 302132 201408 302144
rect 201460 302132 201466 302184
rect 166350 300908 166356 300960
rect 166408 300948 166414 300960
rect 208394 300948 208400 300960
rect 166408 300920 208400 300948
rect 166408 300908 166414 300920
rect 208394 300908 208400 300920
rect 208452 300908 208458 300960
rect 156782 300840 156788 300892
rect 156840 300880 156846 300892
rect 188338 300880 188344 300892
rect 156840 300852 188344 300880
rect 156840 300840 156846 300852
rect 188338 300840 188344 300852
rect 188396 300840 188402 300892
rect 201402 300840 201408 300892
rect 201460 300880 201466 300892
rect 276658 300880 276664 300892
rect 201460 300852 276664 300880
rect 201460 300840 201466 300852
rect 276658 300840 276664 300852
rect 276716 300840 276722 300892
rect 193950 299548 193956 299600
rect 194008 299588 194014 299600
rect 258258 299588 258264 299600
rect 194008 299560 258264 299588
rect 194008 299548 194014 299560
rect 258258 299548 258264 299560
rect 258316 299548 258322 299600
rect 56410 299480 56416 299532
rect 56468 299520 56474 299532
rect 66898 299520 66904 299532
rect 56468 299492 66904 299520
rect 56468 299480 56474 299492
rect 66898 299480 66904 299492
rect 66956 299480 66962 299532
rect 157150 299480 157156 299532
rect 157208 299520 157214 299532
rect 244918 299520 244924 299532
rect 157208 299492 244924 299520
rect 157208 299480 157214 299492
rect 244918 299480 244924 299492
rect 244976 299480 244982 299532
rect 157242 299412 157248 299464
rect 157300 299452 157306 299464
rect 166994 299452 167000 299464
rect 157300 299424 167000 299452
rect 157300 299412 157306 299424
rect 166994 299412 167000 299424
rect 167052 299412 167058 299464
rect 169202 298800 169208 298852
rect 169260 298840 169266 298852
rect 186958 298840 186964 298852
rect 169260 298812 186964 298840
rect 169260 298800 169266 298812
rect 186958 298800 186964 298812
rect 187016 298800 187022 298852
rect 166994 298732 167000 298784
rect 167052 298772 167058 298784
rect 225322 298772 225328 298784
rect 167052 298744 225328 298772
rect 167052 298732 167058 298744
rect 225322 298732 225328 298744
rect 225380 298732 225386 298784
rect 228358 298732 228364 298784
rect 228416 298772 228422 298784
rect 236178 298772 236184 298784
rect 228416 298744 236184 298772
rect 228416 298732 228422 298744
rect 236178 298732 236184 298744
rect 236236 298732 236242 298784
rect 195330 298188 195336 298240
rect 195388 298228 195394 298240
rect 252738 298228 252744 298240
rect 195388 298200 252744 298228
rect 195388 298188 195394 298200
rect 252738 298188 252744 298200
rect 252796 298188 252802 298240
rect 236178 298120 236184 298172
rect 236236 298160 236242 298172
rect 574738 298160 574744 298172
rect 236236 298132 574744 298160
rect 236236 298120 236242 298132
rect 574738 298120 574744 298132
rect 574796 298120 574802 298172
rect 236086 297304 236092 297356
rect 236144 297344 236150 297356
rect 236638 297344 236644 297356
rect 236144 297316 236644 297344
rect 236144 297304 236150 297316
rect 236638 297304 236644 297316
rect 236696 297304 236702 297356
rect 236638 296760 236644 296812
rect 236696 296800 236702 296812
rect 282914 296800 282920 296812
rect 236696 296772 282920 296800
rect 236696 296760 236702 296772
rect 282914 296760 282920 296772
rect 282972 296760 282978 296812
rect 163498 296692 163504 296744
rect 163556 296732 163562 296744
rect 238478 296732 238484 296744
rect 163556 296704 238484 296732
rect 163556 296692 163562 296704
rect 238478 296692 238484 296704
rect 238536 296692 238542 296744
rect 57698 296624 57704 296676
rect 57756 296664 57762 296676
rect 66898 296664 66904 296676
rect 57756 296636 66904 296664
rect 57756 296624 57762 296636
rect 66898 296624 66904 296636
rect 66956 296624 66962 296676
rect 156414 295944 156420 295996
rect 156472 295984 156478 295996
rect 244366 295984 244372 295996
rect 156472 295956 244372 295984
rect 156472 295944 156478 295956
rect 244366 295944 244372 295956
rect 244424 295944 244430 295996
rect 160002 295332 160008 295384
rect 160060 295372 160066 295384
rect 161566 295372 161572 295384
rect 160060 295344 161572 295372
rect 160060 295332 160066 295344
rect 161566 295332 161572 295344
rect 161624 295332 161630 295384
rect 196802 295332 196808 295384
rect 196860 295372 196866 295384
rect 259546 295372 259552 295384
rect 196860 295344 259552 295372
rect 196860 295332 196866 295344
rect 259546 295332 259552 295344
rect 259604 295332 259610 295384
rect 156322 295264 156328 295316
rect 156380 295304 156386 295316
rect 166350 295304 166356 295316
rect 156380 295276 166356 295304
rect 156380 295264 156386 295276
rect 166350 295264 166356 295276
rect 166408 295264 166414 295316
rect 166534 294584 166540 294636
rect 166592 294624 166598 294636
rect 245930 294624 245936 294636
rect 166592 294596 245936 294624
rect 166592 294584 166598 294596
rect 245930 294584 245936 294596
rect 245988 294584 245994 294636
rect 154850 293972 154856 294024
rect 154908 294012 154914 294024
rect 248690 294012 248696 294024
rect 154908 293984 248696 294012
rect 154908 293972 154914 293984
rect 248690 293972 248696 293984
rect 248748 293972 248754 294024
rect 59078 293904 59084 293956
rect 59136 293944 59142 293956
rect 66990 293944 66996 293956
rect 59136 293916 66996 293944
rect 59136 293904 59142 293916
rect 66990 293904 66996 293916
rect 67048 293904 67054 293956
rect 213178 293224 213184 293276
rect 213236 293264 213242 293276
rect 235994 293264 236000 293276
rect 213236 293236 236000 293264
rect 213236 293224 213242 293236
rect 235994 293224 236000 293236
rect 236052 293224 236058 293276
rect 2774 292816 2780 292868
rect 2832 292856 2838 292868
rect 4798 292856 4804 292868
rect 2832 292828 4804 292856
rect 2832 292816 2838 292828
rect 4798 292816 4804 292828
rect 4856 292816 4862 292868
rect 48038 292544 48044 292596
rect 48096 292584 48102 292596
rect 66714 292584 66720 292596
rect 48096 292556 66720 292584
rect 48096 292544 48102 292556
rect 66714 292544 66720 292556
rect 66772 292544 66778 292596
rect 157242 292544 157248 292596
rect 157300 292584 157306 292596
rect 220630 292584 220636 292596
rect 157300 292556 220636 292584
rect 157300 292544 157306 292556
rect 220630 292544 220636 292556
rect 220688 292584 220694 292596
rect 255314 292584 255320 292596
rect 220688 292556 255320 292584
rect 220688 292544 220694 292556
rect 255314 292544 255320 292556
rect 255372 292544 255378 292596
rect 14458 292476 14464 292528
rect 14516 292516 14522 292528
rect 62022 292516 62028 292528
rect 14516 292488 62028 292516
rect 14516 292476 14522 292488
rect 62022 292476 62028 292488
rect 62080 292516 62086 292528
rect 66898 292516 66904 292528
rect 62080 292488 66904 292516
rect 62080 292476 62086 292488
rect 66898 292476 66904 292488
rect 66956 292476 66962 292528
rect 162210 291796 162216 291848
rect 162268 291836 162274 291848
rect 173434 291836 173440 291848
rect 162268 291808 173440 291836
rect 162268 291796 162274 291808
rect 173434 291796 173440 291808
rect 173492 291796 173498 291848
rect 201402 291796 201408 291848
rect 201460 291836 201466 291848
rect 218054 291836 218060 291848
rect 201460 291808 218060 291836
rect 201460 291796 201466 291808
rect 218054 291796 218060 291808
rect 218112 291796 218118 291848
rect 217870 291252 217876 291304
rect 217928 291292 217934 291304
rect 218146 291292 218152 291304
rect 217928 291264 218152 291292
rect 217928 291252 217934 291264
rect 218146 291252 218152 291264
rect 218204 291252 218210 291304
rect 233970 291252 233976 291304
rect 234028 291292 234034 291304
rect 289906 291292 289912 291304
rect 234028 291264 289912 291292
rect 234028 291252 234034 291264
rect 289906 291252 289912 291264
rect 289964 291252 289970 291304
rect 156782 291184 156788 291236
rect 156840 291224 156846 291236
rect 159634 291224 159640 291236
rect 156840 291196 159640 291224
rect 156840 291184 156846 291196
rect 159634 291184 159640 291196
rect 159692 291184 159698 291236
rect 167822 291184 167828 291236
rect 167880 291224 167886 291236
rect 256786 291224 256792 291236
rect 167880 291196 256792 291224
rect 167880 291184 167886 291196
rect 256786 291184 256792 291196
rect 256844 291184 256850 291236
rect 200390 291116 200396 291168
rect 200448 291156 200454 291168
rect 204254 291156 204260 291168
rect 200448 291128 204260 291156
rect 200448 291116 200454 291128
rect 204254 291116 204260 291128
rect 204312 291156 204318 291168
rect 582558 291156 582564 291168
rect 204312 291128 582564 291156
rect 204312 291116 204318 291128
rect 582558 291116 582564 291128
rect 582616 291116 582622 291168
rect 239398 291048 239404 291100
rect 239456 291088 239462 291100
rect 242342 291088 242348 291100
rect 239456 291060 242348 291088
rect 239456 291048 239462 291060
rect 242342 291048 242348 291060
rect 242400 291048 242406 291100
rect 182910 290436 182916 290488
rect 182968 290476 182974 290488
rect 193950 290476 193956 290488
rect 182968 290448 193956 290476
rect 182968 290436 182974 290448
rect 193950 290436 193956 290448
rect 194008 290436 194014 290488
rect 197354 290436 197360 290488
rect 197412 290476 197418 290488
rect 239950 290476 239956 290488
rect 197412 290448 239956 290476
rect 197412 290436 197418 290448
rect 239950 290436 239956 290448
rect 240008 290436 240014 290488
rect 63310 289892 63316 289944
rect 63368 289932 63374 289944
rect 66898 289932 66904 289944
rect 63368 289904 66904 289932
rect 63368 289892 63374 289904
rect 66898 289892 66904 289904
rect 66956 289892 66962 289944
rect 242342 289824 242348 289876
rect 242400 289864 242406 289876
rect 264238 289864 264244 289876
rect 242400 289836 264244 289864
rect 242400 289824 242406 289836
rect 264238 289824 264244 289836
rect 264296 289824 264302 289876
rect 232498 289756 232504 289808
rect 232556 289796 232562 289808
rect 234614 289796 234620 289808
rect 232556 289768 234620 289796
rect 232556 289756 232562 289768
rect 234614 289756 234620 289768
rect 234672 289756 234678 289808
rect 242158 289756 242164 289808
rect 242216 289796 242222 289808
rect 242894 289796 242900 289808
rect 242216 289768 242900 289796
rect 242216 289756 242222 289768
rect 242894 289756 242900 289768
rect 242952 289756 242958 289808
rect 60550 289348 60556 289400
rect 60608 289388 60614 289400
rect 66898 289388 66904 289400
rect 60608 289360 66904 289388
rect 60608 289348 60614 289360
rect 66898 289348 66904 289360
rect 66956 289348 66962 289400
rect 52178 289076 52184 289128
rect 52236 289116 52242 289128
rect 67174 289116 67180 289128
rect 52236 289088 67180 289116
rect 52236 289076 52242 289088
rect 67174 289076 67180 289088
rect 67232 289076 67238 289128
rect 187142 288464 187148 288516
rect 187200 288504 187206 288516
rect 230566 288504 230572 288516
rect 187200 288476 230572 288504
rect 187200 288464 187206 288476
rect 230566 288464 230572 288476
rect 230624 288464 230630 288516
rect 156782 288396 156788 288448
rect 156840 288436 156846 288448
rect 224494 288436 224500 288448
rect 156840 288408 224500 288436
rect 156840 288396 156846 288408
rect 224494 288396 224500 288408
rect 224552 288396 224558 288448
rect 237926 288396 237932 288448
rect 237984 288436 237990 288448
rect 238110 288436 238116 288448
rect 237984 288408 238116 288436
rect 237984 288396 237990 288408
rect 238110 288396 238116 288408
rect 238168 288436 238174 288448
rect 264330 288436 264336 288448
rect 238168 288408 264336 288436
rect 238168 288396 238174 288408
rect 264330 288396 264336 288408
rect 264388 288396 264394 288448
rect 156230 287104 156236 287156
rect 156288 287144 156294 287156
rect 231302 287144 231308 287156
rect 156288 287116 231308 287144
rect 156288 287104 156294 287116
rect 231302 287104 231308 287116
rect 231360 287104 231366 287156
rect 238110 287104 238116 287156
rect 238168 287144 238174 287156
rect 267090 287144 267096 287156
rect 238168 287116 267096 287144
rect 238168 287104 238174 287116
rect 267090 287104 267096 287116
rect 267148 287104 267154 287156
rect 64690 287036 64696 287088
rect 64748 287076 64754 287088
rect 66714 287076 66720 287088
rect 64748 287048 66720 287076
rect 64748 287036 64754 287048
rect 66714 287036 66720 287048
rect 66772 287036 66778 287088
rect 156322 287036 156328 287088
rect 156380 287076 156386 287088
rect 244458 287076 244464 287088
rect 156380 287048 244464 287076
rect 156380 287036 156386 287048
rect 244458 287036 244464 287048
rect 244516 287036 244522 287088
rect 240778 286492 240784 286544
rect 240836 286532 240842 286544
rect 241974 286532 241980 286544
rect 240836 286504 241980 286532
rect 240836 286492 240842 286504
rect 241974 286492 241980 286504
rect 242032 286492 242038 286544
rect 217962 286424 217968 286476
rect 218020 286464 218026 286476
rect 221550 286464 221556 286476
rect 218020 286436 221556 286464
rect 218020 286424 218026 286436
rect 221550 286424 221556 286436
rect 221608 286424 221614 286476
rect 224218 286220 224224 286272
rect 224276 286260 224282 286272
rect 225046 286260 225052 286272
rect 224276 286232 225052 286260
rect 224276 286220 224282 286232
rect 225046 286220 225052 286232
rect 225104 286220 225110 286272
rect 63402 285744 63408 285796
rect 63460 285784 63466 285796
rect 66898 285784 66904 285796
rect 63460 285756 66904 285784
rect 63460 285744 63466 285756
rect 66898 285744 66904 285756
rect 66956 285744 66962 285796
rect 199378 285744 199384 285796
rect 199436 285784 199442 285796
rect 205542 285784 205548 285796
rect 199436 285756 205548 285784
rect 199436 285744 199442 285756
rect 205542 285744 205548 285756
rect 205600 285744 205606 285796
rect 213822 285744 213828 285796
rect 213880 285784 213886 285796
rect 215386 285784 215392 285796
rect 213880 285756 215392 285784
rect 213880 285744 213886 285756
rect 215386 285744 215392 285756
rect 215444 285744 215450 285796
rect 223574 285784 223580 285796
rect 219406 285756 223580 285784
rect 55122 285676 55128 285728
rect 55180 285716 55186 285728
rect 66806 285716 66812 285728
rect 55180 285688 66812 285716
rect 55180 285676 55186 285688
rect 66806 285676 66812 285688
rect 66864 285676 66870 285728
rect 157242 285676 157248 285728
rect 157300 285716 157306 285728
rect 166350 285716 166356 285728
rect 157300 285688 166356 285716
rect 157300 285676 157306 285688
rect 166350 285676 166356 285688
rect 166408 285676 166414 285728
rect 169294 285676 169300 285728
rect 169352 285716 169358 285728
rect 173250 285716 173256 285728
rect 169352 285688 173256 285716
rect 169352 285676 169358 285688
rect 173250 285676 173256 285688
rect 173308 285676 173314 285728
rect 194042 285676 194048 285728
rect 194100 285716 194106 285728
rect 204622 285716 204628 285728
rect 194100 285688 204628 285716
rect 194100 285676 194106 285688
rect 204622 285676 204628 285688
rect 204680 285676 204686 285728
rect 206370 285676 206376 285728
rect 206428 285716 206434 285728
rect 207014 285716 207020 285728
rect 206428 285688 207020 285716
rect 206428 285676 206434 285688
rect 207014 285676 207020 285688
rect 207072 285676 207078 285728
rect 214558 285676 214564 285728
rect 214616 285716 214622 285728
rect 219406 285716 219434 285756
rect 223574 285744 223580 285756
rect 223632 285744 223638 285796
rect 227622 285744 227628 285796
rect 227680 285784 227686 285796
rect 228910 285784 228916 285796
rect 227680 285756 228916 285784
rect 227680 285744 227686 285756
rect 228910 285744 228916 285756
rect 228968 285744 228974 285796
rect 231118 285744 231124 285796
rect 231176 285784 231182 285796
rect 232222 285784 232228 285796
rect 231176 285756 232228 285784
rect 231176 285744 231182 285756
rect 232222 285744 232228 285756
rect 232280 285784 232286 285796
rect 251818 285784 251824 285796
rect 232280 285756 251824 285784
rect 232280 285744 232286 285756
rect 251818 285744 251824 285756
rect 251876 285744 251882 285796
rect 214616 285688 219434 285716
rect 214616 285676 214622 285688
rect 219710 285676 219716 285728
rect 219768 285716 219774 285728
rect 220722 285716 220728 285728
rect 219768 285688 220728 285716
rect 219768 285676 219774 285688
rect 220722 285676 220728 285688
rect 220780 285676 220786 285728
rect 222838 285676 222844 285728
rect 222896 285716 222902 285728
rect 226518 285716 226524 285728
rect 222896 285688 226524 285716
rect 222896 285676 222902 285688
rect 226518 285676 226524 285688
rect 226576 285676 226582 285728
rect 228450 285676 228456 285728
rect 228508 285716 228514 285728
rect 229278 285716 229284 285728
rect 228508 285688 229284 285716
rect 228508 285676 228514 285688
rect 229278 285676 229284 285688
rect 229336 285676 229342 285728
rect 233142 285676 233148 285728
rect 233200 285716 233206 285728
rect 233878 285716 233884 285728
rect 233200 285688 233884 285716
rect 233200 285676 233206 285688
rect 233878 285676 233884 285688
rect 233936 285676 233942 285728
rect 200114 285268 200120 285320
rect 200172 285308 200178 285320
rect 200482 285308 200488 285320
rect 200172 285280 200488 285308
rect 200172 285268 200178 285280
rect 200482 285268 200488 285280
rect 200540 285268 200546 285320
rect 208394 285268 208400 285320
rect 208452 285308 208458 285320
rect 208670 285308 208676 285320
rect 208452 285280 208676 285308
rect 208452 285268 208458 285280
rect 208670 285268 208676 285280
rect 208728 285268 208734 285320
rect 218146 285268 218152 285320
rect 218204 285308 218210 285320
rect 218330 285308 218336 285320
rect 218204 285280 218336 285308
rect 218204 285268 218210 285280
rect 218330 285268 218336 285280
rect 218388 285268 218394 285320
rect 192570 284928 192576 284980
rect 192628 284968 192634 284980
rect 214558 284968 214564 284980
rect 192628 284940 214564 284968
rect 192628 284928 192634 284940
rect 214558 284928 214564 284940
rect 214616 284928 214622 284980
rect 216766 284384 216772 284436
rect 216824 284424 216830 284436
rect 248414 284424 248420 284436
rect 216824 284396 248420 284424
rect 216824 284384 216830 284396
rect 248414 284384 248420 284396
rect 248472 284384 248478 284436
rect 157242 284316 157248 284368
rect 157300 284356 157306 284368
rect 247034 284356 247040 284368
rect 157300 284328 247040 284356
rect 157300 284316 157306 284328
rect 247034 284316 247040 284328
rect 247092 284316 247098 284368
rect 180150 284248 180156 284300
rect 180208 284288 180214 284300
rect 197354 284288 197360 284300
rect 180208 284260 197360 284288
rect 180208 284248 180214 284260
rect 197354 284248 197360 284260
rect 197412 284248 197418 284300
rect 242250 283908 242256 283960
rect 242308 283948 242314 283960
rect 242308 283920 248414 283948
rect 242308 283908 242314 283920
rect 248386 283880 248414 283920
rect 313274 283880 313280 283892
rect 248386 283852 313280 283880
rect 313274 283840 313280 283852
rect 313332 283840 313338 283892
rect 177298 283568 177304 283620
rect 177356 283608 177362 283620
rect 185762 283608 185768 283620
rect 177356 283580 185768 283608
rect 177356 283568 177362 283580
rect 185762 283568 185768 283580
rect 185820 283568 185826 283620
rect 246390 283568 246396 283620
rect 246448 283608 246454 283620
rect 247310 283608 247316 283620
rect 246448 283580 247316 283608
rect 246448 283568 246454 283580
rect 247310 283568 247316 283580
rect 247368 283608 247374 283620
rect 252830 283608 252836 283620
rect 247368 283580 252836 283608
rect 247368 283568 247374 283580
rect 252830 283568 252836 283580
rect 252888 283568 252894 283620
rect 39942 282888 39948 282940
rect 40000 282928 40006 282940
rect 66714 282928 66720 282940
rect 40000 282900 66720 282928
rect 40000 282888 40006 282900
rect 66714 282888 66720 282900
rect 66772 282888 66778 282940
rect 157242 282888 157248 282940
rect 157300 282928 157306 282940
rect 179506 282928 179512 282940
rect 157300 282900 179512 282928
rect 157300 282888 157306 282900
rect 179506 282888 179512 282900
rect 179564 282888 179570 282940
rect 157150 282820 157156 282872
rect 157208 282860 157214 282872
rect 182910 282860 182916 282872
rect 157208 282832 182916 282860
rect 157208 282820 157214 282832
rect 182910 282820 182916 282832
rect 182968 282820 182974 282872
rect 246114 282820 246120 282872
rect 246172 282860 246178 282872
rect 252554 282860 252560 282872
rect 246172 282832 252560 282860
rect 246172 282820 246178 282832
rect 252554 282820 252560 282832
rect 252612 282860 252618 282872
rect 582742 282860 582748 282872
rect 252612 282832 582748 282860
rect 252612 282820 252618 282832
rect 582742 282820 582748 282832
rect 582800 282820 582806 282872
rect 179506 282140 179512 282192
rect 179564 282180 179570 282192
rect 180702 282180 180708 282192
rect 179564 282152 180708 282180
rect 179564 282140 179570 282152
rect 180702 282140 180708 282152
rect 180760 282180 180766 282192
rect 197354 282180 197360 282192
rect 180760 282152 197360 282180
rect 180760 282140 180766 282152
rect 197354 282140 197360 282152
rect 197412 282140 197418 282192
rect 245930 281664 245936 281716
rect 245988 281704 245994 281716
rect 250070 281704 250076 281716
rect 245988 281676 250076 281704
rect 245988 281664 245994 281676
rect 250070 281664 250076 281676
rect 250128 281664 250134 281716
rect 52270 281528 52276 281580
rect 52328 281568 52334 281580
rect 66346 281568 66352 281580
rect 52328 281540 66352 281568
rect 52328 281528 52334 281540
rect 66346 281528 66352 281540
rect 66404 281528 66410 281580
rect 157242 281460 157248 281512
rect 157300 281500 157306 281512
rect 196802 281500 196808 281512
rect 157300 281472 196808 281500
rect 157300 281460 157306 281472
rect 196802 281460 196808 281472
rect 196860 281460 196866 281512
rect 246114 281460 246120 281512
rect 246172 281500 246178 281512
rect 258350 281500 258356 281512
rect 246172 281472 258356 281500
rect 246172 281460 246178 281472
rect 258350 281460 258356 281472
rect 258408 281500 258414 281512
rect 259362 281500 259368 281512
rect 258408 281472 259368 281500
rect 258408 281460 258414 281472
rect 259362 281460 259368 281472
rect 259420 281460 259426 281512
rect 171870 281392 171876 281444
rect 171928 281432 171934 281444
rect 177298 281432 177304 281444
rect 171928 281404 177304 281432
rect 171928 281392 171934 281404
rect 177298 281392 177304 281404
rect 177356 281392 177362 281444
rect 191190 281392 191196 281444
rect 191248 281432 191254 281444
rect 197354 281432 197360 281444
rect 191248 281404 197360 281432
rect 191248 281392 191254 281404
rect 197354 281392 197360 281404
rect 197412 281392 197418 281444
rect 259362 280848 259368 280900
rect 259420 280888 259426 280900
rect 271138 280888 271144 280900
rect 259420 280860 271144 280888
rect 259420 280848 259426 280860
rect 271138 280848 271144 280860
rect 271196 280848 271202 280900
rect 157058 280780 157064 280832
rect 157116 280820 157122 280832
rect 167822 280820 167828 280832
rect 157116 280792 167828 280820
rect 157116 280780 157122 280792
rect 167822 280780 167828 280792
rect 167880 280780 167886 280832
rect 245930 280780 245936 280832
rect 245988 280820 245994 280832
rect 248506 280820 248512 280832
rect 245988 280792 248512 280820
rect 245988 280780 245994 280792
rect 248506 280780 248512 280792
rect 248564 280820 248570 280832
rect 273898 280820 273904 280832
rect 248564 280792 273904 280820
rect 248564 280780 248570 280792
rect 273898 280780 273904 280792
rect 273956 280780 273962 280832
rect 59078 280168 59084 280220
rect 59136 280208 59142 280220
rect 66806 280208 66812 280220
rect 59136 280180 66812 280208
rect 59136 280168 59142 280180
rect 66806 280168 66812 280180
rect 66864 280168 66870 280220
rect 245930 279828 245936 279880
rect 245988 279868 245994 279880
rect 249886 279868 249892 279880
rect 245988 279840 249892 279868
rect 245988 279828 245994 279840
rect 249886 279828 249892 279840
rect 249944 279868 249950 279880
rect 251082 279868 251088 279880
rect 249944 279840 251088 279868
rect 249944 279828 249950 279840
rect 251082 279828 251088 279840
rect 251140 279828 251146 279880
rect 162302 279420 162308 279472
rect 162360 279460 162366 279472
rect 191742 279460 191748 279472
rect 162360 279432 191748 279460
rect 162360 279420 162366 279432
rect 191742 279420 191748 279432
rect 191800 279460 191806 279472
rect 197446 279460 197452 279472
rect 191800 279432 197452 279460
rect 191800 279420 191806 279432
rect 197446 279420 197452 279432
rect 197504 279420 197510 279472
rect 251082 279420 251088 279472
rect 251140 279460 251146 279472
rect 583570 279460 583576 279472
rect 251140 279432 583576 279460
rect 251140 279420 251146 279432
rect 583570 279420 583576 279432
rect 583628 279420 583634 279472
rect 157242 279012 157248 279064
rect 157300 279052 157306 279064
rect 161382 279052 161388 279064
rect 157300 279024 161388 279052
rect 157300 279012 157306 279024
rect 161382 279012 161388 279024
rect 161440 279012 161446 279064
rect 156966 278808 156972 278860
rect 157024 278848 157030 278860
rect 160094 278848 160100 278860
rect 157024 278820 160100 278848
rect 157024 278808 157030 278820
rect 160094 278808 160100 278820
rect 160152 278808 160158 278860
rect 14458 278740 14464 278792
rect 14516 278780 14522 278792
rect 60458 278780 60464 278792
rect 14516 278752 60464 278780
rect 14516 278740 14522 278752
rect 60458 278740 60464 278752
rect 60516 278780 60522 278792
rect 67266 278780 67272 278792
rect 60516 278752 67272 278780
rect 60516 278740 60522 278752
rect 67266 278740 67272 278752
rect 67324 278740 67330 278792
rect 245930 278672 245936 278724
rect 245988 278712 245994 278724
rect 254118 278712 254124 278724
rect 245988 278684 254124 278712
rect 245988 278672 245994 278684
rect 254118 278672 254124 278684
rect 254176 278672 254182 278724
rect 181438 277992 181444 278044
rect 181496 278032 181502 278044
rect 197354 278032 197360 278044
rect 181496 278004 197360 278032
rect 181496 277992 181502 278004
rect 197354 277992 197360 278004
rect 197412 277992 197418 278044
rect 254118 277992 254124 278044
rect 254176 278032 254182 278044
rect 583294 278032 583300 278044
rect 254176 278004 583300 278032
rect 254176 277992 254182 278004
rect 583294 277992 583300 278004
rect 583352 277992 583358 278044
rect 191834 277788 191840 277840
rect 191892 277828 191898 277840
rect 197446 277828 197452 277840
rect 191892 277800 197452 277828
rect 191892 277788 191898 277800
rect 197446 277788 197452 277800
rect 197504 277788 197510 277840
rect 54846 277380 54852 277432
rect 54904 277420 54910 277432
rect 66714 277420 66720 277432
rect 54904 277392 66720 277420
rect 54904 277380 54910 277392
rect 66714 277380 66720 277392
rect 66772 277380 66778 277432
rect 157242 277380 157248 277432
rect 157300 277420 157306 277432
rect 166534 277420 166540 277432
rect 157300 277392 166540 277420
rect 157300 277380 157306 277392
rect 166534 277380 166540 277392
rect 166592 277380 166598 277432
rect 186958 277380 186964 277432
rect 187016 277420 187022 277432
rect 191834 277420 191840 277432
rect 187016 277392 191840 277420
rect 187016 277380 187022 277392
rect 191834 277380 191840 277392
rect 191892 277380 191898 277432
rect 185762 276700 185768 276752
rect 185820 276740 185826 276752
rect 197538 276740 197544 276752
rect 185820 276712 197544 276740
rect 185820 276700 185826 276712
rect 197538 276700 197544 276712
rect 197596 276700 197602 276752
rect 160094 276632 160100 276684
rect 160152 276672 160158 276684
rect 194502 276672 194508 276684
rect 160152 276644 194508 276672
rect 160152 276632 160158 276644
rect 194502 276632 194508 276644
rect 194560 276672 194566 276684
rect 197354 276672 197360 276684
rect 194560 276644 197360 276672
rect 194560 276632 194566 276644
rect 197354 276632 197360 276644
rect 197412 276632 197418 276684
rect 245746 276632 245752 276684
rect 245804 276672 245810 276684
rect 278038 276672 278044 276684
rect 245804 276644 278044 276672
rect 245804 276632 245810 276644
rect 278038 276632 278044 276644
rect 278096 276632 278102 276684
rect 177482 276496 177488 276548
rect 177540 276536 177546 276548
rect 181530 276536 181536 276548
rect 177540 276508 181536 276536
rect 177540 276496 177546 276508
rect 181530 276496 181536 276508
rect 181588 276496 181594 276548
rect 156874 276020 156880 276072
rect 156932 276060 156938 276072
rect 167822 276060 167828 276072
rect 156932 276032 167828 276060
rect 156932 276020 156938 276032
rect 167822 276020 167828 276032
rect 167880 276020 167886 276072
rect 245930 275952 245936 276004
rect 245988 275992 245994 276004
rect 253934 275992 253940 276004
rect 245988 275964 253940 275992
rect 245988 275952 245994 275964
rect 253934 275952 253940 275964
rect 253992 275992 253998 276004
rect 582650 275992 582656 276004
rect 253992 275964 582656 275992
rect 253992 275952 253998 275964
rect 582650 275952 582656 275964
rect 582708 275952 582714 276004
rect 186958 275340 186964 275392
rect 187016 275380 187022 275392
rect 199654 275380 199660 275392
rect 187016 275352 199660 275380
rect 187016 275340 187022 275352
rect 199654 275340 199660 275352
rect 199712 275340 199718 275392
rect 166442 275272 166448 275324
rect 166500 275312 166506 275324
rect 188614 275312 188620 275324
rect 166500 275284 188620 275312
rect 166500 275272 166506 275284
rect 188614 275272 188620 275284
rect 188672 275272 188678 275324
rect 61746 274660 61752 274712
rect 61804 274700 61810 274712
rect 66806 274700 66812 274712
rect 61804 274672 66812 274700
rect 61804 274660 61810 274672
rect 66806 274660 66812 274672
rect 66864 274660 66870 274712
rect 162210 274660 162216 274712
rect 162268 274700 162274 274712
rect 169294 274700 169300 274712
rect 162268 274672 169300 274700
rect 162268 274660 162274 274672
rect 169294 274660 169300 274672
rect 169352 274660 169358 274712
rect 156506 274592 156512 274644
rect 156564 274632 156570 274644
rect 167730 274632 167736 274644
rect 156564 274604 167736 274632
rect 156564 274592 156570 274604
rect 167730 274592 167736 274604
rect 167788 274592 167794 274644
rect 264330 273980 264336 274032
rect 264388 274020 264394 274032
rect 280798 274020 280804 274032
rect 264388 273992 280804 274020
rect 264388 273980 264394 273992
rect 280798 273980 280804 273992
rect 280856 273980 280862 274032
rect 57698 273912 57704 273964
rect 57756 273952 57762 273964
rect 66898 273952 66904 273964
rect 57756 273924 66904 273952
rect 57756 273912 57762 273924
rect 66898 273912 66904 273924
rect 66956 273912 66962 273964
rect 159450 273912 159456 273964
rect 159508 273952 159514 273964
rect 187142 273952 187148 273964
rect 159508 273924 187148 273952
rect 159508 273912 159514 273924
rect 187142 273912 187148 273924
rect 187200 273912 187206 273964
rect 245838 273912 245844 273964
rect 245896 273952 245902 273964
rect 311894 273952 311900 273964
rect 245896 273924 311900 273952
rect 245896 273912 245902 273924
rect 311894 273912 311900 273924
rect 311952 273912 311958 273964
rect 62022 273232 62028 273284
rect 62080 273272 62086 273284
rect 66806 273272 66812 273284
rect 62080 273244 66812 273272
rect 62080 273232 62086 273244
rect 66806 273232 66812 273244
rect 66864 273232 66870 273284
rect 187050 273232 187056 273284
rect 187108 273272 187114 273284
rect 197354 273272 197360 273284
rect 187108 273244 197360 273272
rect 187108 273232 187114 273244
rect 197354 273232 197360 273244
rect 197412 273232 197418 273284
rect 245838 273232 245844 273284
rect 245896 273272 245902 273284
rect 249886 273272 249892 273284
rect 245896 273244 249892 273272
rect 245896 273232 245902 273244
rect 249886 273232 249892 273244
rect 249944 273232 249950 273284
rect 164970 272552 164976 272604
rect 165028 272592 165034 272604
rect 177482 272592 177488 272604
rect 165028 272564 177488 272592
rect 165028 272552 165034 272564
rect 177482 272552 177488 272564
rect 177540 272552 177546 272604
rect 165062 272484 165068 272536
rect 165120 272524 165126 272536
rect 197446 272524 197452 272536
rect 165120 272496 197452 272524
rect 165120 272484 165126 272496
rect 197446 272484 197452 272496
rect 197504 272484 197510 272536
rect 245746 272484 245752 272536
rect 245804 272524 245810 272536
rect 252646 272524 252652 272536
rect 245804 272496 252652 272524
rect 245804 272484 245810 272496
rect 252646 272484 252652 272496
rect 252704 272524 252710 272536
rect 253842 272524 253848 272536
rect 252704 272496 253848 272524
rect 252704 272484 252710 272496
rect 253842 272484 253848 272496
rect 253900 272484 253906 272536
rect 197354 271912 197360 271924
rect 183480 271884 197360 271912
rect 176102 271804 176108 271856
rect 176160 271844 176166 271856
rect 182910 271844 182916 271856
rect 176160 271816 182916 271844
rect 176160 271804 176166 271816
rect 182910 271804 182916 271816
rect 182968 271844 182974 271856
rect 183480 271844 183508 271884
rect 197354 271872 197360 271884
rect 197412 271872 197418 271924
rect 182968 271816 183508 271844
rect 182968 271804 182974 271816
rect 245838 271464 245844 271516
rect 245896 271504 245902 271516
rect 248598 271504 248604 271516
rect 245896 271476 248604 271504
rect 245896 271464 245902 271476
rect 248598 271464 248604 271476
rect 248656 271464 248662 271516
rect 157150 271124 157156 271176
rect 157208 271164 157214 271176
rect 191190 271164 191196 271176
rect 157208 271136 191196 271164
rect 157208 271124 157214 271136
rect 191190 271124 191196 271136
rect 191248 271124 191254 271176
rect 195514 270580 195520 270632
rect 195572 270620 195578 270632
rect 197814 270620 197820 270632
rect 195572 270592 197820 270620
rect 195572 270580 195578 270592
rect 197814 270580 197820 270592
rect 197872 270580 197878 270632
rect 48222 270512 48228 270564
rect 48280 270552 48286 270564
rect 66898 270552 66904 270564
rect 48280 270524 66904 270552
rect 48280 270512 48286 270524
rect 66898 270512 66904 270524
rect 66956 270512 66962 270564
rect 157242 270512 157248 270564
rect 157300 270552 157306 270564
rect 175918 270552 175924 270564
rect 157300 270524 175924 270552
rect 157300 270512 157306 270524
rect 175918 270512 175924 270524
rect 175976 270512 175982 270564
rect 186222 270512 186228 270564
rect 186280 270552 186286 270564
rect 197354 270552 197360 270564
rect 186280 270524 197360 270552
rect 186280 270512 186286 270524
rect 197354 270512 197360 270524
rect 197412 270512 197418 270564
rect 245930 270444 245936 270496
rect 245988 270484 245994 270496
rect 251174 270484 251180 270496
rect 245988 270456 251180 270484
rect 245988 270444 245994 270456
rect 251174 270444 251180 270456
rect 251232 270484 251238 270496
rect 252646 270484 252652 270496
rect 251232 270456 252652 270484
rect 251232 270444 251238 270456
rect 252646 270444 252652 270456
rect 252704 270444 252710 270496
rect 256878 270444 256884 270496
rect 256936 270484 256942 270496
rect 583386 270484 583392 270496
rect 256936 270456 583392 270484
rect 256936 270444 256942 270456
rect 583386 270444 583392 270456
rect 583444 270444 583450 270496
rect 194870 269832 194876 269884
rect 194928 269872 194934 269884
rect 197446 269872 197452 269884
rect 194928 269844 197452 269872
rect 194928 269832 194934 269844
rect 197446 269832 197452 269844
rect 197504 269832 197510 269884
rect 246574 269764 246580 269816
rect 246632 269804 246638 269816
rect 256878 269804 256884 269816
rect 246632 269776 256884 269804
rect 246632 269764 246638 269776
rect 256878 269764 256884 269776
rect 256936 269764 256942 269816
rect 181622 269152 181628 269204
rect 181680 269192 181686 269204
rect 197354 269192 197360 269204
rect 181680 269164 197360 269192
rect 181680 269152 181686 269164
rect 197354 269152 197360 269164
rect 197412 269152 197418 269204
rect 64506 269084 64512 269136
rect 64564 269124 64570 269136
rect 66714 269124 66720 269136
rect 64564 269096 66720 269124
rect 64564 269084 64570 269096
rect 66714 269084 66720 269096
rect 66772 269084 66778 269136
rect 157242 269084 157248 269136
rect 157300 269124 157306 269136
rect 195422 269124 195428 269136
rect 157300 269096 195428 269124
rect 157300 269084 157306 269096
rect 195422 269084 195428 269096
rect 195480 269084 195486 269136
rect 171962 269016 171968 269068
rect 172020 269056 172026 269068
rect 197354 269056 197360 269068
rect 172020 269028 197360 269056
rect 172020 269016 172026 269028
rect 197354 269016 197360 269028
rect 197412 269016 197418 269068
rect 245746 269016 245752 269068
rect 245804 269056 245810 269068
rect 263594 269056 263600 269068
rect 245804 269028 263600 269056
rect 245804 269016 245810 269028
rect 263594 269016 263600 269028
rect 263652 269016 263658 269068
rect 157242 268336 157248 268388
rect 157300 268376 157306 268388
rect 192570 268376 192576 268388
rect 157300 268348 192576 268376
rect 157300 268336 157306 268348
rect 192570 268336 192576 268348
rect 192628 268336 192634 268388
rect 263594 268336 263600 268388
rect 263652 268376 263658 268388
rect 582650 268376 582656 268388
rect 263652 268348 582656 268376
rect 263652 268336 263658 268348
rect 582650 268336 582656 268348
rect 582708 268336 582714 268388
rect 38654 267724 38660 267776
rect 38712 267764 38718 267776
rect 40678 267764 40684 267776
rect 38712 267736 40684 267764
rect 38712 267724 38718 267736
rect 40678 267724 40684 267736
rect 40736 267724 40742 267776
rect 157242 267656 157248 267708
rect 157300 267696 157306 267708
rect 195330 267696 195336 267708
rect 157300 267668 195336 267696
rect 157300 267656 157306 267668
rect 195330 267656 195336 267668
rect 195388 267656 195394 267708
rect 38654 267588 38660 267640
rect 38712 267628 38718 267640
rect 43438 267628 43444 267640
rect 38712 267600 43444 267628
rect 38712 267588 38718 267600
rect 43438 267588 43444 267600
rect 43496 267588 43502 267640
rect 3510 266976 3516 267028
rect 3568 267016 3574 267028
rect 38654 267016 38660 267028
rect 3568 266988 38660 267016
rect 3568 266976 3574 266988
rect 38654 266976 38660 266988
rect 38712 266976 38718 267028
rect 159634 266976 159640 267028
rect 159692 267016 159698 267028
rect 193950 267016 193956 267028
rect 159692 266988 193956 267016
rect 159692 266976 159698 266988
rect 193950 266976 193956 266988
rect 194008 266976 194014 267028
rect 246482 266976 246488 267028
rect 246540 267016 246546 267028
rect 294046 267016 294052 267028
rect 246540 266988 294052 267016
rect 246540 266976 246546 266988
rect 294046 266976 294052 266988
rect 294104 266976 294110 267028
rect 195882 266364 195888 266416
rect 195940 266404 195946 266416
rect 197998 266404 198004 266416
rect 195940 266376 198004 266404
rect 195940 266364 195946 266376
rect 197998 266364 198004 266376
rect 198056 266364 198062 266416
rect 245838 266364 245844 266416
rect 245896 266404 245902 266416
rect 276014 266404 276020 266416
rect 245896 266376 276020 266404
rect 245896 266364 245902 266376
rect 276014 266364 276020 266376
rect 276072 266364 276078 266416
rect 157242 266296 157248 266348
rect 157300 266336 157306 266348
rect 198090 266336 198096 266348
rect 157300 266308 198096 266336
rect 157300 266296 157306 266308
rect 198090 266296 198096 266308
rect 198148 266296 198154 266348
rect 245930 266296 245936 266348
rect 245988 266336 245994 266348
rect 267734 266336 267740 266348
rect 245988 266308 267740 266336
rect 245988 266296 245994 266308
rect 267734 266296 267740 266308
rect 267792 266336 267798 266348
rect 269022 266336 269028 266348
rect 267792 266308 269028 266336
rect 267792 266296 267798 266308
rect 269022 266296 269028 266308
rect 269080 266296 269086 266348
rect 191098 266228 191104 266280
rect 191156 266268 191162 266280
rect 197354 266268 197360 266280
rect 191156 266240 197360 266268
rect 191156 266228 191162 266240
rect 197354 266228 197360 266240
rect 197412 266228 197418 266280
rect 245930 265752 245936 265804
rect 245988 265792 245994 265804
rect 249978 265792 249984 265804
rect 245988 265764 249984 265792
rect 245988 265752 245994 265764
rect 249978 265752 249984 265764
rect 250036 265752 250042 265804
rect 269022 265616 269028 265668
rect 269080 265656 269086 265668
rect 583018 265656 583024 265668
rect 269080 265628 583024 265656
rect 269080 265616 269086 265628
rect 583018 265616 583024 265628
rect 583076 265616 583082 265668
rect 41322 264936 41328 264988
rect 41380 264976 41386 264988
rect 66806 264976 66812 264988
rect 41380 264948 66812 264976
rect 41380 264936 41386 264948
rect 66806 264936 66812 264948
rect 66864 264936 66870 264988
rect 50982 264188 50988 264240
rect 51040 264228 51046 264240
rect 65978 264228 65984 264240
rect 51040 264200 65984 264228
rect 51040 264188 51046 264200
rect 65978 264188 65984 264200
rect 66036 264228 66042 264240
rect 66530 264228 66536 264240
rect 66036 264200 66536 264228
rect 66036 264188 66042 264200
rect 66530 264188 66536 264200
rect 66588 264188 66594 264240
rect 156874 264188 156880 264240
rect 156932 264228 156938 264240
rect 174722 264228 174728 264240
rect 156932 264200 174728 264228
rect 156932 264188 156938 264200
rect 174722 264188 174728 264200
rect 174780 264188 174786 264240
rect 189902 264188 189908 264240
rect 189960 264228 189966 264240
rect 199562 264228 199568 264240
rect 189960 264200 199568 264228
rect 189960 264188 189966 264200
rect 199562 264188 199568 264200
rect 199620 264188 199626 264240
rect 246022 264188 246028 264240
rect 246080 264228 246086 264240
rect 296714 264228 296720 264240
rect 246080 264200 296720 264228
rect 246080 264188 246086 264200
rect 296714 264188 296720 264200
rect 296772 264188 296778 264240
rect 56318 263576 56324 263628
rect 56376 263616 56382 263628
rect 66806 263616 66812 263628
rect 56376 263588 66812 263616
rect 56376 263576 56382 263588
rect 66806 263576 66812 263588
rect 66864 263576 66870 263628
rect 164142 263576 164148 263628
rect 164200 263616 164206 263628
rect 197354 263616 197360 263628
rect 164200 263588 197360 263616
rect 164200 263576 164206 263588
rect 197354 263576 197360 263588
rect 197412 263576 197418 263628
rect 247126 263304 247132 263356
rect 247184 263304 247190 263356
rect 247034 263100 247040 263152
rect 247092 263140 247098 263152
rect 247144 263140 247172 263304
rect 247092 263112 247172 263140
rect 247092 263100 247098 263112
rect 52362 262828 52368 262880
rect 52420 262868 52426 262880
rect 63494 262868 63500 262880
rect 52420 262840 63500 262868
rect 52420 262828 52426 262840
rect 63494 262828 63500 262840
rect 63552 262828 63558 262880
rect 169294 262828 169300 262880
rect 169352 262868 169358 262880
rect 185670 262868 185676 262880
rect 169352 262840 185676 262868
rect 169352 262828 169358 262840
rect 185670 262828 185676 262840
rect 185728 262828 185734 262880
rect 246666 262828 246672 262880
rect 246724 262868 246730 262880
rect 310606 262868 310612 262880
rect 246724 262840 310612 262868
rect 246724 262828 246730 262840
rect 310606 262828 310612 262840
rect 310664 262828 310670 262880
rect 63494 262216 63500 262268
rect 63552 262256 63558 262268
rect 64598 262256 64604 262268
rect 63552 262228 64604 262256
rect 63552 262216 63558 262228
rect 64598 262216 64604 262228
rect 64656 262256 64662 262268
rect 66438 262256 66444 262268
rect 64656 262228 66444 262256
rect 64656 262216 64662 262228
rect 66438 262216 66444 262228
rect 66496 262216 66502 262268
rect 157242 262216 157248 262268
rect 157300 262256 157306 262268
rect 178770 262256 178776 262268
rect 157300 262228 178776 262256
rect 157300 262216 157306 262228
rect 178770 262216 178776 262228
rect 178828 262216 178834 262268
rect 185762 262216 185768 262268
rect 185820 262256 185826 262268
rect 197354 262256 197360 262268
rect 185820 262228 197360 262256
rect 185820 262216 185826 262228
rect 197354 262216 197360 262228
rect 197412 262216 197418 262268
rect 245930 262216 245936 262268
rect 245988 262256 245994 262268
rect 251450 262256 251456 262268
rect 245988 262228 251456 262256
rect 245988 262216 245994 262228
rect 251450 262216 251456 262228
rect 251508 262216 251514 262268
rect 160922 261536 160928 261588
rect 160980 261576 160986 261588
rect 169754 261576 169760 261588
rect 160980 261548 169760 261576
rect 160980 261536 160986 261548
rect 169754 261536 169760 261548
rect 169812 261536 169818 261588
rect 189902 261536 189908 261588
rect 189960 261576 189966 261588
rect 199378 261576 199384 261588
rect 189960 261548 199384 261576
rect 189960 261536 189966 261548
rect 199378 261536 199384 261548
rect 199436 261536 199442 261588
rect 29638 261468 29644 261520
rect 29696 261508 29702 261520
rect 52454 261508 52460 261520
rect 29696 261480 52460 261508
rect 29696 261468 29702 261480
rect 52454 261468 52460 261480
rect 52512 261468 52518 261520
rect 167730 261468 167736 261520
rect 167788 261508 167794 261520
rect 195514 261508 195520 261520
rect 167788 261480 195520 261508
rect 167788 261468 167794 261480
rect 195514 261468 195520 261480
rect 195572 261468 195578 261520
rect 246390 261468 246396 261520
rect 246448 261508 246454 261520
rect 247310 261508 247316 261520
rect 246448 261480 247316 261508
rect 246448 261468 246454 261480
rect 247310 261468 247316 261480
rect 247368 261508 247374 261520
rect 251174 261508 251180 261520
rect 247368 261480 251180 261508
rect 247368 261468 247374 261480
rect 251174 261468 251180 261480
rect 251232 261468 251238 261520
rect 251818 261468 251824 261520
rect 251876 261508 251882 261520
rect 281902 261508 281908 261520
rect 251876 261480 281908 261508
rect 251876 261468 251882 261480
rect 281902 261468 281908 261480
rect 281960 261468 281966 261520
rect 52454 260856 52460 260908
rect 52512 260896 52518 260908
rect 53466 260896 53472 260908
rect 52512 260868 53472 260896
rect 52512 260856 52518 260868
rect 53466 260856 53472 260868
rect 53524 260896 53530 260908
rect 66806 260896 66812 260908
rect 53524 260868 66812 260896
rect 53524 260856 53530 260868
rect 66806 260856 66812 260868
rect 66864 260856 66870 260908
rect 245930 260176 245936 260228
rect 245988 260216 245994 260228
rect 248690 260216 248696 260228
rect 245988 260188 248696 260216
rect 245988 260176 245994 260188
rect 248690 260176 248696 260188
rect 248748 260176 248754 260228
rect 160830 260108 160836 260160
rect 160888 260148 160894 260160
rect 171962 260148 171968 260160
rect 160888 260120 171968 260148
rect 160888 260108 160894 260120
rect 171962 260108 171968 260120
rect 172020 260108 172026 260160
rect 60550 259428 60556 259480
rect 60608 259468 60614 259480
rect 66806 259468 66812 259480
rect 60608 259440 66812 259468
rect 60608 259428 60614 259440
rect 66806 259428 66812 259440
rect 66864 259428 66870 259480
rect 188522 259428 188528 259480
rect 188580 259468 188586 259480
rect 197446 259468 197452 259480
rect 188580 259440 197452 259468
rect 188580 259428 188586 259440
rect 197446 259428 197452 259440
rect 197504 259428 197510 259480
rect 244366 259428 244372 259480
rect 244424 259468 244430 259480
rect 291194 259468 291200 259480
rect 244424 259440 291200 259468
rect 244424 259428 244430 259440
rect 291194 259428 291200 259440
rect 291252 259428 291258 259480
rect 184290 259360 184296 259412
rect 184348 259400 184354 259412
rect 197354 259400 197360 259412
rect 184348 259372 197360 259400
rect 184348 259360 184354 259372
rect 197354 259360 197360 259372
rect 197412 259360 197418 259412
rect 245930 259360 245936 259412
rect 245988 259400 245994 259412
rect 259546 259400 259552 259412
rect 245988 259372 259552 259400
rect 245988 259360 245994 259372
rect 259546 259360 259552 259372
rect 259604 259400 259610 259412
rect 260742 259400 260748 259412
rect 259604 259372 260748 259400
rect 259604 259360 259610 259372
rect 260742 259360 260748 259372
rect 260800 259360 260806 259412
rect 171870 258680 171876 258732
rect 171928 258720 171934 258732
rect 197906 258720 197912 258732
rect 171928 258692 197912 258720
rect 171928 258680 171934 258692
rect 197906 258680 197912 258692
rect 197964 258680 197970 258732
rect 260742 258680 260748 258732
rect 260800 258720 260806 258732
rect 300946 258720 300952 258732
rect 260800 258692 300952 258720
rect 260800 258680 260806 258692
rect 300946 258680 300952 258692
rect 301004 258680 301010 258732
rect 53742 258068 53748 258120
rect 53800 258108 53806 258120
rect 66714 258108 66720 258120
rect 53800 258080 66720 258108
rect 53800 258068 53806 258080
rect 66714 258068 66720 258080
rect 66772 258068 66778 258120
rect 156414 258068 156420 258120
rect 156472 258108 156478 258120
rect 170490 258108 170496 258120
rect 156472 258080 170496 258108
rect 156472 258068 156478 258080
rect 170490 258068 170496 258080
rect 170548 258068 170554 258120
rect 67450 258000 67456 258052
rect 67508 258040 67514 258052
rect 68186 258040 68192 258052
rect 67508 258012 68192 258040
rect 67508 258000 67514 258012
rect 68186 258000 68192 258012
rect 68244 258000 68250 258052
rect 156874 257932 156880 257984
rect 156932 257972 156938 257984
rect 159542 257972 159548 257984
rect 156932 257944 159548 257972
rect 156932 257932 156938 257944
rect 159542 257932 159548 257944
rect 159600 257932 159606 257984
rect 198642 257456 198648 257508
rect 198700 257496 198706 257508
rect 199378 257496 199384 257508
rect 198700 257468 199384 257496
rect 198700 257456 198706 257468
rect 199378 257456 199384 257468
rect 199436 257456 199442 257508
rect 195422 257388 195428 257440
rect 195480 257428 195486 257440
rect 200022 257428 200028 257440
rect 195480 257400 200028 257428
rect 195480 257388 195486 257400
rect 200022 257388 200028 257400
rect 200080 257388 200086 257440
rect 260190 257320 260196 257372
rect 260248 257360 260254 257372
rect 580350 257360 580356 257372
rect 260248 257332 580356 257360
rect 260248 257320 260254 257332
rect 580350 257320 580356 257332
rect 580408 257320 580414 257372
rect 157242 256776 157248 256828
rect 157300 256816 157306 256828
rect 177942 256816 177948 256828
rect 157300 256788 177948 256816
rect 157300 256776 157306 256788
rect 177942 256776 177948 256788
rect 178000 256816 178006 256828
rect 181438 256816 181444 256828
rect 178000 256788 181444 256816
rect 178000 256776 178006 256788
rect 181438 256776 181444 256788
rect 181496 256776 181502 256828
rect 197354 256816 197360 256828
rect 190426 256788 197360 256816
rect 158714 256708 158720 256760
rect 158772 256748 158778 256760
rect 184842 256748 184848 256760
rect 158772 256720 184848 256748
rect 158772 256708 158778 256720
rect 184842 256708 184848 256720
rect 184900 256748 184906 256760
rect 190426 256748 190454 256788
rect 197354 256776 197360 256788
rect 197412 256776 197418 256828
rect 184900 256720 190454 256748
rect 184900 256708 184906 256720
rect 188430 256640 188436 256692
rect 188488 256680 188494 256692
rect 197354 256680 197360 256692
rect 188488 256652 197360 256680
rect 188488 256640 188494 256652
rect 197354 256640 197360 256652
rect 197412 256640 197418 256692
rect 192570 256368 192576 256420
rect 192628 256408 192634 256420
rect 193858 256408 193864 256420
rect 192628 256380 193864 256408
rect 192628 256368 192634 256380
rect 193858 256368 193864 256380
rect 193916 256368 193922 256420
rect 245654 256028 245660 256080
rect 245712 256068 245718 256080
rect 260834 256068 260840 256080
rect 245712 256040 260840 256068
rect 245712 256028 245718 256040
rect 260834 256028 260840 256040
rect 260892 256028 260898 256080
rect 247126 255960 247132 256012
rect 247184 256000 247190 256012
rect 288434 256000 288440 256012
rect 247184 255972 288440 256000
rect 247184 255960 247190 255972
rect 288434 255960 288440 255972
rect 288492 255960 288498 256012
rect 60366 255688 60372 255740
rect 60424 255728 60430 255740
rect 66990 255728 66996 255740
rect 60424 255700 66996 255728
rect 60424 255688 60430 255700
rect 66990 255688 66996 255700
rect 67048 255688 67054 255740
rect 157242 255280 157248 255332
rect 157300 255320 157306 255332
rect 168374 255320 168380 255332
rect 157300 255292 168380 255320
rect 157300 255280 157306 255292
rect 168374 255280 168380 255292
rect 168432 255280 168438 255332
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 11698 255252 11704 255264
rect 3200 255224 11704 255252
rect 3200 255212 3206 255224
rect 11698 255212 11704 255224
rect 11756 255212 11762 255264
rect 178034 255212 178040 255264
rect 178092 255252 178098 255264
rect 195974 255252 195980 255264
rect 178092 255224 195980 255252
rect 178092 255212 178098 255224
rect 195974 255212 195980 255224
rect 196032 255212 196038 255264
rect 159542 254532 159548 254584
rect 159600 254572 159606 254584
rect 178034 254572 178040 254584
rect 159600 254544 178040 254572
rect 159600 254532 159606 254544
rect 178034 254532 178040 254544
rect 178092 254532 178098 254584
rect 260834 254532 260840 254584
rect 260892 254572 260898 254584
rect 295426 254572 295432 254584
rect 260892 254544 295432 254572
rect 260892 254532 260898 254544
rect 295426 254532 295432 254544
rect 295484 254532 295490 254584
rect 63126 253920 63132 253972
rect 63184 253960 63190 253972
rect 66898 253960 66904 253972
rect 63184 253932 66904 253960
rect 63184 253920 63190 253932
rect 66898 253920 66904 253932
rect 66956 253920 66962 253972
rect 157242 253920 157248 253972
rect 157300 253960 157306 253972
rect 179322 253960 179328 253972
rect 157300 253932 179328 253960
rect 157300 253920 157306 253932
rect 179322 253920 179328 253932
rect 179380 253920 179386 253972
rect 192662 253920 192668 253972
rect 192720 253960 192726 253972
rect 197354 253960 197360 253972
rect 192720 253932 197360 253960
rect 192720 253920 192726 253932
rect 197354 253920 197360 253932
rect 197412 253920 197418 253972
rect 245930 253852 245936 253904
rect 245988 253892 245994 253904
rect 258258 253892 258264 253904
rect 245988 253864 258264 253892
rect 245988 253852 245994 253864
rect 258258 253852 258264 253864
rect 258316 253892 258322 253904
rect 259362 253892 259368 253904
rect 258316 253864 259368 253892
rect 258316 253852 258322 253864
rect 259362 253852 259368 253864
rect 259420 253852 259426 253904
rect 156414 253580 156420 253632
rect 156472 253620 156478 253632
rect 158714 253620 158720 253632
rect 156472 253592 158720 253620
rect 156472 253580 156478 253592
rect 158714 253580 158720 253592
rect 158772 253580 158778 253632
rect 177482 253240 177488 253292
rect 177540 253280 177546 253292
rect 186314 253280 186320 253292
rect 177540 253252 186320 253280
rect 177540 253240 177546 253252
rect 186314 253240 186320 253252
rect 186372 253240 186378 253292
rect 158162 253172 158168 253224
rect 158220 253212 158226 253224
rect 165154 253212 165160 253224
rect 158220 253184 165160 253212
rect 158220 253172 158226 253184
rect 165154 253172 165160 253184
rect 165212 253172 165218 253224
rect 166534 253172 166540 253224
rect 166592 253212 166598 253224
rect 180334 253212 180340 253224
rect 166592 253184 180340 253212
rect 166592 253172 166598 253184
rect 180334 253172 180340 253184
rect 180392 253172 180398 253224
rect 245654 253172 245660 253224
rect 245712 253212 245718 253224
rect 256786 253212 256792 253224
rect 245712 253184 256792 253212
rect 245712 253172 245718 253184
rect 256786 253172 256792 253184
rect 256844 253172 256850 253224
rect 259362 253172 259368 253224
rect 259420 253212 259426 253224
rect 296806 253212 296812 253224
rect 259420 253184 296812 253212
rect 259420 253172 259426 253184
rect 296806 253172 296812 253184
rect 296864 253172 296870 253224
rect 186314 252628 186320 252680
rect 186372 252668 186378 252680
rect 187602 252668 187608 252680
rect 186372 252640 187608 252668
rect 186372 252628 186378 252640
rect 187602 252628 187608 252640
rect 187660 252668 187666 252680
rect 197446 252668 197452 252680
rect 187660 252640 197452 252668
rect 187660 252628 187666 252640
rect 197446 252628 197452 252640
rect 197504 252628 197510 252680
rect 55030 252560 55036 252612
rect 55088 252600 55094 252612
rect 57606 252600 57612 252612
rect 55088 252572 57612 252600
rect 55088 252560 55094 252572
rect 57606 252560 57612 252572
rect 57664 252600 57670 252612
rect 66898 252600 66904 252612
rect 57664 252572 66904 252600
rect 57664 252560 57670 252572
rect 66898 252560 66904 252572
rect 66956 252560 66962 252612
rect 179874 252560 179880 252612
rect 179932 252600 179938 252612
rect 197354 252600 197360 252612
rect 179932 252572 197360 252600
rect 179932 252560 179938 252572
rect 197354 252560 197360 252572
rect 197412 252560 197418 252612
rect 246022 252492 246028 252544
rect 246080 252532 246086 252544
rect 259454 252532 259460 252544
rect 246080 252504 259460 252532
rect 246080 252492 246086 252504
rect 259454 252492 259460 252504
rect 259512 252532 259518 252544
rect 260742 252532 260748 252544
rect 259512 252504 260748 252532
rect 259512 252492 259518 252504
rect 260742 252492 260748 252504
rect 260800 252492 260806 252544
rect 245930 252424 245936 252476
rect 245988 252464 245994 252476
rect 251358 252464 251364 252476
rect 245988 252436 251364 252464
rect 245988 252424 245994 252436
rect 251358 252424 251364 252436
rect 251416 252424 251422 252476
rect 58986 252084 58992 252136
rect 59044 252124 59050 252136
rect 66806 252124 66812 252136
rect 59044 252096 66812 252124
rect 59044 252084 59050 252096
rect 66806 252084 66812 252096
rect 66864 252084 66870 252136
rect 159358 251880 159364 251932
rect 159416 251920 159422 251932
rect 170398 251920 170404 251932
rect 159416 251892 170404 251920
rect 159416 251880 159422 251892
rect 170398 251880 170404 251892
rect 170456 251880 170462 251932
rect 168374 251812 168380 251864
rect 168432 251852 168438 251864
rect 195790 251852 195796 251864
rect 168432 251824 195796 251852
rect 168432 251812 168438 251824
rect 195790 251812 195796 251824
rect 195848 251852 195854 251864
rect 197446 251852 197452 251864
rect 195848 251824 197452 251852
rect 195848 251812 195854 251824
rect 197446 251812 197452 251824
rect 197504 251812 197510 251864
rect 260742 251812 260748 251864
rect 260800 251852 260806 251864
rect 583662 251852 583668 251864
rect 260800 251824 583668 251852
rect 260800 251812 260806 251824
rect 583662 251812 583668 251824
rect 583720 251812 583726 251864
rect 156874 251336 156880 251388
rect 156932 251376 156938 251388
rect 162210 251376 162216 251388
rect 156932 251348 162216 251376
rect 156932 251336 156938 251348
rect 162210 251336 162216 251348
rect 162268 251336 162274 251388
rect 191098 251200 191104 251252
rect 191156 251240 191162 251252
rect 197354 251240 197360 251252
rect 191156 251212 197360 251240
rect 191156 251200 191162 251212
rect 197354 251200 197360 251212
rect 197412 251200 197418 251252
rect 245654 250452 245660 250504
rect 245712 250492 245718 250504
rect 252738 250492 252744 250504
rect 245712 250464 252744 250492
rect 245712 250452 245718 250464
rect 252738 250452 252744 250464
rect 252796 250492 252802 250504
rect 253014 250492 253020 250504
rect 252796 250464 253020 250492
rect 252796 250452 252802 250464
rect 253014 250452 253020 250464
rect 253072 250452 253078 250504
rect 256786 250452 256792 250504
rect 256844 250492 256850 250504
rect 287054 250492 287060 250504
rect 256844 250464 287060 250492
rect 256844 250452 256850 250464
rect 287054 250452 287060 250464
rect 287112 250452 287118 250504
rect 164142 249840 164148 249892
rect 164200 249880 164206 249892
rect 169018 249880 169024 249892
rect 164200 249852 169024 249880
rect 164200 249840 164206 249852
rect 169018 249840 169024 249852
rect 169076 249840 169082 249892
rect 185670 249840 185676 249892
rect 185728 249880 185734 249892
rect 197354 249880 197360 249892
rect 185728 249852 197360 249880
rect 185728 249840 185734 249852
rect 197354 249840 197360 249852
rect 197412 249840 197418 249892
rect 157242 249772 157248 249824
rect 157300 249812 157306 249824
rect 196342 249812 196348 249824
rect 157300 249784 196348 249812
rect 157300 249772 157306 249784
rect 196342 249772 196348 249784
rect 196400 249772 196406 249824
rect 157150 249704 157156 249756
rect 157208 249744 157214 249756
rect 164142 249744 164148 249756
rect 157208 249716 164148 249744
rect 157208 249704 157214 249716
rect 164142 249704 164148 249716
rect 164200 249704 164206 249756
rect 167822 249704 167828 249756
rect 167880 249744 167886 249756
rect 169202 249744 169208 249756
rect 167880 249716 169208 249744
rect 167880 249704 167886 249716
rect 169202 249704 169208 249716
rect 169260 249704 169266 249756
rect 191190 249704 191196 249756
rect 191248 249744 191254 249756
rect 195698 249744 195704 249756
rect 191248 249716 195704 249744
rect 191248 249704 191254 249716
rect 195698 249704 195704 249716
rect 195756 249744 195762 249756
rect 197354 249744 197360 249756
rect 195756 249716 197360 249744
rect 195756 249704 195762 249716
rect 197354 249704 197360 249716
rect 197412 249704 197418 249756
rect 178862 249296 178868 249348
rect 178920 249336 178926 249348
rect 179874 249336 179880 249348
rect 178920 249308 179880 249336
rect 178920 249296 178926 249308
rect 179874 249296 179880 249308
rect 179932 249296 179938 249348
rect 169754 249024 169760 249076
rect 169812 249064 169818 249076
rect 199470 249064 199476 249076
rect 169812 249036 199476 249064
rect 169812 249024 169818 249036
rect 199470 249024 199476 249036
rect 199528 249024 199534 249076
rect 253014 249024 253020 249076
rect 253072 249064 253078 249076
rect 285674 249064 285680 249076
rect 253072 249036 285680 249064
rect 253072 249024 253078 249036
rect 285674 249024 285680 249036
rect 285732 249024 285738 249076
rect 61930 248412 61936 248464
rect 61988 248452 61994 248464
rect 66806 248452 66812 248464
rect 61988 248424 66812 248452
rect 61988 248412 61994 248424
rect 66806 248412 66812 248424
rect 66864 248412 66870 248464
rect 156414 248412 156420 248464
rect 156472 248452 156478 248464
rect 177850 248452 177856 248464
rect 156472 248424 177856 248452
rect 156472 248412 156478 248424
rect 177850 248412 177856 248424
rect 177908 248412 177914 248464
rect 67450 248276 67456 248328
rect 67508 248316 67514 248328
rect 67910 248316 67916 248328
rect 67508 248288 67916 248316
rect 67508 248276 67514 248288
rect 67910 248276 67916 248288
rect 67968 248276 67974 248328
rect 171778 247732 171784 247784
rect 171836 247772 171842 247784
rect 194410 247772 194416 247784
rect 171836 247744 194416 247772
rect 171836 247732 171842 247744
rect 194410 247732 194416 247744
rect 194468 247732 194474 247784
rect 158622 247664 158628 247716
rect 158680 247704 158686 247716
rect 182726 247704 182732 247716
rect 158680 247676 182732 247704
rect 158680 247664 158686 247676
rect 182726 247664 182732 247676
rect 182784 247664 182790 247716
rect 245930 247664 245936 247716
rect 245988 247704 245994 247716
rect 248690 247704 248696 247716
rect 245988 247676 248696 247704
rect 245988 247664 245994 247676
rect 248690 247664 248696 247676
rect 248748 247704 248754 247716
rect 582834 247704 582840 247716
rect 248748 247676 582840 247704
rect 248748 247664 248754 247676
rect 582834 247664 582840 247676
rect 582892 247664 582898 247716
rect 50982 247052 50988 247104
rect 51040 247092 51046 247104
rect 66622 247092 66628 247104
rect 51040 247064 66628 247092
rect 51040 247052 51046 247064
rect 66622 247052 66628 247064
rect 66680 247052 66686 247104
rect 191190 247052 191196 247104
rect 191248 247092 191254 247104
rect 197446 247092 197452 247104
rect 191248 247064 197452 247092
rect 191248 247052 191254 247064
rect 197446 247052 197452 247064
rect 197504 247052 197510 247104
rect 195238 246984 195244 247036
rect 195296 247024 195302 247036
rect 197354 247024 197360 247036
rect 195296 246996 197360 247024
rect 195296 246984 195302 246996
rect 197354 246984 197360 246996
rect 197412 246984 197418 247036
rect 245930 246372 245936 246424
rect 245988 246412 245994 246424
rect 254026 246412 254032 246424
rect 245988 246384 254032 246412
rect 245988 246372 245994 246384
rect 254026 246372 254032 246384
rect 254084 246372 254090 246424
rect 245010 246304 245016 246356
rect 245068 246344 245074 246356
rect 306558 246344 306564 246356
rect 245068 246316 306564 246344
rect 245068 246304 245074 246316
rect 306558 246304 306564 246316
rect 306616 246304 306622 246356
rect 194502 246032 194508 246084
rect 194560 246072 194566 246084
rect 195330 246072 195336 246084
rect 194560 246044 195336 246072
rect 194560 246032 194566 246044
rect 195330 246032 195336 246044
rect 195388 246032 195394 246084
rect 156782 245692 156788 245744
rect 156840 245732 156846 245744
rect 185762 245732 185768 245744
rect 156840 245704 185768 245732
rect 156840 245692 156846 245704
rect 185762 245692 185768 245704
rect 185820 245692 185826 245744
rect 154850 245624 154856 245676
rect 154908 245664 154914 245676
rect 187050 245664 187056 245676
rect 154908 245636 187056 245664
rect 154908 245624 154914 245636
rect 187050 245624 187056 245636
rect 187108 245624 187114 245676
rect 254026 245624 254032 245676
rect 254084 245664 254090 245676
rect 254578 245664 254584 245676
rect 254084 245636 254584 245664
rect 254084 245624 254090 245636
rect 254578 245624 254584 245636
rect 254636 245624 254642 245676
rect 53558 245556 53564 245608
rect 53616 245596 53622 245608
rect 66622 245596 66628 245608
rect 53616 245568 66628 245596
rect 53616 245556 53622 245568
rect 66622 245556 66628 245568
rect 66680 245556 66686 245608
rect 190362 245420 190368 245472
rect 190420 245460 190426 245472
rect 191834 245460 191840 245472
rect 190420 245432 191840 245460
rect 190420 245420 190426 245432
rect 191834 245420 191840 245432
rect 191892 245420 191898 245472
rect 194410 245148 194416 245200
rect 194468 245188 194474 245200
rect 197354 245188 197360 245200
rect 194468 245160 197360 245188
rect 194468 245148 194474 245160
rect 197354 245148 197360 245160
rect 197412 245148 197418 245200
rect 196342 245012 196348 245064
rect 196400 245052 196406 245064
rect 198734 245052 198740 245064
rect 196400 245024 198740 245052
rect 196400 245012 196406 245024
rect 198734 245012 198740 245024
rect 198792 245012 198798 245064
rect 177850 244876 177856 244928
rect 177908 244916 177914 244928
rect 189994 244916 190000 244928
rect 177908 244888 190000 244916
rect 177908 244876 177914 244888
rect 189994 244876 190000 244888
rect 190052 244876 190058 244928
rect 280890 244876 280896 244928
rect 280948 244916 280954 244928
rect 310514 244916 310520 244928
rect 280948 244888 310520 244916
rect 280948 244876 280954 244888
rect 310514 244876 310520 244888
rect 310572 244876 310578 244928
rect 155310 244332 155316 244384
rect 155368 244372 155374 244384
rect 155368 244344 161474 244372
rect 155368 244332 155374 244344
rect 156966 244264 156972 244316
rect 157024 244304 157030 244316
rect 160830 244304 160836 244316
rect 157024 244276 160836 244304
rect 157024 244264 157030 244276
rect 160830 244264 160836 244276
rect 160888 244264 160894 244316
rect 161446 244304 161474 244344
rect 192570 244304 192576 244316
rect 161446 244276 192576 244304
rect 192570 244264 192576 244276
rect 192628 244304 192634 244316
rect 192754 244304 192760 244316
rect 192628 244276 192760 244304
rect 192628 244264 192634 244276
rect 192754 244264 192760 244276
rect 192812 244264 192818 244316
rect 155402 243380 155408 243432
rect 155460 243420 155466 243432
rect 155862 243420 155868 243432
rect 155460 243392 155868 243420
rect 155460 243380 155466 243392
rect 155862 243380 155868 243392
rect 155920 243380 155926 243432
rect 155862 242972 155868 243024
rect 155920 243012 155926 243024
rect 174630 243012 174636 243024
rect 155920 242984 174636 243012
rect 155920 242972 155926 242984
rect 174630 242972 174636 242984
rect 174688 242972 174694 243024
rect 156046 242904 156052 242956
rect 156104 242944 156110 242956
rect 188430 242944 188436 242956
rect 156104 242916 188436 242944
rect 156104 242904 156110 242916
rect 188430 242904 188436 242916
rect 188488 242904 188494 242956
rect 245930 242904 245936 242956
rect 245988 242944 245994 242956
rect 271322 242944 271328 242956
rect 245988 242916 271328 242944
rect 245988 242904 245994 242916
rect 271322 242904 271328 242916
rect 271380 242904 271386 242956
rect 265618 242224 265624 242276
rect 265676 242264 265682 242276
rect 278866 242264 278872 242276
rect 265676 242236 278872 242264
rect 265676 242224 265682 242236
rect 278866 242224 278872 242236
rect 278924 242224 278930 242276
rect 169754 242196 169760 242208
rect 151786 242168 169760 242196
rect 67450 242020 67456 242072
rect 67508 242060 67514 242072
rect 73890 242060 73896 242072
rect 67508 242032 73896 242060
rect 67508 242020 67514 242032
rect 73890 242020 73896 242032
rect 73948 242020 73954 242072
rect 150066 242020 150072 242072
rect 150124 242060 150130 242072
rect 151786 242060 151814 242168
rect 169754 242156 169760 242168
rect 169812 242156 169818 242208
rect 173802 242156 173808 242208
rect 173860 242196 173866 242208
rect 197354 242196 197360 242208
rect 173860 242168 197360 242196
rect 173860 242156 173866 242168
rect 197354 242156 197360 242168
rect 197412 242156 197418 242208
rect 271230 242156 271236 242208
rect 271288 242196 271294 242208
rect 298278 242196 298284 242208
rect 271288 242168 298284 242196
rect 271288 242156 271294 242168
rect 298278 242156 298284 242168
rect 298336 242156 298342 242208
rect 150124 242032 151814 242060
rect 150124 242020 150130 242032
rect 70302 241884 70308 241936
rect 70360 241924 70366 241936
rect 76374 241924 76380 241936
rect 70360 241896 76380 241924
rect 70360 241884 70366 241896
rect 76374 241884 76380 241896
rect 76432 241884 76438 241936
rect 192754 241516 192760 241528
rect 151786 241488 192760 241516
rect 3510 241408 3516 241460
rect 3568 241448 3574 241460
rect 36538 241448 36544 241460
rect 3568 241420 36544 241448
rect 3568 241408 3574 241420
rect 36538 241408 36544 241420
rect 36596 241408 36602 241460
rect 43438 241408 43444 241460
rect 43496 241448 43502 241460
rect 92888 241448 92894 241460
rect 43496 241420 92894 241448
rect 43496 241408 43502 241420
rect 92888 241408 92894 241420
rect 92946 241408 92952 241460
rect 144224 241408 144230 241460
rect 144282 241448 144288 241460
rect 151786 241448 151814 241488
rect 192754 241476 192760 241488
rect 192812 241476 192818 241528
rect 246390 241476 246396 241528
rect 246448 241516 246454 241528
rect 247218 241516 247224 241528
rect 246448 241488 247224 241516
rect 246448 241476 246454 241488
rect 247218 241476 247224 241488
rect 247276 241516 247282 241528
rect 268378 241516 268384 241528
rect 247276 241488 268384 241516
rect 247276 241476 247282 241488
rect 268378 241476 268384 241488
rect 268436 241476 268442 241528
rect 144282 241420 151814 241448
rect 144282 241408 144288 241420
rect 106090 240796 106096 240848
rect 106148 240836 106154 240848
rect 124858 240836 124864 240848
rect 106148 240808 124864 240836
rect 106148 240796 106154 240808
rect 124858 240796 124864 240808
rect 124916 240796 124922 240848
rect 152458 240796 152464 240848
rect 152516 240836 152522 240848
rect 162302 240836 162308 240848
rect 152516 240808 162308 240836
rect 152516 240796 152522 240808
rect 162302 240796 162308 240808
rect 162360 240796 162366 240848
rect 67542 240728 67548 240780
rect 67600 240768 67606 240780
rect 74718 240768 74724 240780
rect 67600 240740 74724 240768
rect 67600 240728 67606 240740
rect 74718 240728 74724 240740
rect 74776 240728 74782 240780
rect 82538 240728 82544 240780
rect 82596 240768 82602 240780
rect 116578 240768 116584 240780
rect 82596 240740 116584 240768
rect 82596 240728 82602 240740
rect 116578 240728 116584 240740
rect 116636 240728 116642 240780
rect 138842 240728 138848 240780
rect 138900 240768 138906 240780
rect 147674 240768 147680 240780
rect 138900 240740 147680 240768
rect 138900 240728 138906 240740
rect 147674 240728 147680 240740
rect 147732 240728 147738 240780
rect 149514 240728 149520 240780
rect 149572 240768 149578 240780
rect 149572 240740 209774 240768
rect 149572 240728 149578 240740
rect 195698 240456 195704 240508
rect 195756 240496 195762 240508
rect 200114 240496 200120 240508
rect 195756 240468 200120 240496
rect 195756 240456 195762 240468
rect 200114 240456 200120 240468
rect 200172 240456 200178 240508
rect 69014 240116 69020 240168
rect 69072 240156 69078 240168
rect 69750 240156 69756 240168
rect 69072 240128 69756 240156
rect 69072 240116 69078 240128
rect 69750 240116 69756 240128
rect 69808 240116 69814 240168
rect 115934 240116 115940 240168
rect 115992 240156 115998 240168
rect 116854 240156 116860 240168
rect 115992 240128 116860 240156
rect 115992 240116 115998 240128
rect 116854 240116 116860 240128
rect 116912 240116 116918 240168
rect 120718 240116 120724 240168
rect 120776 240156 120782 240168
rect 136082 240156 136088 240168
rect 120776 240128 136088 240156
rect 120776 240116 120782 240128
rect 136082 240116 136088 240128
rect 136140 240116 136146 240168
rect 198642 240116 198648 240168
rect 198700 240156 198706 240168
rect 200298 240156 200304 240168
rect 198700 240128 200304 240156
rect 198700 240116 198706 240128
rect 200298 240116 200304 240128
rect 200356 240116 200362 240168
rect 209746 240156 209774 240740
rect 218146 240156 218152 240168
rect 209746 240128 218152 240156
rect 218146 240116 218152 240128
rect 218204 240116 218210 240168
rect 224954 240116 224960 240168
rect 225012 240156 225018 240168
rect 227806 240156 227812 240168
rect 225012 240128 227812 240156
rect 225012 240116 225018 240128
rect 227806 240116 227812 240128
rect 227864 240116 227870 240168
rect 242802 240116 242808 240168
rect 242860 240156 242866 240168
rect 302326 240156 302332 240168
rect 242860 240128 302332 240156
rect 242860 240116 242866 240128
rect 302326 240116 302332 240128
rect 302384 240116 302390 240168
rect 68922 240048 68928 240100
rect 68980 240088 68986 240100
rect 71406 240088 71412 240100
rect 68980 240060 71412 240088
rect 68980 240048 68986 240060
rect 71406 240048 71412 240060
rect 71464 240048 71470 240100
rect 76558 240048 76564 240100
rect 76616 240088 76622 240100
rect 77294 240088 77300 240100
rect 76616 240060 77300 240088
rect 76616 240048 76622 240060
rect 77294 240048 77300 240060
rect 77352 240048 77358 240100
rect 86034 240048 86040 240100
rect 86092 240088 86098 240100
rect 86862 240088 86868 240100
rect 86092 240060 86868 240088
rect 86092 240048 86098 240060
rect 86862 240048 86868 240060
rect 86920 240048 86926 240100
rect 90450 240048 90456 240100
rect 90508 240088 90514 240100
rect 90910 240088 90916 240100
rect 90508 240060 90916 240088
rect 90508 240048 90514 240060
rect 90910 240048 90916 240060
rect 90968 240048 90974 240100
rect 91922 240048 91928 240100
rect 91980 240088 91986 240100
rect 92382 240088 92388 240100
rect 91980 240060 92388 240088
rect 91980 240048 91986 240060
rect 92382 240048 92388 240060
rect 92440 240048 92446 240100
rect 99374 240048 99380 240100
rect 99432 240088 99438 240100
rect 100662 240088 100668 240100
rect 99432 240060 100668 240088
rect 99432 240048 99438 240060
rect 100662 240048 100668 240060
rect 100720 240048 100726 240100
rect 115290 240048 115296 240100
rect 115348 240088 115354 240100
rect 115842 240088 115848 240100
rect 115348 240060 115848 240088
rect 115348 240048 115354 240060
rect 115842 240048 115848 240060
rect 115900 240048 115906 240100
rect 120442 240048 120448 240100
rect 120500 240088 120506 240100
rect 121362 240088 121368 240100
rect 120500 240060 121368 240088
rect 120500 240048 120506 240060
rect 121362 240048 121368 240060
rect 121420 240048 121426 240100
rect 121730 240048 121736 240100
rect 121788 240088 121794 240100
rect 122742 240088 122748 240100
rect 121788 240060 122748 240088
rect 121788 240048 121794 240060
rect 122742 240048 122748 240060
rect 122800 240048 122806 240100
rect 124674 240048 124680 240100
rect 124732 240088 124738 240100
rect 125410 240088 125416 240100
rect 124732 240060 125416 240088
rect 124732 240048 124738 240060
rect 125410 240048 125416 240060
rect 125468 240048 125474 240100
rect 126974 240048 126980 240100
rect 127032 240088 127038 240100
rect 127526 240088 127532 240100
rect 127032 240060 127532 240088
rect 127032 240048 127038 240060
rect 127526 240048 127532 240060
rect 127584 240048 127590 240100
rect 130378 240048 130384 240100
rect 130436 240088 130442 240100
rect 130930 240088 130936 240100
rect 130436 240060 130936 240088
rect 130436 240048 130442 240060
rect 130930 240048 130936 240060
rect 130988 240048 130994 240100
rect 131850 240048 131856 240100
rect 131908 240088 131914 240100
rect 132402 240088 132408 240100
rect 131908 240060 132408 240088
rect 131908 240048 131914 240060
rect 132402 240048 132408 240060
rect 132460 240048 132466 240100
rect 134610 240048 134616 240100
rect 134668 240088 134674 240100
rect 135162 240088 135168 240100
rect 134668 240060 135168 240088
rect 134668 240048 134674 240060
rect 135162 240048 135168 240060
rect 135220 240048 135226 240100
rect 138014 240048 138020 240100
rect 138072 240088 138078 240100
rect 138934 240088 138940 240100
rect 138072 240060 138940 240088
rect 138072 240048 138078 240060
rect 138934 240048 138940 240060
rect 138992 240048 138998 240100
rect 143994 240048 144000 240100
rect 144052 240088 144058 240100
rect 144822 240088 144828 240100
rect 144052 240060 144828 240088
rect 144052 240048 144058 240060
rect 144822 240048 144828 240060
rect 144880 240048 144886 240100
rect 147674 240048 147680 240100
rect 147732 240088 147738 240100
rect 165062 240088 165068 240100
rect 147732 240060 165068 240088
rect 147732 240048 147738 240060
rect 165062 240048 165068 240060
rect 165120 240048 165126 240100
rect 242250 240048 242256 240100
rect 242308 240088 242314 240100
rect 245654 240088 245660 240100
rect 242308 240060 245660 240088
rect 242308 240048 242314 240060
rect 245654 240048 245660 240060
rect 245712 240048 245718 240100
rect 74810 239980 74816 240032
rect 74868 240020 74874 240032
rect 83458 240020 83464 240032
rect 74868 239992 83464 240020
rect 74868 239980 74874 239992
rect 83458 239980 83464 239992
rect 83516 239980 83522 240032
rect 127434 239980 127440 240032
rect 127492 240020 127498 240032
rect 128262 240020 128268 240032
rect 127492 239992 128268 240020
rect 127492 239980 127498 239992
rect 128262 239980 128268 239992
rect 128320 239980 128326 240032
rect 106826 239912 106832 239964
rect 106884 239952 106890 239964
rect 107562 239952 107568 239964
rect 106884 239924 107568 239952
rect 106884 239912 106890 239924
rect 107562 239912 107568 239924
rect 107620 239912 107626 239964
rect 111058 239912 111064 239964
rect 111116 239952 111122 239964
rect 111610 239952 111616 239964
rect 111116 239924 111616 239952
rect 111116 239912 111122 239924
rect 111610 239912 111616 239924
rect 111668 239912 111674 239964
rect 120994 239912 121000 239964
rect 121052 239952 121058 239964
rect 122926 239952 122932 239964
rect 121052 239924 122932 239952
rect 121052 239912 121058 239924
rect 122926 239912 122932 239924
rect 122984 239912 122990 239964
rect 133138 239912 133144 239964
rect 133196 239952 133202 239964
rect 133782 239952 133788 239964
rect 133196 239924 133788 239952
rect 133196 239912 133202 239924
rect 133782 239912 133788 239924
rect 133840 239912 133846 239964
rect 142246 239912 142252 239964
rect 142304 239952 142310 239964
rect 143442 239952 143448 239964
rect 142304 239924 143448 239952
rect 142304 239912 142310 239924
rect 143442 239912 143448 239924
rect 143500 239912 143506 239964
rect 88978 239776 88984 239828
rect 89036 239816 89042 239828
rect 89622 239816 89628 239828
rect 89036 239788 89628 239816
rect 89036 239776 89042 239788
rect 89622 239776 89628 239788
rect 89680 239776 89686 239828
rect 148226 239776 148232 239828
rect 148284 239816 148290 239828
rect 148962 239816 148968 239828
rect 148284 239788 148968 239816
rect 148284 239776 148290 239788
rect 148962 239776 148968 239788
rect 149020 239776 149026 239828
rect 71682 239640 71688 239692
rect 71740 239680 71746 239692
rect 73798 239680 73804 239692
rect 71740 239652 73804 239680
rect 71740 239640 71746 239652
rect 73798 239640 73804 239652
rect 73856 239640 73862 239692
rect 75362 239640 75368 239692
rect 75420 239680 75426 239692
rect 75822 239680 75828 239692
rect 75420 239652 75828 239680
rect 75420 239640 75426 239652
rect 75822 239640 75828 239652
rect 75880 239640 75886 239692
rect 101122 239640 101128 239692
rect 101180 239680 101186 239692
rect 102042 239680 102048 239692
rect 101180 239652 102048 239680
rect 101180 239640 101186 239652
rect 102042 239640 102048 239652
rect 102100 239640 102106 239692
rect 149054 239572 149060 239624
rect 149112 239612 149118 239624
rect 149606 239612 149612 239624
rect 149112 239584 149612 239612
rect 149112 239572 149118 239584
rect 149606 239572 149612 239584
rect 149664 239572 149670 239624
rect 79042 239504 79048 239556
rect 79100 239544 79106 239556
rect 79962 239544 79968 239556
rect 79100 239516 79968 239544
rect 79100 239504 79106 239516
rect 79962 239504 79968 239516
rect 80020 239504 80026 239556
rect 141050 239504 141056 239556
rect 141108 239544 141114 239556
rect 142062 239544 142068 239556
rect 141108 239516 142068 239544
rect 141108 239504 141114 239516
rect 142062 239504 142068 239516
rect 142120 239504 142126 239556
rect 200114 239504 200120 239556
rect 200172 239544 200178 239556
rect 236730 239544 236736 239556
rect 200172 239516 236736 239544
rect 200172 239504 200178 239516
rect 236730 239504 236736 239516
rect 236788 239504 236794 239556
rect 198734 239436 198740 239488
rect 198792 239476 198798 239488
rect 238754 239476 238760 239488
rect 198792 239448 238760 239476
rect 198792 239436 198798 239448
rect 238754 239436 238760 239448
rect 238812 239436 238818 239488
rect 81802 239368 81808 239420
rect 81860 239408 81866 239420
rect 82722 239408 82728 239420
rect 81860 239380 82728 239408
rect 81860 239368 81866 239380
rect 82722 239368 82728 239380
rect 82780 239368 82786 239420
rect 84746 239368 84752 239420
rect 84804 239408 84810 239420
rect 200114 239408 200120 239420
rect 84804 239380 200120 239408
rect 84804 239368 84810 239380
rect 200114 239368 200120 239380
rect 200172 239368 200178 239420
rect 80514 239232 80520 239284
rect 80572 239272 80578 239284
rect 81250 239272 81256 239284
rect 80572 239244 81256 239272
rect 80572 239232 80578 239244
rect 81250 239232 81256 239244
rect 81308 239232 81314 239284
rect 109586 239232 109592 239284
rect 109644 239272 109650 239284
rect 110322 239272 110328 239284
rect 109644 239244 110328 239272
rect 109644 239232 109650 239244
rect 110322 239232 110328 239244
rect 110380 239232 110386 239284
rect 128906 239232 128912 239284
rect 128964 239272 128970 239284
rect 129642 239272 129648 239284
rect 128964 239244 129648 239272
rect 128964 239232 128970 239244
rect 129642 239232 129648 239244
rect 129700 239232 129706 239284
rect 153930 239232 153936 239284
rect 153988 239272 153994 239284
rect 154482 239272 154488 239284
rect 153988 239244 154488 239272
rect 153988 239232 153994 239244
rect 154482 239232 154488 239244
rect 154540 239232 154546 239284
rect 69474 238824 69480 238876
rect 69532 238864 69538 238876
rect 75270 238864 75276 238876
rect 69532 238836 75276 238864
rect 69532 238824 69538 238836
rect 75270 238824 75276 238836
rect 75328 238824 75334 238876
rect 240134 238756 240140 238808
rect 240192 238796 240198 238808
rect 241238 238796 241244 238808
rect 240192 238768 241244 238796
rect 240192 238756 240198 238768
rect 241238 238756 241244 238768
rect 241296 238796 241302 238808
rect 257430 238796 257436 238808
rect 241296 238768 257436 238796
rect 241296 238756 241302 238768
rect 257430 238756 257436 238768
rect 257488 238756 257494 238808
rect 96614 238688 96620 238740
rect 96672 238728 96678 238740
rect 214190 238728 214196 238740
rect 96672 238700 214196 238728
rect 96672 238688 96678 238700
rect 214190 238688 214196 238700
rect 214248 238688 214254 238740
rect 218146 238688 218152 238740
rect 218204 238728 218210 238740
rect 240318 238728 240324 238740
rect 218204 238700 240324 238728
rect 218204 238688 218210 238700
rect 240318 238688 240324 238700
rect 240376 238688 240382 238740
rect 241790 238688 241796 238740
rect 241848 238728 241854 238740
rect 258166 238728 258172 238740
rect 241848 238700 258172 238728
rect 241848 238688 241854 238700
rect 258166 238688 258172 238700
rect 258224 238688 258230 238740
rect 107654 238620 107660 238672
rect 107712 238660 107718 238672
rect 219894 238660 219900 238672
rect 107712 238632 219900 238660
rect 107712 238620 107718 238632
rect 219894 238620 219900 238632
rect 219952 238620 219958 238672
rect 221090 238620 221096 238672
rect 221148 238660 221154 238672
rect 227622 238660 227628 238672
rect 221148 238632 227628 238660
rect 221148 238620 221154 238632
rect 227622 238620 227628 238632
rect 227680 238620 227686 238672
rect 238754 238620 238760 238672
rect 238812 238660 238818 238672
rect 243906 238660 243912 238672
rect 238812 238632 243912 238660
rect 238812 238620 238818 238632
rect 243906 238620 243912 238632
rect 243964 238620 243970 238672
rect 231118 238552 231124 238604
rect 231176 238592 231182 238604
rect 234706 238592 234712 238604
rect 231176 238564 234712 238592
rect 231176 238552 231182 238564
rect 234706 238552 234712 238564
rect 234764 238552 234770 238604
rect 229094 238076 229100 238128
rect 229152 238116 229158 238128
rect 230474 238116 230480 238128
rect 229152 238088 230480 238116
rect 229152 238076 229158 238088
rect 230474 238076 230480 238088
rect 230532 238076 230538 238128
rect 61746 238008 61752 238060
rect 61804 238048 61810 238060
rect 108298 238048 108304 238060
rect 61804 238020 108304 238048
rect 61804 238008 61810 238020
rect 108298 238008 108304 238020
rect 108356 238008 108362 238060
rect 241790 237804 241796 237856
rect 241848 237844 241854 237856
rect 242434 237844 242440 237856
rect 241848 237816 242440 237844
rect 241848 237804 241854 237816
rect 242434 237804 242440 237816
rect 242492 237804 242498 237856
rect 65886 237532 65892 237584
rect 65944 237572 65950 237584
rect 72510 237572 72516 237584
rect 65944 237544 72516 237572
rect 65944 237532 65950 237544
rect 72510 237532 72516 237544
rect 72568 237532 72574 237584
rect 214190 237464 214196 237516
rect 214248 237504 214254 237516
rect 214650 237504 214656 237516
rect 214248 237476 214656 237504
rect 214248 237464 214254 237476
rect 214650 237464 214656 237476
rect 214708 237464 214714 237516
rect 214558 237396 214564 237448
rect 214616 237436 214622 237448
rect 216030 237436 216036 237448
rect 214616 237408 216036 237436
rect 214616 237396 214622 237408
rect 216030 237396 216036 237408
rect 216088 237396 216094 237448
rect 240318 237396 240324 237448
rect 240376 237436 240382 237448
rect 240778 237436 240784 237448
rect 240376 237408 240784 237436
rect 240376 237396 240382 237408
rect 240778 237396 240784 237408
rect 240836 237396 240842 237448
rect 115934 237328 115940 237380
rect 115992 237368 115998 237380
rect 224310 237368 224316 237380
rect 115992 237340 224316 237368
rect 115992 237328 115998 237340
rect 224310 237328 224316 237340
rect 224368 237328 224374 237380
rect 231762 237328 231768 237380
rect 231820 237368 231826 237380
rect 247218 237368 247224 237380
rect 231820 237340 247224 237368
rect 231820 237328 231826 237340
rect 247218 237328 247224 237340
rect 247276 237328 247282 237380
rect 54846 237260 54852 237312
rect 54904 237300 54910 237312
rect 120718 237300 120724 237312
rect 54904 237272 120724 237300
rect 54904 237260 54910 237272
rect 120718 237260 120724 237272
rect 120776 237260 120782 237312
rect 136082 237260 136088 237312
rect 136140 237300 136146 237312
rect 149698 237300 149704 237312
rect 136140 237272 149704 237300
rect 136140 237260 136146 237272
rect 149698 237260 149704 237272
rect 149756 237260 149762 237312
rect 151906 237260 151912 237312
rect 151964 237300 151970 237312
rect 170582 237300 170588 237312
rect 151964 237272 170588 237300
rect 151964 237260 151970 237272
rect 170582 237260 170588 237272
rect 170640 237260 170646 237312
rect 169754 236648 169760 236700
rect 169812 236688 169818 236700
rect 202782 236688 202788 236700
rect 169812 236660 202788 236688
rect 169812 236648 169818 236660
rect 202782 236648 202788 236660
rect 202840 236648 202846 236700
rect 204162 236648 204168 236700
rect 204220 236688 204226 236700
rect 214742 236688 214748 236700
rect 204220 236660 214748 236688
rect 204220 236648 204226 236660
rect 214742 236648 214748 236660
rect 214800 236648 214806 236700
rect 224310 236648 224316 236700
rect 224368 236688 224374 236700
rect 303798 236688 303804 236700
rect 224368 236660 303804 236688
rect 224368 236648 224374 236660
rect 303798 236648 303804 236660
rect 303856 236648 303862 236700
rect 225690 236036 225696 236088
rect 225748 236076 225754 236088
rect 229646 236076 229652 236088
rect 225748 236048 229652 236076
rect 225748 236036 225754 236048
rect 229646 236036 229652 236048
rect 229704 236036 229710 236088
rect 65978 235900 65984 235952
rect 66036 235940 66042 235952
rect 167638 235940 167644 235952
rect 66036 235912 167644 235940
rect 66036 235900 66042 235912
rect 167638 235900 167644 235912
rect 167696 235900 167702 235952
rect 48130 235832 48136 235884
rect 48188 235872 48194 235884
rect 118878 235872 118884 235884
rect 48188 235844 118884 235872
rect 48188 235832 48194 235844
rect 118878 235832 118884 235844
rect 118936 235832 118942 235884
rect 138014 235832 138020 235884
rect 138072 235872 138078 235884
rect 155402 235872 155408 235884
rect 138072 235844 155408 235872
rect 138072 235832 138078 235844
rect 155402 235832 155408 235844
rect 155460 235832 155466 235884
rect 155678 235764 155684 235816
rect 155736 235804 155742 235816
rect 159542 235804 159548 235816
rect 155736 235776 159548 235804
rect 155736 235764 155742 235776
rect 159542 235764 159548 235776
rect 159600 235764 159606 235816
rect 199930 235288 199936 235340
rect 199988 235328 199994 235340
rect 204990 235328 204996 235340
rect 199988 235300 204996 235328
rect 199988 235288 199994 235300
rect 204990 235288 204996 235300
rect 205048 235288 205054 235340
rect 124122 235220 124128 235272
rect 124180 235260 124186 235272
rect 135346 235260 135352 235272
rect 124180 235232 135352 235260
rect 124180 235220 124186 235232
rect 135346 235220 135352 235232
rect 135404 235220 135410 235272
rect 173434 235220 173440 235272
rect 173492 235260 173498 235272
rect 198826 235260 198832 235272
rect 173492 235232 198832 235260
rect 173492 235220 173498 235232
rect 198826 235220 198832 235232
rect 198884 235220 198890 235272
rect 205082 235220 205088 235272
rect 205140 235260 205146 235272
rect 582742 235260 582748 235272
rect 205140 235232 582748 235260
rect 205140 235220 205146 235232
rect 582742 235220 582748 235232
rect 582800 235220 582806 235272
rect 118878 234608 118884 234660
rect 118936 234648 118942 234660
rect 119338 234648 119344 234660
rect 118936 234620 119344 234648
rect 118936 234608 118942 234620
rect 119338 234608 119344 234620
rect 119396 234608 119402 234660
rect 200298 234608 200304 234660
rect 200356 234648 200362 234660
rect 202138 234648 202144 234660
rect 200356 234620 202144 234648
rect 200356 234608 200362 234620
rect 202138 234608 202144 234620
rect 202196 234608 202202 234660
rect 225598 234608 225604 234660
rect 225656 234648 225662 234660
rect 226150 234648 226156 234660
rect 225656 234620 226156 234648
rect 225656 234608 225662 234620
rect 226150 234608 226156 234620
rect 226208 234648 226214 234660
rect 292574 234648 292580 234660
rect 226208 234620 292580 234648
rect 226208 234608 226214 234620
rect 292574 234608 292580 234620
rect 292632 234608 292638 234660
rect 60366 234540 60372 234592
rect 60424 234580 60430 234592
rect 153838 234580 153844 234592
rect 60424 234552 153844 234580
rect 60424 234540 60430 234552
rect 153838 234540 153844 234552
rect 153896 234540 153902 234592
rect 188430 234540 188436 234592
rect 188488 234580 188494 234592
rect 240134 234580 240140 234592
rect 188488 234552 240140 234580
rect 188488 234540 188494 234552
rect 240134 234540 240140 234552
rect 240192 234540 240198 234592
rect 123018 234472 123024 234524
rect 123076 234512 123082 234524
rect 181622 234512 181628 234524
rect 123076 234484 181628 234512
rect 123076 234472 123082 234484
rect 181622 234472 181628 234484
rect 181680 234472 181686 234524
rect 209130 233248 209136 233300
rect 209188 233288 209194 233300
rect 220998 233288 221004 233300
rect 209188 233260 221004 233288
rect 209188 233248 209194 233260
rect 220998 233248 221004 233260
rect 221056 233288 221062 233300
rect 222102 233288 222108 233300
rect 221056 233260 222108 233288
rect 221056 233248 221062 233260
rect 222102 233248 222108 233260
rect 222160 233248 222166 233300
rect 233970 233248 233976 233300
rect 234028 233288 234034 233300
rect 295518 233288 295524 233300
rect 234028 233260 295524 233288
rect 234028 233248 234034 233260
rect 295518 233248 295524 233260
rect 295576 233248 295582 233300
rect 126974 233180 126980 233232
rect 127032 233220 127038 233232
rect 230474 233220 230480 233232
rect 127032 233192 230480 233220
rect 127032 233180 127038 233192
rect 230474 233180 230480 233192
rect 230532 233220 230538 233232
rect 231762 233220 231768 233232
rect 230532 233192 231768 233220
rect 230532 233180 230538 233192
rect 231762 233180 231768 233192
rect 231820 233180 231826 233232
rect 108298 233112 108304 233164
rect 108356 233152 108362 233164
rect 156782 233152 156788 233164
rect 108356 233124 156788 233152
rect 108356 233112 108362 233124
rect 156782 233112 156788 233124
rect 156840 233112 156846 233164
rect 180058 233112 180064 233164
rect 180116 233152 180122 233164
rect 203610 233152 203616 233164
rect 180116 233124 203616 233152
rect 180116 233112 180122 233124
rect 203610 233112 203616 233124
rect 203668 233152 203674 233164
rect 204070 233152 204076 233164
rect 203668 233124 204076 233152
rect 203668 233112 203674 233124
rect 204070 233112 204076 233124
rect 204128 233112 204134 233164
rect 218974 233112 218980 233164
rect 219032 233152 219038 233164
rect 220354 233152 220360 233164
rect 219032 233124 220360 233152
rect 219032 233112 219038 233124
rect 220354 233112 220360 233124
rect 220412 233112 220418 233164
rect 53466 232500 53472 232552
rect 53524 232540 53530 232552
rect 106734 232540 106740 232552
rect 53524 232512 106740 232540
rect 53524 232500 53530 232512
rect 106734 232500 106740 232512
rect 106792 232500 106798 232552
rect 102134 231820 102140 231872
rect 102192 231860 102198 231872
rect 104158 231860 104164 231872
rect 102192 231832 104164 231860
rect 102192 231820 102198 231832
rect 104158 231820 104164 231832
rect 104216 231820 104222 231872
rect 219526 231820 219532 231872
rect 219584 231860 219590 231872
rect 220354 231860 220360 231872
rect 219584 231832 220360 231860
rect 219584 231820 219590 231832
rect 220354 231820 220360 231832
rect 220412 231860 220418 231872
rect 292666 231860 292672 231872
rect 220412 231832 292672 231860
rect 220412 231820 220418 231832
rect 292666 231820 292672 231832
rect 292724 231820 292730 231872
rect 124858 231752 124864 231804
rect 124916 231792 124922 231804
rect 189902 231792 189908 231804
rect 124916 231764 189908 231792
rect 124916 231752 124922 231764
rect 189902 231752 189908 231764
rect 189960 231752 189966 231804
rect 189994 231752 190000 231804
rect 190052 231792 190058 231804
rect 243630 231792 243636 231804
rect 190052 231764 243636 231792
rect 190052 231752 190058 231764
rect 243630 231752 243636 231764
rect 243688 231752 243694 231804
rect 114370 231684 114376 231736
rect 114428 231724 114434 231736
rect 133506 231724 133512 231736
rect 114428 231696 133512 231724
rect 114428 231684 114434 231696
rect 133506 231684 133512 231696
rect 133564 231684 133570 231736
rect 147582 231684 147588 231736
rect 147640 231724 147646 231736
rect 159450 231724 159456 231736
rect 147640 231696 159456 231724
rect 147640 231684 147646 231696
rect 159450 231684 159456 231696
rect 159508 231684 159514 231736
rect 48038 231616 48044 231668
rect 48096 231656 48102 231668
rect 125318 231656 125324 231668
rect 48096 231628 125324 231656
rect 48096 231616 48102 231628
rect 125318 231616 125324 231628
rect 125376 231616 125382 231668
rect 217134 231480 217140 231532
rect 217192 231520 217198 231532
rect 221458 231520 221464 231532
rect 217192 231492 221464 231520
rect 217192 231480 217198 231492
rect 221458 231480 221464 231492
rect 221516 231480 221522 231532
rect 198734 231072 198740 231124
rect 198792 231112 198798 231124
rect 217318 231112 217324 231124
rect 198792 231084 217324 231112
rect 198792 231072 198798 231084
rect 217318 231072 217324 231084
rect 217376 231072 217382 231124
rect 231762 231072 231768 231124
rect 231820 231112 231826 231124
rect 311986 231112 311992 231124
rect 231820 231084 311992 231112
rect 231820 231072 231826 231084
rect 311986 231072 311992 231084
rect 312044 231072 312050 231124
rect 133598 230460 133604 230512
rect 133656 230500 133662 230512
rect 146110 230500 146116 230512
rect 133656 230472 146116 230500
rect 133656 230460 133662 230472
rect 146110 230460 146116 230472
rect 146168 230460 146174 230512
rect 142062 230392 142068 230444
rect 142120 230432 142126 230444
rect 233970 230432 233976 230444
rect 142120 230404 233976 230432
rect 142120 230392 142126 230404
rect 233970 230392 233976 230404
rect 234028 230392 234034 230444
rect 144822 230324 144828 230376
rect 144880 230364 144886 230376
rect 148318 230364 148324 230376
rect 144880 230336 148324 230364
rect 144880 230324 144886 230336
rect 148318 230324 148324 230336
rect 148376 230324 148382 230376
rect 166902 230324 166908 230376
rect 166960 230364 166966 230376
rect 167730 230364 167736 230376
rect 166960 230336 167736 230364
rect 166960 230324 166966 230336
rect 167730 230324 167736 230336
rect 167788 230324 167794 230376
rect 198826 230324 198832 230376
rect 198884 230364 198890 230376
rect 222838 230364 222844 230376
rect 198884 230336 222844 230364
rect 198884 230324 198890 230336
rect 222838 230324 222844 230336
rect 222896 230324 222902 230376
rect 85574 229712 85580 229764
rect 85632 229752 85638 229764
rect 144178 229752 144184 229764
rect 85632 229724 144184 229752
rect 85632 229712 85638 229724
rect 144178 229712 144184 229724
rect 144236 229712 144242 229764
rect 148870 229712 148876 229764
rect 148928 229752 148934 229764
rect 166902 229752 166908 229764
rect 148928 229724 166908 229752
rect 148928 229712 148934 229724
rect 166902 229712 166908 229724
rect 166960 229712 166966 229764
rect 181530 229712 181536 229764
rect 181588 229752 181594 229764
rect 195606 229752 195612 229764
rect 181588 229724 195612 229752
rect 181588 229712 181594 229724
rect 195606 229712 195612 229724
rect 195664 229712 195670 229764
rect 146110 229032 146116 229084
rect 146168 229072 146174 229084
rect 156874 229072 156880 229084
rect 146168 229044 156880 229072
rect 146168 229032 146174 229044
rect 156874 229032 156880 229044
rect 156932 229032 156938 229084
rect 180334 229032 180340 229084
rect 180392 229072 180398 229084
rect 220446 229072 220452 229084
rect 180392 229044 220452 229072
rect 180392 229032 180398 229044
rect 220446 229032 220452 229044
rect 220504 229032 220510 229084
rect 227254 228420 227260 228472
rect 227312 228460 227318 228472
rect 309226 228460 309232 228472
rect 227312 228432 309232 228460
rect 227312 228420 227318 228432
rect 309226 228420 309232 228432
rect 309284 228420 309290 228472
rect 63310 228352 63316 228404
rect 63368 228392 63374 228404
rect 106918 228392 106924 228404
rect 63368 228364 106924 228392
rect 63368 228352 63374 228364
rect 106918 228352 106924 228364
rect 106976 228352 106982 228404
rect 125410 228352 125416 228404
rect 125468 228392 125474 228404
rect 190822 228392 190828 228404
rect 125468 228364 190828 228392
rect 125468 228352 125474 228364
rect 190822 228352 190828 228364
rect 190880 228352 190886 228404
rect 195790 228352 195796 228404
rect 195848 228392 195854 228404
rect 299750 228392 299756 228404
rect 195848 228364 299756 228392
rect 195848 228352 195854 228364
rect 299750 228352 299756 228364
rect 299808 228352 299814 228404
rect 220262 227808 220268 227860
rect 220320 227848 220326 227860
rect 227254 227848 227260 227860
rect 220320 227820 227260 227848
rect 220320 227808 220326 227820
rect 227254 227808 227260 227820
rect 227312 227808 227318 227860
rect 220078 227740 220084 227792
rect 220136 227780 220142 227792
rect 220446 227780 220452 227792
rect 220136 227752 220452 227780
rect 220136 227740 220142 227752
rect 220446 227740 220452 227752
rect 220504 227740 220510 227792
rect 151078 227672 151084 227724
rect 151136 227712 151142 227724
rect 249978 227712 249984 227724
rect 151136 227684 249984 227712
rect 151136 227672 151142 227684
rect 249978 227672 249984 227684
rect 250036 227672 250042 227724
rect 66070 227604 66076 227656
rect 66128 227644 66134 227656
rect 155310 227644 155316 227656
rect 66128 227616 155316 227644
rect 66128 227604 66134 227616
rect 155310 227604 155316 227616
rect 155368 227604 155374 227656
rect 63218 226992 63224 227044
rect 63276 227032 63282 227044
rect 134518 227032 134524 227044
rect 63276 227004 134524 227032
rect 63276 226992 63282 227004
rect 134518 226992 134524 227004
rect 134576 226992 134582 227044
rect 214742 226992 214748 227044
rect 214800 227032 214806 227044
rect 272518 227032 272524 227044
rect 214800 227004 272524 227032
rect 214800 226992 214806 227004
rect 272518 226992 272524 227004
rect 272576 226992 272582 227044
rect 276658 226992 276664 227044
rect 276716 227032 276722 227044
rect 305086 227032 305092 227044
rect 276716 227004 305092 227032
rect 276716 226992 276722 227004
rect 305086 226992 305092 227004
rect 305144 226992 305150 227044
rect 160738 226312 160744 226364
rect 160796 226352 160802 226364
rect 160796 226324 207060 226352
rect 160796 226312 160802 226324
rect 116578 226244 116584 226296
rect 116636 226284 116642 226296
rect 185670 226284 185676 226296
rect 116636 226256 185676 226284
rect 116636 226244 116642 226256
rect 185670 226244 185676 226256
rect 185728 226244 185734 226296
rect 188614 226244 188620 226296
rect 188672 226284 188678 226296
rect 206830 226284 206836 226296
rect 188672 226256 206836 226284
rect 188672 226244 188678 226256
rect 206830 226244 206836 226256
rect 206888 226244 206894 226296
rect 207032 226284 207060 226324
rect 240686 226284 240692 226296
rect 207032 226256 240692 226284
rect 240686 226244 240692 226256
rect 240744 226244 240750 226296
rect 151078 225564 151084 225616
rect 151136 225604 151142 225616
rect 162394 225604 162400 225616
rect 151136 225576 162400 225604
rect 151136 225564 151142 225576
rect 162394 225564 162400 225576
rect 162452 225564 162458 225616
rect 201402 225292 201408 225344
rect 201460 225332 201466 225344
rect 203610 225332 203616 225344
rect 201460 225304 203616 225332
rect 201460 225292 201466 225304
rect 203610 225292 203616 225304
rect 203668 225292 203674 225344
rect 206278 225156 206284 225208
rect 206336 225196 206342 225208
rect 206830 225196 206836 225208
rect 206336 225168 206836 225196
rect 206336 225156 206342 225168
rect 206830 225156 206836 225168
rect 206888 225156 206894 225208
rect 203518 224952 203524 225004
rect 203576 224992 203582 225004
rect 214742 224992 214748 225004
rect 203576 224964 214748 224992
rect 203576 224952 203582 224964
rect 214742 224952 214748 224964
rect 214800 224952 214806 225004
rect 240962 224952 240968 225004
rect 241020 224992 241026 225004
rect 243262 224992 243268 225004
rect 241020 224964 243268 224992
rect 241020 224952 241026 224964
rect 243262 224952 243268 224964
rect 243320 224952 243326 225004
rect 70394 224884 70400 224936
rect 70452 224924 70458 224936
rect 215938 224924 215944 224936
rect 70452 224896 215944 224924
rect 70452 224884 70458 224896
rect 215938 224884 215944 224896
rect 215996 224884 216002 224936
rect 110230 224816 110236 224868
rect 110288 224856 110294 224868
rect 178862 224856 178868 224868
rect 110288 224828 178868 224856
rect 110288 224816 110294 224828
rect 178862 224816 178868 224828
rect 178920 224816 178926 224868
rect 195606 224816 195612 224868
rect 195664 224856 195670 224868
rect 224310 224856 224316 224868
rect 195664 224828 224316 224856
rect 195664 224816 195670 224828
rect 224310 224816 224316 224828
rect 224368 224856 224374 224868
rect 224862 224856 224868 224868
rect 224368 224828 224868 224856
rect 224368 224816 224374 224828
rect 224862 224816 224868 224828
rect 224920 224816 224926 224868
rect 229002 224204 229008 224256
rect 229060 224244 229066 224256
rect 307846 224244 307852 224256
rect 229060 224216 307852 224244
rect 229060 224204 229066 224216
rect 307846 224204 307852 224216
rect 307904 224204 307910 224256
rect 82722 223524 82728 223576
rect 82780 223564 82786 223576
rect 248506 223564 248512 223576
rect 82780 223536 248512 223564
rect 82780 223524 82786 223536
rect 248506 223524 248512 223536
rect 248564 223524 248570 223576
rect 155218 222844 155224 222896
rect 155276 222884 155282 222896
rect 195238 222884 195244 222896
rect 155276 222856 195244 222884
rect 155276 222844 155282 222856
rect 195238 222844 195244 222856
rect 195296 222844 195302 222896
rect 201586 222844 201592 222896
rect 201644 222884 201650 222896
rect 226978 222884 226984 222896
rect 201644 222856 226984 222884
rect 201644 222844 201650 222856
rect 226978 222844 226984 222856
rect 227036 222844 227042 222896
rect 72510 222096 72516 222148
rect 72568 222136 72574 222148
rect 159358 222136 159364 222148
rect 72568 222108 159364 222136
rect 72568 222096 72574 222108
rect 159358 222096 159364 222108
rect 159416 222096 159422 222148
rect 174722 222096 174728 222148
rect 174780 222136 174786 222148
rect 247034 222136 247040 222148
rect 174780 222108 247040 222136
rect 174780 222096 174786 222108
rect 247034 222096 247040 222108
rect 247092 222096 247098 222148
rect 133874 221416 133880 221468
rect 133932 221456 133938 221468
rect 191834 221456 191840 221468
rect 133932 221428 191840 221456
rect 133932 221416 133938 221428
rect 191834 221416 191840 221428
rect 191892 221416 191898 221468
rect 202138 221416 202144 221468
rect 202196 221456 202202 221468
rect 294138 221456 294144 221468
rect 202196 221428 294144 221456
rect 202196 221416 202202 221428
rect 294138 221416 294144 221428
rect 294196 221416 294202 221468
rect 580902 221144 580908 221196
rect 580960 221184 580966 221196
rect 583570 221184 583576 221196
rect 580960 221156 583576 221184
rect 580960 221144 580966 221156
rect 583570 221144 583576 221156
rect 583628 221144 583634 221196
rect 4798 220804 4804 220856
rect 4856 220844 4862 220856
rect 93762 220844 93768 220856
rect 4856 220816 93768 220844
rect 4856 220804 4862 220816
rect 93762 220804 93768 220816
rect 93820 220804 93826 220856
rect 148318 220736 148324 220788
rect 148376 220776 148382 220788
rect 236914 220776 236920 220788
rect 148376 220748 236920 220776
rect 148376 220736 148382 220748
rect 236914 220736 236920 220748
rect 236972 220736 236978 220788
rect 107470 220668 107476 220720
rect 107528 220708 107534 220720
rect 158070 220708 158076 220720
rect 107528 220680 158076 220708
rect 107528 220668 107534 220680
rect 158070 220668 158076 220680
rect 158128 220668 158134 220720
rect 166350 220668 166356 220720
rect 166408 220708 166414 220720
rect 223758 220708 223764 220720
rect 166408 220680 223764 220708
rect 166408 220668 166414 220680
rect 223758 220668 223764 220680
rect 223816 220668 223822 220720
rect 236914 220056 236920 220108
rect 236972 220096 236978 220108
rect 306650 220096 306656 220108
rect 236972 220068 306656 220096
rect 236972 220056 236978 220068
rect 306650 220056 306656 220068
rect 306708 220056 306714 220108
rect 223758 219920 223764 219972
rect 223816 219960 223822 219972
rect 224218 219960 224224 219972
rect 223816 219932 224224 219960
rect 223816 219920 223822 219932
rect 224218 219920 224224 219932
rect 224276 219920 224282 219972
rect 130930 219376 130936 219428
rect 130988 219416 130994 219428
rect 186958 219416 186964 219428
rect 130988 219388 186964 219416
rect 130988 219376 130994 219388
rect 186958 219376 186964 219388
rect 187016 219376 187022 219428
rect 565078 219376 565084 219428
rect 565136 219416 565142 219428
rect 580166 219416 580172 219428
rect 565136 219388 580172 219416
rect 565136 219376 565142 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 171962 219308 171968 219360
rect 172020 219348 172026 219360
rect 223390 219348 223396 219360
rect 172020 219320 223396 219348
rect 172020 219308 172026 219320
rect 223390 219308 223396 219320
rect 223448 219308 223454 219360
rect 81250 218764 81256 218816
rect 81308 218804 81314 218816
rect 128354 218804 128360 218816
rect 81308 218776 128360 218804
rect 81308 218764 81314 218776
rect 128354 218764 128360 218776
rect 128412 218764 128418 218816
rect 21358 218696 21364 218748
rect 21416 218736 21422 218748
rect 156598 218736 156604 218748
rect 21416 218708 156604 218736
rect 21416 218696 21422 218708
rect 156598 218696 156604 218708
rect 156656 218696 156662 218748
rect 224402 218696 224408 218748
rect 224460 218736 224466 218748
rect 238846 218736 238852 218748
rect 224460 218708 238852 218736
rect 224460 218696 224466 218708
rect 238846 218696 238852 218708
rect 238904 218696 238910 218748
rect 222930 218084 222936 218136
rect 222988 218124 222994 218136
rect 223390 218124 223396 218136
rect 222988 218096 223396 218124
rect 222988 218084 222994 218096
rect 223390 218084 223396 218096
rect 223448 218084 223454 218136
rect 186958 218016 186964 218068
rect 187016 218056 187022 218068
rect 187142 218056 187148 218068
rect 187016 218028 187148 218056
rect 187016 218016 187022 218028
rect 187142 218016 187148 218028
rect 187200 218016 187206 218068
rect 104802 217268 104808 217320
rect 104860 217308 104866 217320
rect 172790 217308 172796 217320
rect 104860 217280 172796 217308
rect 104860 217268 104866 217280
rect 172790 217268 172796 217280
rect 172848 217268 172854 217320
rect 187510 217268 187516 217320
rect 187568 217308 187574 217320
rect 197998 217308 198004 217320
rect 187568 217280 198004 217308
rect 187568 217268 187574 217280
rect 197998 217268 198004 217280
rect 198056 217268 198062 217320
rect 206278 217268 206284 217320
rect 206336 217308 206342 217320
rect 236638 217308 236644 217320
rect 206336 217280 236644 217308
rect 206336 217268 206342 217280
rect 236638 217268 236644 217280
rect 236696 217268 236702 217320
rect 236730 217268 236736 217320
rect 236788 217308 236794 217320
rect 254026 217308 254032 217320
rect 236788 217280 254032 217308
rect 236788 217268 236794 217280
rect 254026 217268 254032 217280
rect 254084 217268 254090 217320
rect 254578 217268 254584 217320
rect 254636 217308 254642 217320
rect 317414 217308 317420 217320
rect 254636 217280 317420 217308
rect 254636 217268 254642 217280
rect 317414 217268 317420 217280
rect 317472 217268 317478 217320
rect 142798 216656 142804 216708
rect 142856 216696 142862 216708
rect 234614 216696 234620 216708
rect 142856 216668 234620 216696
rect 142856 216656 142862 216668
rect 234614 216656 234620 216668
rect 234672 216656 234678 216708
rect 131022 216588 131028 216640
rect 131080 216628 131086 216640
rect 191190 216628 191196 216640
rect 131080 216600 191196 216628
rect 131080 216588 131086 216600
rect 191190 216588 191196 216600
rect 191248 216588 191254 216640
rect 191834 216588 191840 216640
rect 191892 216628 191898 216640
rect 241514 216628 241520 216640
rect 191892 216600 241520 216628
rect 191892 216588 191898 216600
rect 241514 216588 241520 216600
rect 241572 216628 241578 216640
rect 242250 216628 242256 216640
rect 241572 216600 242256 216628
rect 241572 216588 241578 216600
rect 242250 216588 242256 216600
rect 242308 216588 242314 216640
rect 111794 215908 111800 215960
rect 111852 215948 111858 215960
rect 191650 215948 191656 215960
rect 111852 215920 191656 215948
rect 111852 215908 111858 215920
rect 191650 215908 191656 215920
rect 191708 215908 191714 215960
rect 200022 215908 200028 215960
rect 200080 215948 200086 215960
rect 230474 215948 230480 215960
rect 200080 215920 230480 215948
rect 200080 215908 200086 215920
rect 230474 215908 230480 215920
rect 230532 215908 230538 215960
rect 67726 215228 67732 215280
rect 67784 215268 67790 215280
rect 206462 215268 206468 215280
rect 67784 215240 206468 215268
rect 67784 215228 67790 215240
rect 206462 215228 206468 215240
rect 206520 215228 206526 215280
rect 73890 215160 73896 215212
rect 73948 215200 73954 215212
rect 151078 215200 151084 215212
rect 73948 215172 151084 215200
rect 73948 215160 73954 215172
rect 151078 215160 151084 215172
rect 151136 215160 151142 215212
rect 205082 214616 205088 214668
rect 205140 214656 205146 214668
rect 245654 214656 245660 214668
rect 205140 214628 245660 214656
rect 205140 214616 205146 214628
rect 245654 214616 245660 214628
rect 245712 214616 245718 214668
rect 238110 214548 238116 214600
rect 238168 214588 238174 214600
rect 309318 214588 309324 214600
rect 238168 214560 309324 214588
rect 238168 214548 238174 214560
rect 309318 214548 309324 214560
rect 309376 214548 309382 214600
rect 233234 214344 233240 214396
rect 233292 214384 233298 214396
rect 234430 214384 234436 214396
rect 233292 214356 234436 214384
rect 233292 214344 233298 214356
rect 234430 214344 234436 214356
rect 234488 214344 234494 214396
rect 212994 213936 213000 213988
rect 213052 213976 213058 213988
rect 233234 213976 233240 213988
rect 213052 213948 233240 213976
rect 213052 213936 213058 213948
rect 233234 213936 233240 213948
rect 233292 213936 233298 213988
rect 64690 213868 64696 213920
rect 64748 213908 64754 213920
rect 191926 213908 191932 213920
rect 64748 213880 191932 213908
rect 64748 213868 64754 213880
rect 191926 213868 191932 213880
rect 191984 213868 191990 213920
rect 191650 213800 191656 213852
rect 191708 213840 191714 213852
rect 222286 213840 222292 213852
rect 191708 213812 222292 213840
rect 191708 213800 191714 213812
rect 222286 213800 222292 213812
rect 222344 213840 222350 213852
rect 223022 213840 223028 213852
rect 222344 213812 223028 213840
rect 222344 213800 222350 213812
rect 223022 213800 223028 213812
rect 223080 213800 223086 213852
rect 197354 213256 197360 213308
rect 197412 213296 197418 213308
rect 214834 213296 214840 213308
rect 197412 213268 214840 213296
rect 197412 213256 197418 213268
rect 214834 213256 214840 213268
rect 214892 213256 214898 213308
rect 134518 213188 134524 213240
rect 134576 213228 134582 213240
rect 186958 213228 186964 213240
rect 134576 213200 186964 213228
rect 134576 213188 134582 213200
rect 186958 213188 186964 213200
rect 187016 213188 187022 213240
rect 214650 213188 214656 213240
rect 214708 213228 214714 213240
rect 302510 213228 302516 213240
rect 214708 213200 302516 213228
rect 214708 213188 214714 213200
rect 302510 213188 302516 213200
rect 302568 213188 302574 213240
rect 249058 212780 249064 212832
rect 249116 212820 249122 212832
rect 251266 212820 251272 212832
rect 249116 212792 251272 212820
rect 249116 212780 249122 212792
rect 251266 212780 251272 212792
rect 251324 212780 251330 212832
rect 122834 212440 122840 212492
rect 122892 212480 122898 212492
rect 227806 212480 227812 212492
rect 122892 212452 227812 212480
rect 122892 212440 122898 212452
rect 227806 212440 227812 212452
rect 227864 212480 227870 212492
rect 228358 212480 228364 212492
rect 227864 212452 228364 212480
rect 227864 212440 227870 212452
rect 228358 212440 228364 212452
rect 228416 212440 228422 212492
rect 77386 212372 77392 212424
rect 77444 212412 77450 212424
rect 147674 212412 147680 212424
rect 77444 212384 147680 212412
rect 77444 212372 77450 212384
rect 147674 212372 147680 212384
rect 147732 212372 147738 212424
rect 195238 212372 195244 212424
rect 195296 212412 195302 212424
rect 245746 212412 245752 212424
rect 195296 212384 245752 212412
rect 195296 212372 195302 212384
rect 245746 212372 245752 212384
rect 245804 212372 245810 212424
rect 148962 211760 148968 211812
rect 149020 211800 149026 211812
rect 171778 211800 171784 211812
rect 149020 211772 171784 211800
rect 149020 211760 149026 211772
rect 171778 211760 171784 211772
rect 171836 211760 171842 211812
rect 172422 211148 172428 211200
rect 172480 211188 172486 211200
rect 192478 211188 192484 211200
rect 172480 211160 192484 211188
rect 172480 211148 172486 211160
rect 192478 211148 192484 211160
rect 192536 211148 192542 211200
rect 237374 211148 237380 211200
rect 237432 211188 237438 211200
rect 238294 211188 238300 211200
rect 237432 211160 238300 211188
rect 237432 211148 237438 211160
rect 238294 211148 238300 211160
rect 238352 211188 238358 211200
rect 246298 211188 246304 211200
rect 238352 211160 246304 211188
rect 238352 211148 238358 211160
rect 246298 211148 246304 211160
rect 246356 211148 246362 211200
rect 76650 211080 76656 211132
rect 76708 211120 76714 211132
rect 212994 211120 213000 211132
rect 76708 211092 213000 211120
rect 76708 211080 76714 211092
rect 212994 211080 213000 211092
rect 213052 211080 213058 211132
rect 104894 211012 104900 211064
rect 104952 211052 104958 211064
rect 188522 211052 188528 211064
rect 104952 211024 188528 211052
rect 104952 211012 104958 211024
rect 188522 211012 188528 211024
rect 188580 211012 188586 211064
rect 214834 210468 214840 210520
rect 214892 210508 214898 210520
rect 251266 210508 251272 210520
rect 214892 210480 251272 210508
rect 214892 210468 214898 210480
rect 251266 210468 251272 210480
rect 251324 210468 251330 210520
rect 214742 210400 214748 210452
rect 214800 210440 214806 210452
rect 302418 210440 302424 210452
rect 214800 210412 302424 210440
rect 214800 210400 214806 210412
rect 302418 210400 302424 210412
rect 302476 210400 302482 210452
rect 132402 209720 132408 209772
rect 132460 209760 132466 209772
rect 244458 209760 244464 209772
rect 132460 209732 244464 209760
rect 132460 209720 132466 209732
rect 244458 209720 244464 209732
rect 244516 209720 244522 209772
rect 75270 209652 75276 209704
rect 75328 209692 75334 209704
rect 142798 209692 142804 209704
rect 75328 209664 142804 209692
rect 75328 209652 75334 209664
rect 142798 209652 142804 209664
rect 142856 209652 142862 209704
rect 144178 209040 144184 209092
rect 144236 209080 144242 209092
rect 213730 209080 213736 209092
rect 144236 209052 213736 209080
rect 144236 209040 144242 209052
rect 213730 209040 213736 209052
rect 213788 209040 213794 209092
rect 213730 208360 213736 208412
rect 213788 208400 213794 208412
rect 238110 208400 238116 208412
rect 213788 208372 238116 208400
rect 213788 208360 213794 208372
rect 238110 208360 238116 208372
rect 238168 208360 238174 208412
rect 113082 208292 113088 208344
rect 113140 208332 113146 208344
rect 247126 208332 247132 208344
rect 113140 208304 247132 208332
rect 113140 208292 113146 208304
rect 247126 208292 247132 208304
rect 247184 208292 247190 208344
rect 69014 207612 69020 207664
rect 69072 207652 69078 207664
rect 200022 207652 200028 207664
rect 69072 207624 200028 207652
rect 69072 207612 69078 207624
rect 200022 207612 200028 207624
rect 200080 207612 200086 207664
rect 57698 206932 57704 206984
rect 57756 206972 57762 206984
rect 209038 206972 209044 206984
rect 57756 206944 209044 206972
rect 57756 206932 57762 206944
rect 209038 206932 209044 206944
rect 209096 206932 209102 206984
rect 99466 206864 99472 206916
rect 99524 206904 99530 206916
rect 211798 206904 211804 206916
rect 99524 206876 211804 206904
rect 99524 206864 99530 206876
rect 211798 206864 211804 206876
rect 211856 206904 211862 206916
rect 212442 206904 212448 206916
rect 211856 206876 212448 206904
rect 211856 206864 211862 206876
rect 212442 206864 212448 206876
rect 212500 206864 212506 206916
rect 212442 206320 212448 206372
rect 212500 206360 212506 206372
rect 231118 206360 231124 206372
rect 212500 206332 231124 206360
rect 212500 206320 212506 206332
rect 231118 206320 231124 206332
rect 231176 206320 231182 206372
rect 220170 206252 220176 206304
rect 220228 206292 220234 206304
rect 295610 206292 295616 206304
rect 220228 206264 295616 206292
rect 220228 206252 220234 206264
rect 295610 206252 295616 206264
rect 295668 206252 295674 206304
rect 95234 205572 95240 205624
rect 95292 205612 95298 205624
rect 244274 205612 244280 205624
rect 95292 205584 244280 205612
rect 95292 205572 95298 205584
rect 244274 205572 244280 205584
rect 244332 205572 244338 205624
rect 195330 204960 195336 205012
rect 195388 205000 195394 205012
rect 218882 205000 218888 205012
rect 195388 204972 218888 205000
rect 195388 204960 195394 204972
rect 218882 204960 218888 204972
rect 218940 204960 218946 205012
rect 83458 204892 83464 204944
rect 83516 204932 83522 204944
rect 166994 204932 167000 204944
rect 83516 204904 167000 204932
rect 83516 204892 83522 204904
rect 166994 204892 167000 204904
rect 167052 204892 167058 204944
rect 218790 204892 218796 204944
rect 218848 204932 218854 204944
rect 283006 204932 283012 204944
rect 218848 204904 283012 204932
rect 218848 204892 218854 204904
rect 283006 204892 283012 204904
rect 283064 204892 283070 204944
rect 137922 204212 137928 204264
rect 137980 204252 137986 204264
rect 232130 204252 232136 204264
rect 137980 204224 232136 204252
rect 137980 204212 137986 204224
rect 232130 204212 232136 204224
rect 232188 204252 232194 204264
rect 233142 204252 233148 204264
rect 232188 204224 233148 204252
rect 232188 204212 232194 204224
rect 233142 204212 233148 204224
rect 233200 204212 233206 204264
rect 191190 203668 191196 203720
rect 191248 203708 191254 203720
rect 231946 203708 231952 203720
rect 191248 203680 231952 203708
rect 191248 203668 191254 203680
rect 231946 203668 231952 203680
rect 232004 203668 232010 203720
rect 146202 203532 146208 203584
rect 146260 203572 146266 203584
rect 191282 203572 191288 203584
rect 146260 203544 191288 203572
rect 146260 203532 146266 203544
rect 191282 203532 191288 203544
rect 191340 203532 191346 203584
rect 233142 203532 233148 203584
rect 233200 203572 233206 203584
rect 303706 203572 303712 203584
rect 233200 203544 303712 203572
rect 233200 203532 233206 203544
rect 303706 203532 303712 203544
rect 303764 203532 303770 203584
rect 3050 202784 3056 202836
rect 3108 202824 3114 202836
rect 124122 202824 124128 202836
rect 3108 202796 124128 202824
rect 3108 202784 3114 202796
rect 124122 202784 124128 202796
rect 124180 202784 124186 202836
rect 125502 202784 125508 202836
rect 125560 202824 125566 202836
rect 251450 202824 251456 202836
rect 125560 202796 251456 202824
rect 125560 202784 125566 202796
rect 251450 202784 251456 202796
rect 251508 202784 251514 202836
rect 166994 202716 167000 202768
rect 167052 202756 167058 202768
rect 202874 202756 202880 202768
rect 167052 202728 202880 202756
rect 167052 202716 167058 202728
rect 202874 202716 202880 202728
rect 202932 202756 202938 202768
rect 203518 202756 203524 202768
rect 202932 202728 203524 202756
rect 202932 202716 202938 202728
rect 203518 202716 203524 202728
rect 203576 202716 203582 202768
rect 83090 202104 83096 202156
rect 83148 202144 83154 202156
rect 166810 202144 166816 202156
rect 83148 202116 166816 202144
rect 83148 202104 83154 202116
rect 166810 202104 166816 202116
rect 166868 202104 166874 202156
rect 282178 201532 282184 201544
rect 224972 201504 282184 201532
rect 200022 201424 200028 201476
rect 200080 201464 200086 201476
rect 224972 201464 225000 201504
rect 282178 201492 282184 201504
rect 282236 201492 282242 201544
rect 200080 201436 225000 201464
rect 200080 201424 200086 201436
rect 76558 201356 76564 201408
rect 76616 201396 76622 201408
rect 200850 201396 200856 201408
rect 76616 201368 200856 201396
rect 76616 201356 76622 201368
rect 200850 201356 200856 201368
rect 200908 201356 200914 201408
rect 225690 200812 225696 200864
rect 225748 200852 225754 200864
rect 291286 200852 291292 200864
rect 225748 200824 291292 200852
rect 225748 200812 225754 200824
rect 291286 200812 291292 200824
rect 291344 200812 291350 200864
rect 86862 200744 86868 200796
rect 86920 200784 86926 200796
rect 189718 200784 189724 200796
rect 86920 200756 189724 200784
rect 86920 200744 86926 200756
rect 189718 200744 189724 200756
rect 189776 200744 189782 200796
rect 204990 200744 204996 200796
rect 205048 200784 205054 200796
rect 285766 200784 285772 200796
rect 205048 200756 285772 200784
rect 205048 200744 205054 200756
rect 285766 200744 285772 200756
rect 285824 200744 285830 200796
rect 93118 200064 93124 200116
rect 93176 200104 93182 200116
rect 198734 200104 198740 200116
rect 93176 200076 198740 200104
rect 93176 200064 93182 200076
rect 198734 200064 198740 200076
rect 198792 200064 198798 200116
rect 223022 199452 223028 199504
rect 223080 199492 223086 199504
rect 279050 199492 279056 199504
rect 223080 199464 279056 199492
rect 223080 199452 223086 199464
rect 279050 199452 279056 199464
rect 279108 199452 279114 199504
rect 118602 199384 118608 199436
rect 118660 199424 118666 199436
rect 202138 199424 202144 199436
rect 118660 199396 202144 199424
rect 118660 199384 118666 199396
rect 202138 199384 202144 199396
rect 202196 199384 202202 199436
rect 211890 199384 211896 199436
rect 211948 199424 211954 199436
rect 305178 199424 305184 199436
rect 211948 199396 305184 199424
rect 211948 199384 211954 199396
rect 305178 199384 305184 199396
rect 305236 199384 305242 199436
rect 50798 198636 50804 198688
rect 50856 198676 50862 198688
rect 180242 198676 180248 198688
rect 50856 198648 180248 198676
rect 50856 198636 50862 198648
rect 180242 198636 180248 198648
rect 180300 198636 180306 198688
rect 191282 198636 191288 198688
rect 191340 198676 191346 198688
rect 191340 198648 238754 198676
rect 191340 198636 191346 198648
rect 97810 198568 97816 198620
rect 97868 198608 97874 198620
rect 158714 198608 158720 198620
rect 97868 198580 158720 198608
rect 97868 198568 97874 198580
rect 158714 198568 158720 198580
rect 158772 198568 158778 198620
rect 166810 198568 166816 198620
rect 166868 198608 166874 198620
rect 207658 198608 207664 198620
rect 166868 198580 207664 198608
rect 166868 198568 166874 198580
rect 207658 198568 207664 198580
rect 207716 198568 207722 198620
rect 238726 198540 238754 198648
rect 244274 198540 244280 198552
rect 238726 198512 244280 198540
rect 244274 198500 244280 198512
rect 244332 198540 244338 198552
rect 244918 198540 244924 198552
rect 244332 198512 244924 198540
rect 244332 198500 244338 198512
rect 244918 198500 244924 198512
rect 244976 198500 244982 198552
rect 46842 197276 46848 197328
rect 46900 197316 46906 197328
rect 173250 197316 173256 197328
rect 46900 197288 173256 197316
rect 46900 197276 46906 197288
rect 173250 197276 173256 197288
rect 173308 197276 173314 197328
rect 143442 197208 143448 197260
rect 143500 197248 143506 197260
rect 163498 197248 163504 197260
rect 143500 197220 163504 197248
rect 143500 197208 143506 197220
rect 163498 197208 163504 197220
rect 163556 197208 163562 197260
rect 174630 196596 174636 196648
rect 174688 196636 174694 196648
rect 212074 196636 212080 196648
rect 174688 196608 212080 196636
rect 174688 196596 174694 196608
rect 212074 196596 212080 196608
rect 212132 196596 212138 196648
rect 213822 196596 213828 196648
rect 213880 196636 213886 196648
rect 226978 196636 226984 196648
rect 213880 196608 226984 196636
rect 213880 196596 213886 196608
rect 226978 196596 226984 196608
rect 227036 196596 227042 196648
rect 223022 195984 223028 196036
rect 223080 196024 223086 196036
rect 249886 196024 249892 196036
rect 223080 195996 249892 196024
rect 223080 195984 223086 195996
rect 249886 195984 249892 195996
rect 249944 195984 249950 196036
rect 79870 195916 79876 195968
rect 79928 195956 79934 195968
rect 226334 195956 226340 195968
rect 79928 195928 226340 195956
rect 79928 195916 79934 195928
rect 226334 195916 226340 195928
rect 226392 195916 226398 195968
rect 106918 195848 106924 195900
rect 106976 195888 106982 195900
rect 214558 195888 214564 195900
rect 106976 195860 214564 195888
rect 106976 195848 106982 195860
rect 214558 195848 214564 195860
rect 214616 195848 214622 195900
rect 218882 195236 218888 195288
rect 218940 195276 218946 195288
rect 237466 195276 237472 195288
rect 218940 195248 237472 195276
rect 218940 195236 218946 195248
rect 237466 195236 237472 195248
rect 237524 195236 237530 195288
rect 63126 194488 63132 194540
rect 63184 194528 63190 194540
rect 210418 194528 210424 194540
rect 63184 194500 210424 194528
rect 63184 194488 63190 194500
rect 210418 194488 210424 194500
rect 210476 194488 210482 194540
rect 212074 193876 212080 193928
rect 212132 193916 212138 193928
rect 232498 193916 232504 193928
rect 212132 193888 232504 193916
rect 212132 193876 212138 193888
rect 232498 193876 232504 193888
rect 232556 193876 232562 193928
rect 81342 193808 81348 193860
rect 81400 193848 81406 193860
rect 176010 193848 176016 193860
rect 81400 193820 176016 193848
rect 81400 193808 81406 193820
rect 176010 193808 176016 193820
rect 176068 193808 176074 193860
rect 199378 193808 199384 193860
rect 199436 193848 199442 193860
rect 230566 193848 230572 193860
rect 199436 193820 230572 193848
rect 199436 193808 199442 193820
rect 230566 193808 230572 193820
rect 230624 193808 230630 193860
rect 238018 193808 238024 193860
rect 238076 193848 238082 193860
rect 281718 193848 281724 193860
rect 238076 193820 281724 193848
rect 238076 193808 238082 193820
rect 281718 193808 281724 193820
rect 281776 193808 281782 193860
rect 166902 192516 166908 192568
rect 166960 192556 166966 192568
rect 237374 192556 237380 192568
rect 166960 192528 237380 192556
rect 166960 192516 166966 192528
rect 237374 192516 237380 192528
rect 237432 192516 237438 192568
rect 72418 192448 72424 192500
rect 72476 192488 72482 192500
rect 171962 192488 171968 192500
rect 72476 192460 171968 192488
rect 72476 192448 72482 192460
rect 171962 192448 171968 192460
rect 172020 192448 172026 192500
rect 207658 192448 207664 192500
rect 207716 192488 207722 192500
rect 287330 192488 287336 192500
rect 207716 192460 287336 192488
rect 207716 192448 207722 192460
rect 287330 192448 287336 192460
rect 287388 192448 287394 192500
rect 73154 191768 73160 191820
rect 73212 191808 73218 191820
rect 202598 191808 202604 191820
rect 73212 191780 202604 191808
rect 73212 191768 73218 191780
rect 202598 191768 202604 191780
rect 202656 191768 202662 191820
rect 206370 191156 206376 191208
rect 206428 191196 206434 191208
rect 301038 191196 301044 191208
rect 206428 191168 301044 191196
rect 206428 191156 206434 191168
rect 301038 191156 301044 191168
rect 301096 191156 301102 191208
rect 192570 191088 192576 191140
rect 192628 191128 192634 191140
rect 292758 191128 292764 191140
rect 192628 191100 292764 191128
rect 192628 191088 192634 191100
rect 292758 191088 292764 191100
rect 292816 191088 292822 191140
rect 133782 190476 133788 190528
rect 133840 190516 133846 190528
rect 192662 190516 192668 190528
rect 133840 190488 192668 190516
rect 133840 190476 133846 190488
rect 192662 190476 192668 190488
rect 192720 190476 192726 190528
rect 89530 189728 89536 189780
rect 89588 189768 89594 189780
rect 191190 189768 191196 189780
rect 89588 189740 191196 189768
rect 89588 189728 89594 189740
rect 191190 189728 191196 189740
rect 191248 189728 191254 189780
rect 194502 189728 194508 189780
rect 194560 189768 194566 189780
rect 220722 189768 220728 189780
rect 194560 189740 220728 189768
rect 194560 189728 194566 189740
rect 220722 189728 220728 189740
rect 220780 189728 220786 189780
rect 266998 189728 267004 189780
rect 267056 189768 267062 189780
rect 307938 189768 307944 189780
rect 267056 189740 307944 189768
rect 267056 189728 267062 189740
rect 307938 189728 307944 189740
rect 307996 189728 308002 189780
rect 170582 189156 170588 189168
rect 161446 189128 170588 189156
rect 113082 189048 113088 189100
rect 113140 189088 113146 189100
rect 161446 189088 161474 189128
rect 170582 189116 170588 189128
rect 170640 189116 170646 189168
rect 221458 189116 221464 189168
rect 221516 189156 221522 189168
rect 234706 189156 234712 189168
rect 221516 189128 234712 189156
rect 221516 189116 221522 189128
rect 234706 189116 234712 189128
rect 234764 189116 234770 189168
rect 113140 189060 161474 189088
rect 113140 189048 113146 189060
rect 169754 189048 169760 189100
rect 169812 189088 169818 189100
rect 335354 189088 335360 189100
rect 169812 189060 335360 189088
rect 169812 189048 169818 189060
rect 335354 189048 335360 189060
rect 335412 189048 335418 189100
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 35158 189020 35164 189032
rect 3568 188992 35164 189020
rect 3568 188980 3574 188992
rect 35158 188980 35164 188992
rect 35216 188980 35222 189032
rect 89622 188980 89628 189032
rect 89680 189020 89686 189032
rect 223022 189020 223028 189032
rect 89680 188992 223028 189020
rect 89680 188980 89686 188992
rect 223022 188980 223028 188992
rect 223080 188980 223086 189032
rect 240778 188368 240784 188420
rect 240836 188408 240842 188420
rect 279142 188408 279148 188420
rect 240836 188380 279148 188408
rect 240836 188368 240842 188380
rect 279142 188368 279148 188380
rect 279200 188368 279206 188420
rect 191742 188300 191748 188352
rect 191800 188340 191806 188352
rect 214558 188340 214564 188352
rect 191800 188312 214564 188340
rect 191800 188300 191806 188312
rect 214558 188300 214564 188312
rect 214616 188300 214622 188352
rect 224310 188300 224316 188352
rect 224368 188340 224374 188352
rect 236086 188340 236092 188352
rect 224368 188312 236092 188340
rect 224368 188300 224374 188312
rect 236086 188300 236092 188312
rect 236144 188300 236150 188352
rect 236730 188300 236736 188352
rect 236788 188340 236794 188352
rect 283190 188340 283196 188352
rect 236788 188312 283196 188340
rect 236788 188300 236794 188312
rect 283190 188300 283196 188312
rect 283248 188300 283254 188352
rect 304258 188300 304264 188352
rect 304316 188340 304322 188352
rect 325694 188340 325700 188352
rect 304316 188312 325700 188340
rect 304316 188300 304322 188312
rect 325694 188300 325700 188312
rect 325752 188300 325758 188352
rect 131022 187688 131028 187740
rect 131080 187728 131086 187740
rect 188614 187728 188620 187740
rect 131080 187700 188620 187728
rect 131080 187688 131086 187700
rect 188614 187688 188620 187700
rect 188672 187688 188678 187740
rect 52270 187620 52276 187672
rect 52328 187660 52334 187672
rect 221458 187660 221464 187672
rect 52328 187632 221464 187660
rect 52328 187620 52334 187632
rect 221458 187620 221464 187632
rect 221516 187620 221522 187672
rect 280798 187620 280804 187672
rect 280856 187660 280862 187672
rect 288618 187660 288624 187672
rect 280856 187632 288624 187660
rect 280856 187620 280862 187632
rect 288618 187620 288624 187632
rect 288676 187620 288682 187672
rect 180702 186940 180708 186992
rect 180760 186980 180766 186992
rect 237558 186980 237564 186992
rect 180760 186952 237564 186980
rect 180760 186940 180766 186952
rect 237558 186940 237564 186952
rect 237616 186940 237622 186992
rect 128262 186328 128268 186380
rect 128320 186368 128326 186380
rect 174630 186368 174636 186380
rect 128320 186340 174636 186368
rect 128320 186328 128326 186340
rect 174630 186328 174636 186340
rect 174688 186328 174694 186380
rect 222102 186328 222108 186380
rect 222160 186368 222166 186380
rect 293954 186368 293960 186380
rect 222160 186340 293960 186368
rect 222160 186328 222166 186340
rect 293954 186328 293960 186340
rect 294012 186328 294018 186380
rect 188522 185648 188528 185700
rect 188580 185688 188586 185700
rect 231210 185688 231216 185700
rect 188580 185660 231216 185688
rect 188580 185648 188586 185660
rect 231210 185648 231216 185660
rect 231268 185648 231274 185700
rect 220262 185580 220268 185632
rect 220320 185620 220326 185632
rect 280154 185620 280160 185632
rect 220320 185592 280160 185620
rect 220320 185580 220326 185592
rect 280154 185580 280160 185592
rect 280212 185580 280218 185632
rect 106182 184968 106188 185020
rect 106240 185008 106246 185020
rect 182910 185008 182916 185020
rect 106240 184980 182916 185008
rect 106240 184968 106246 184980
rect 182910 184968 182916 184980
rect 182968 184968 182974 185020
rect 121362 184900 121368 184952
rect 121420 184940 121426 184952
rect 207658 184940 207664 184952
rect 121420 184912 207664 184940
rect 121420 184900 121426 184912
rect 207658 184900 207664 184912
rect 207716 184900 207722 184952
rect 200758 184220 200764 184272
rect 200816 184260 200822 184272
rect 235994 184260 236000 184272
rect 200816 184232 236000 184260
rect 200816 184220 200822 184232
rect 235994 184220 236000 184232
rect 236052 184220 236058 184272
rect 184842 184152 184848 184204
rect 184900 184192 184906 184204
rect 303890 184192 303896 184204
rect 184900 184164 303896 184192
rect 184900 184152 184906 184164
rect 303890 184152 303896 184164
rect 303948 184152 303954 184204
rect 243814 183744 243820 183796
rect 243872 183784 243878 183796
rect 245746 183784 245752 183796
rect 243872 183756 245752 183784
rect 243872 183744 243878 183756
rect 245746 183744 245752 183756
rect 245804 183744 245810 183796
rect 100662 183608 100668 183660
rect 100720 183648 100726 183660
rect 180242 183648 180248 183660
rect 100720 183620 180248 183648
rect 100720 183608 100726 183620
rect 180242 183608 180248 183620
rect 180300 183608 180306 183660
rect 108942 183540 108948 183592
rect 109000 183580 109006 183592
rect 195330 183580 195336 183592
rect 109000 183552 195336 183580
rect 109000 183540 109006 183552
rect 195330 183540 195336 183552
rect 195388 183540 195394 183592
rect 203610 182860 203616 182912
rect 203668 182900 203674 182912
rect 238754 182900 238760 182912
rect 203668 182872 238760 182900
rect 203668 182860 203674 182872
rect 238754 182860 238760 182872
rect 238812 182860 238818 182912
rect 271322 182860 271328 182912
rect 271380 182900 271386 182912
rect 281810 182900 281816 182912
rect 271380 182872 281816 182900
rect 271380 182860 271386 182872
rect 281810 182860 281816 182872
rect 281868 182860 281874 182912
rect 178862 182792 178868 182844
rect 178920 182832 178926 182844
rect 284478 182832 284484 182844
rect 178920 182804 284484 182832
rect 178920 182792 178926 182804
rect 284478 182792 284484 182804
rect 284536 182792 284542 182844
rect 132402 182248 132408 182300
rect 132460 182288 132466 182300
rect 172054 182288 172060 182300
rect 132460 182260 172060 182288
rect 132460 182248 132466 182260
rect 172054 182248 172060 182260
rect 172112 182248 172118 182300
rect 102042 182180 102048 182232
rect 102100 182220 102106 182232
rect 167730 182220 167736 182232
rect 102100 182192 167736 182220
rect 102100 182180 102106 182192
rect 167730 182180 167736 182192
rect 167788 182180 167794 182232
rect 209130 181500 209136 181552
rect 209188 181540 209194 181552
rect 233326 181540 233332 181552
rect 209188 181512 233332 181540
rect 209188 181500 209194 181512
rect 233326 181500 233332 181512
rect 233384 181500 233390 181552
rect 235994 181500 236000 181552
rect 236052 181540 236058 181552
rect 274542 181540 274548 181552
rect 236052 181512 274548 181540
rect 236052 181500 236058 181512
rect 274542 181500 274548 181512
rect 274600 181500 274606 181552
rect 167638 181432 167644 181484
rect 167696 181472 167702 181484
rect 245746 181472 245752 181484
rect 167696 181444 245752 181472
rect 167696 181432 167702 181444
rect 245746 181432 245752 181444
rect 245804 181432 245810 181484
rect 269850 181432 269856 181484
rect 269908 181472 269914 181484
rect 298370 181472 298376 181484
rect 269908 181444 298376 181472
rect 269908 181432 269914 181444
rect 298370 181432 298376 181444
rect 298428 181432 298434 181484
rect 125962 180888 125968 180940
rect 126020 180928 126026 180940
rect 166442 180928 166448 180940
rect 126020 180900 166448 180928
rect 126020 180888 126026 180900
rect 166442 180888 166448 180900
rect 166500 180888 166506 180940
rect 148226 180820 148232 180872
rect 148284 180860 148290 180872
rect 209038 180860 209044 180872
rect 148284 180832 209044 180860
rect 148284 180820 148290 180832
rect 209038 180820 209044 180832
rect 209096 180820 209102 180872
rect 232498 180208 232504 180260
rect 232556 180248 232562 180260
rect 241698 180248 241704 180260
rect 232556 180220 241704 180248
rect 232556 180208 232562 180220
rect 241698 180208 241704 180220
rect 241756 180208 241762 180260
rect 214558 180140 214564 180192
rect 214616 180180 214622 180192
rect 233142 180180 233148 180192
rect 214616 180152 233148 180180
rect 214616 180140 214622 180152
rect 233142 180140 233148 180152
rect 233200 180140 233206 180192
rect 272518 180140 272524 180192
rect 272576 180180 272582 180192
rect 292850 180180 292856 180192
rect 272576 180152 292856 180180
rect 272576 180140 272582 180152
rect 292850 180140 292856 180152
rect 292908 180140 292914 180192
rect 169018 180072 169024 180124
rect 169076 180112 169082 180124
rect 224218 180112 224224 180124
rect 169076 180084 224224 180112
rect 169076 180072 169082 180084
rect 224218 180072 224224 180084
rect 224276 180072 224282 180124
rect 239398 180072 239404 180124
rect 239456 180112 239462 180124
rect 252646 180112 252652 180124
rect 239456 180084 252652 180112
rect 239456 180072 239462 180084
rect 252646 180072 252652 180084
rect 252704 180072 252710 180124
rect 257430 180072 257436 180124
rect 257488 180112 257494 180124
rect 288526 180112 288532 180124
rect 257488 180084 288532 180112
rect 257488 180072 257494 180084
rect 288526 180072 288532 180084
rect 288584 180072 288590 180124
rect 192478 179868 192484 179920
rect 192536 179908 192542 179920
rect 197998 179908 198004 179920
rect 192536 179880 198004 179908
rect 192536 179868 192542 179880
rect 197998 179868 198004 179880
rect 198056 179868 198062 179920
rect 129458 179460 129464 179512
rect 129516 179500 129522 179512
rect 165430 179500 165436 179512
rect 129516 179472 165436 179500
rect 129516 179460 129522 179472
rect 165430 179460 165436 179472
rect 165488 179460 165494 179512
rect 121914 179392 121920 179444
rect 121972 179432 121978 179444
rect 192570 179432 192576 179444
rect 121972 179404 192576 179432
rect 121972 179392 121978 179404
rect 192570 179392 192576 179404
rect 192628 179392 192634 179444
rect 224310 179392 224316 179444
rect 224368 179432 224374 179444
rect 229462 179432 229468 179444
rect 224368 179404 229468 179432
rect 224368 179392 224374 179404
rect 229462 179392 229468 179404
rect 229520 179392 229526 179444
rect 574738 179324 574744 179376
rect 574796 179364 574802 179376
rect 580166 179364 580172 179376
rect 574796 179336 580172 179364
rect 574796 179324 574802 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 224218 179256 224224 179308
rect 224276 179296 224282 179308
rect 229922 179296 229928 179308
rect 224276 179268 229928 179296
rect 224276 179256 224282 179268
rect 229922 179256 229928 179268
rect 229980 179256 229986 179308
rect 171962 178712 171968 178764
rect 172020 178752 172026 178764
rect 197354 178752 197360 178764
rect 172020 178724 197360 178752
rect 172020 178712 172026 178724
rect 197354 178712 197360 178724
rect 197412 178712 197418 178764
rect 278038 178712 278044 178764
rect 278096 178752 278102 178764
rect 294230 178752 294236 178764
rect 278096 178724 294236 178752
rect 278096 178712 278102 178724
rect 294230 178712 294236 178724
rect 294288 178712 294294 178764
rect 184290 178644 184296 178696
rect 184348 178684 184354 178696
rect 242894 178684 242900 178696
rect 184348 178656 242900 178684
rect 184348 178644 184354 178656
rect 242894 178644 242900 178656
rect 242952 178644 242958 178696
rect 243538 178644 243544 178696
rect 243596 178684 243602 178696
rect 287146 178684 287152 178696
rect 243596 178656 287152 178684
rect 243596 178644 243602 178656
rect 287146 178644 287152 178656
rect 287204 178644 287210 178696
rect 123294 178100 123300 178152
rect 123352 178140 123358 178152
rect 164970 178140 164976 178152
rect 123352 178112 164976 178140
rect 123352 178100 123358 178112
rect 164970 178100 164976 178112
rect 165028 178100 165034 178152
rect 115842 178032 115848 178084
rect 115900 178072 115906 178084
rect 171870 178072 171876 178084
rect 115900 178044 171876 178072
rect 115900 178032 115906 178044
rect 171870 178032 171876 178044
rect 171928 178032 171934 178084
rect 222838 177352 222844 177404
rect 222896 177392 222902 177404
rect 232130 177392 232136 177404
rect 222896 177364 232136 177392
rect 222896 177352 222902 177364
rect 232130 177352 232136 177364
rect 232188 177352 232194 177404
rect 271138 177352 271144 177404
rect 271196 177392 271202 177404
rect 285858 177392 285864 177404
rect 271196 177364 285864 177392
rect 271196 177352 271202 177364
rect 285858 177352 285864 177364
rect 285916 177352 285922 177404
rect 193858 177284 193864 177336
rect 193916 177324 193922 177336
rect 229370 177324 229376 177336
rect 193916 177296 229376 177324
rect 193916 177284 193922 177296
rect 229370 177284 229376 177296
rect 229428 177284 229434 177336
rect 231210 177284 231216 177336
rect 231268 177324 231274 177336
rect 238846 177324 238852 177336
rect 231268 177296 238852 177324
rect 231268 177284 231274 177296
rect 238846 177284 238852 177296
rect 238904 177284 238910 177336
rect 268378 177284 268384 177336
rect 268436 177324 268442 177336
rect 287238 177324 287244 177336
rect 268436 177296 287244 177324
rect 268436 177284 268442 177296
rect 287238 177284 287244 177296
rect 287296 177284 287302 177336
rect 128170 176808 128176 176860
rect 128228 176848 128234 176860
rect 207014 176848 207020 176860
rect 128228 176820 207020 176848
rect 128228 176808 128234 176820
rect 207014 176808 207020 176820
rect 207072 176808 207078 176860
rect 158990 176740 158996 176792
rect 159048 176780 159054 176792
rect 174722 176780 174728 176792
rect 159048 176752 174728 176780
rect 159048 176740 159054 176752
rect 174722 176740 174728 176752
rect 174780 176740 174786 176792
rect 67542 176672 67548 176724
rect 67600 176712 67606 176724
rect 70486 176712 70492 176724
rect 67600 176684 70492 176712
rect 67600 176672 67606 176684
rect 70486 176672 70492 176684
rect 70544 176672 70550 176724
rect 136082 176672 136088 176724
rect 136140 176712 136146 176724
rect 136140 176684 142154 176712
rect 136140 176672 136146 176684
rect 142126 176644 142154 176684
rect 213914 176644 213920 176656
rect 142126 176616 213920 176644
rect 213914 176604 213920 176616
rect 213972 176604 213978 176656
rect 164878 176196 164884 176248
rect 164936 176236 164942 176248
rect 166994 176236 167000 176248
rect 164936 176208 167000 176236
rect 164936 176196 164942 176208
rect 166994 176196 167000 176208
rect 167052 176196 167058 176248
rect 231118 176128 231124 176180
rect 231176 176168 231182 176180
rect 235994 176168 236000 176180
rect 231176 176140 236000 176168
rect 231176 176128 231182 176140
rect 235994 176128 236000 176140
rect 236052 176128 236058 176180
rect 220078 175992 220084 176044
rect 220136 176032 220142 176044
rect 231854 176032 231860 176044
rect 220136 176004 231860 176032
rect 220136 175992 220142 176004
rect 231854 175992 231860 176004
rect 231912 175992 231918 176044
rect 233142 175992 233148 176044
rect 233200 176032 233206 176044
rect 244366 176032 244372 176044
rect 233200 176004 244372 176032
rect 233200 175992 233206 176004
rect 244366 175992 244372 176004
rect 244424 175992 244430 176044
rect 276658 175992 276664 176044
rect 276716 176032 276722 176044
rect 284570 176032 284576 176044
rect 276716 176004 284576 176032
rect 276716 175992 276722 176004
rect 284570 175992 284576 176004
rect 284628 175992 284634 176044
rect 119430 175924 119436 175976
rect 119488 175964 119494 175976
rect 165062 175964 165068 175976
rect 119488 175936 165068 175964
rect 119488 175924 119494 175936
rect 165062 175924 165068 175936
rect 165120 175924 165126 175976
rect 207014 175924 207020 175976
rect 207072 175964 207078 175976
rect 214098 175964 214104 175976
rect 207072 175936 214104 175964
rect 207072 175924 207078 175936
rect 214098 175924 214104 175936
rect 214156 175924 214162 175976
rect 215202 175924 215208 175976
rect 215260 175964 215266 175976
rect 229186 175964 229192 175976
rect 215260 175936 229192 175964
rect 215260 175924 215266 175936
rect 229186 175924 229192 175936
rect 229244 175924 229250 175976
rect 246298 175924 246304 175976
rect 246356 175964 246362 175976
rect 278774 175964 278780 175976
rect 246356 175936 278780 175964
rect 246356 175924 246362 175936
rect 278774 175924 278780 175936
rect 278832 175924 278838 175976
rect 224954 175788 224960 175840
rect 225012 175788 225018 175840
rect 273346 175788 273352 175840
rect 273404 175788 273410 175840
rect 135254 175176 135260 175228
rect 135312 175216 135318 175228
rect 213914 175216 213920 175228
rect 135312 175188 213920 175216
rect 135312 175176 135318 175188
rect 213914 175176 213920 175188
rect 213972 175176 213978 175228
rect 224972 175216 225000 175788
rect 243630 175244 243636 175296
rect 243688 175284 243694 175296
rect 264974 175284 264980 175296
rect 243688 175256 264980 175284
rect 243688 175244 243694 175256
rect 264974 175244 264980 175256
rect 265032 175244 265038 175296
rect 229278 175216 229284 175228
rect 224972 175188 229284 175216
rect 229278 175176 229284 175188
rect 229336 175176 229342 175228
rect 229922 175176 229928 175228
rect 229980 175216 229986 175228
rect 230842 175216 230848 175228
rect 229980 175188 230848 175216
rect 229980 175176 229986 175188
rect 230842 175176 230848 175188
rect 230900 175176 230906 175228
rect 231118 175176 231124 175228
rect 231176 175216 231182 175228
rect 249886 175216 249892 175228
rect 231176 175188 249892 175216
rect 231176 175176 231182 175188
rect 249886 175176 249892 175188
rect 249944 175176 249950 175228
rect 273364 175216 273392 175788
rect 279418 175216 279424 175228
rect 273364 175188 279424 175216
rect 279418 175176 279424 175188
rect 279476 175176 279482 175228
rect 192662 175108 192668 175160
rect 192720 175148 192726 175160
rect 214006 175148 214012 175160
rect 192720 175120 214012 175148
rect 192720 175108 192726 175120
rect 214006 175108 214012 175120
rect 214064 175108 214070 175160
rect 263134 173952 263140 174004
rect 263192 173992 263198 174004
rect 264974 173992 264980 174004
rect 263192 173964 264980 173992
rect 263192 173952 263198 173964
rect 264974 173952 264980 173964
rect 265032 173952 265038 174004
rect 214558 173884 214564 173936
rect 214616 173924 214622 173936
rect 242986 173924 242992 173936
rect 214616 173896 242992 173924
rect 214616 173884 214622 173896
rect 242986 173884 242992 173896
rect 243044 173884 243050 173936
rect 245010 173884 245016 173936
rect 245068 173924 245074 173936
rect 265066 173924 265072 173936
rect 245068 173896 265072 173924
rect 245068 173884 245074 173896
rect 265066 173884 265072 173896
rect 265124 173884 265130 173936
rect 172054 173816 172060 173868
rect 172112 173856 172118 173868
rect 213914 173856 213920 173868
rect 172112 173828 213920 173856
rect 172112 173816 172118 173828
rect 213914 173816 213920 173828
rect 213972 173816 213978 173868
rect 231578 173816 231584 173868
rect 231636 173856 231642 173868
rect 239398 173856 239404 173868
rect 231636 173828 239404 173856
rect 231636 173816 231642 173828
rect 239398 173816 239404 173828
rect 239456 173816 239462 173868
rect 282454 173816 282460 173868
rect 282512 173856 282518 173868
rect 289906 173856 289912 173868
rect 282512 173828 289912 173856
rect 282512 173816 282518 173828
rect 289906 173816 289912 173828
rect 289964 173816 289970 173868
rect 188614 173748 188620 173800
rect 188672 173788 188678 173800
rect 214006 173788 214012 173800
rect 188672 173760 214012 173788
rect 188672 173748 188678 173760
rect 214006 173748 214012 173760
rect 214064 173748 214070 173800
rect 229094 173612 229100 173664
rect 229152 173652 229158 173664
rect 229462 173652 229468 173664
rect 229152 173624 229468 173652
rect 229152 173612 229158 173624
rect 229462 173612 229468 173624
rect 229520 173612 229526 173664
rect 250530 172592 250536 172644
rect 250588 172632 250594 172644
rect 264974 172632 264980 172644
rect 250588 172604 264980 172632
rect 250588 172592 250594 172604
rect 264974 172592 264980 172604
rect 265032 172592 265038 172644
rect 238202 172524 238208 172576
rect 238260 172564 238266 172576
rect 265066 172564 265072 172576
rect 238260 172536 265072 172564
rect 238260 172524 238266 172536
rect 265066 172524 265072 172536
rect 265124 172524 265130 172576
rect 165430 172456 165436 172508
rect 165488 172496 165494 172508
rect 213914 172496 213920 172508
rect 165488 172468 213920 172496
rect 165488 172456 165494 172468
rect 213914 172456 213920 172468
rect 213972 172456 213978 172508
rect 231578 172456 231584 172508
rect 231636 172496 231642 172508
rect 240226 172496 240232 172508
rect 231636 172468 240232 172496
rect 231636 172456 231642 172468
rect 240226 172456 240232 172468
rect 240284 172456 240290 172508
rect 282086 172456 282092 172508
rect 282144 172496 282150 172508
rect 295610 172496 295616 172508
rect 282144 172468 295616 172496
rect 282144 172456 282150 172468
rect 295610 172456 295616 172468
rect 295668 172456 295674 172508
rect 240226 171776 240232 171828
rect 240284 171816 240290 171828
rect 248414 171816 248420 171828
rect 240284 171788 248420 171816
rect 240284 171776 240290 171788
rect 248414 171776 248420 171788
rect 248472 171776 248478 171828
rect 258810 171232 258816 171284
rect 258868 171272 258874 171284
rect 264974 171272 264980 171284
rect 258868 171244 264980 171272
rect 258868 171232 258874 171244
rect 264974 171232 264980 171244
rect 265032 171232 265038 171284
rect 240778 171096 240784 171148
rect 240836 171136 240842 171148
rect 265066 171136 265072 171148
rect 240836 171108 265072 171136
rect 240836 171096 240842 171108
rect 265066 171096 265072 171108
rect 265124 171096 265130 171148
rect 166442 171028 166448 171080
rect 166500 171068 166506 171080
rect 214006 171068 214012 171080
rect 166500 171040 214012 171068
rect 166500 171028 166506 171040
rect 214006 171028 214012 171040
rect 214064 171028 214070 171080
rect 231118 171028 231124 171080
rect 231176 171068 231182 171080
rect 233510 171068 233516 171080
rect 231176 171040 233516 171068
rect 231176 171028 231182 171040
rect 233510 171028 233516 171040
rect 233568 171028 233574 171080
rect 282822 171028 282828 171080
rect 282880 171068 282886 171080
rect 298186 171068 298192 171080
rect 282880 171040 298192 171068
rect 282880 171028 282886 171040
rect 298186 171028 298192 171040
rect 298244 171028 298250 171080
rect 174630 170960 174636 171012
rect 174688 171000 174694 171012
rect 213914 171000 213920 171012
rect 174688 170972 213920 171000
rect 174688 170960 174694 170972
rect 213914 170960 213920 170972
rect 213972 170960 213978 171012
rect 236822 169804 236828 169856
rect 236880 169844 236886 169856
rect 264974 169844 264980 169856
rect 236880 169816 264980 169844
rect 236880 169804 236886 169816
rect 264974 169804 264980 169816
rect 265032 169804 265038 169856
rect 233970 169736 233976 169788
rect 234028 169776 234034 169788
rect 265066 169776 265072 169788
rect 234028 169748 265072 169776
rect 234028 169736 234034 169748
rect 265066 169736 265072 169748
rect 265124 169736 265130 169788
rect 164970 169668 164976 169720
rect 165028 169708 165034 169720
rect 214006 169708 214012 169720
rect 165028 169680 214012 169708
rect 165028 169668 165034 169680
rect 214006 169668 214012 169680
rect 214064 169668 214070 169720
rect 167822 169600 167828 169652
rect 167880 169640 167886 169652
rect 213914 169640 213920 169652
rect 167880 169612 213920 169640
rect 167880 169600 167886 169612
rect 213914 169600 213920 169612
rect 213972 169600 213978 169652
rect 281534 169464 281540 169516
rect 281592 169504 281598 169516
rect 283190 169504 283196 169516
rect 281592 169476 283196 169504
rect 281592 169464 281598 169476
rect 283190 169464 283196 169476
rect 283248 169464 283254 169516
rect 282822 169396 282828 169448
rect 282880 169436 282886 169448
rect 287330 169436 287336 169448
rect 282880 169408 287336 169436
rect 282880 169396 282886 169408
rect 287330 169396 287336 169408
rect 287388 169396 287394 169448
rect 238386 169056 238392 169108
rect 238444 169096 238450 169108
rect 241606 169096 241612 169108
rect 238444 169068 241612 169096
rect 238444 169056 238450 169068
rect 241606 169056 241612 169068
rect 241664 169056 241670 169108
rect 231670 168988 231676 169040
rect 231728 169028 231734 169040
rect 247034 169028 247040 169040
rect 231728 169000 247040 169028
rect 231728 168988 231734 169000
rect 247034 168988 247040 169000
rect 247092 168988 247098 169040
rect 247770 168444 247776 168496
rect 247828 168484 247834 168496
rect 264974 168484 264980 168496
rect 247828 168456 264980 168484
rect 247828 168444 247834 168456
rect 264974 168444 264980 168456
rect 265032 168444 265038 168496
rect 242250 168376 242256 168428
rect 242308 168416 242314 168428
rect 265066 168416 265072 168428
rect 242308 168388 265072 168416
rect 242308 168376 242314 168388
rect 265066 168376 265072 168388
rect 265124 168376 265130 168428
rect 192570 168308 192576 168360
rect 192628 168348 192634 168360
rect 213914 168348 213920 168360
rect 192628 168320 213920 168348
rect 192628 168308 192634 168320
rect 213914 168308 213920 168320
rect 213972 168308 213978 168360
rect 231762 168308 231768 168360
rect 231820 168348 231826 168360
rect 240226 168348 240232 168360
rect 231820 168320 240232 168348
rect 231820 168308 231826 168320
rect 240226 168308 240232 168320
rect 240284 168308 240290 168360
rect 282822 167696 282828 167748
rect 282880 167736 282886 167748
rect 288710 167736 288716 167748
rect 282880 167708 288716 167736
rect 282880 167696 282886 167708
rect 288710 167696 288716 167708
rect 288768 167696 288774 167748
rect 174722 167628 174728 167680
rect 174780 167668 174786 167680
rect 214558 167668 214564 167680
rect 174780 167640 214564 167668
rect 174780 167628 174786 167640
rect 214558 167628 214564 167640
rect 214616 167628 214622 167680
rect 229738 167628 229744 167680
rect 229796 167668 229802 167680
rect 239030 167668 239036 167680
rect 229796 167640 239036 167668
rect 229796 167628 229802 167640
rect 239030 167628 239036 167640
rect 239088 167628 239094 167680
rect 248046 167084 248052 167136
rect 248104 167124 248110 167136
rect 264974 167124 264980 167136
rect 248104 167096 264980 167124
rect 248104 167084 248110 167096
rect 264974 167084 264980 167096
rect 265032 167084 265038 167136
rect 239490 167016 239496 167068
rect 239548 167056 239554 167068
rect 265066 167056 265072 167068
rect 239548 167028 265072 167056
rect 239548 167016 239554 167028
rect 265066 167016 265072 167028
rect 265124 167016 265130 167068
rect 280062 167016 280068 167068
rect 280120 167056 280126 167068
rect 280430 167056 280436 167068
rect 280120 167028 280436 167056
rect 280120 167016 280126 167028
rect 280430 167016 280436 167028
rect 280488 167016 280494 167068
rect 165062 166948 165068 167000
rect 165120 166988 165126 167000
rect 213914 166988 213920 167000
rect 165120 166960 213920 166988
rect 165120 166948 165126 166960
rect 213914 166948 213920 166960
rect 213972 166948 213978 167000
rect 282822 166948 282828 167000
rect 282880 166988 282886 167000
rect 291378 166988 291384 167000
rect 282880 166960 291384 166988
rect 282880 166948 282886 166960
rect 291378 166948 291384 166960
rect 291436 166948 291442 167000
rect 170490 166880 170496 166932
rect 170548 166920 170554 166932
rect 214006 166920 214012 166932
rect 170548 166892 214012 166920
rect 170548 166880 170554 166892
rect 214006 166880 214012 166892
rect 214064 166880 214070 166932
rect 231762 166676 231768 166728
rect 231820 166716 231826 166728
rect 234890 166716 234896 166728
rect 231820 166688 234896 166716
rect 231820 166676 231826 166688
rect 234890 166676 234896 166688
rect 234948 166676 234954 166728
rect 230474 166268 230480 166320
rect 230532 166308 230538 166320
rect 230842 166308 230848 166320
rect 230532 166280 230848 166308
rect 230532 166268 230538 166280
rect 230842 166268 230848 166280
rect 230900 166268 230906 166320
rect 236086 166268 236092 166320
rect 236144 166308 236150 166320
rect 258074 166308 258080 166320
rect 236144 166280 258080 166308
rect 236144 166268 236150 166280
rect 258074 166268 258080 166280
rect 258132 166268 258138 166320
rect 262858 165656 262864 165708
rect 262916 165696 262922 165708
rect 265342 165696 265348 165708
rect 262916 165668 265348 165696
rect 262916 165656 262922 165668
rect 265342 165656 265348 165668
rect 265400 165656 265406 165708
rect 232774 165588 232780 165640
rect 232832 165628 232838 165640
rect 264974 165628 264980 165640
rect 232832 165600 264980 165628
rect 232832 165588 232838 165600
rect 264974 165588 264980 165600
rect 265032 165588 265038 165640
rect 166534 165520 166540 165572
rect 166592 165560 166598 165572
rect 214006 165560 214012 165572
rect 166592 165532 214012 165560
rect 166592 165520 166598 165532
rect 214006 165520 214012 165532
rect 214064 165520 214070 165572
rect 231486 165520 231492 165572
rect 231544 165560 231550 165572
rect 244366 165560 244372 165572
rect 231544 165532 244372 165560
rect 231544 165520 231550 165532
rect 244366 165520 244372 165532
rect 244424 165520 244430 165572
rect 281994 165520 282000 165572
rect 282052 165560 282058 165572
rect 284570 165560 284576 165572
rect 282052 165532 284576 165560
rect 282052 165520 282058 165532
rect 284570 165520 284576 165532
rect 284628 165520 284634 165572
rect 171870 165452 171876 165504
rect 171928 165492 171934 165504
rect 213914 165492 213920 165504
rect 171928 165464 213920 165492
rect 171928 165452 171934 165464
rect 213914 165452 213920 165464
rect 213972 165452 213978 165504
rect 231118 164840 231124 164892
rect 231176 164880 231182 164892
rect 248506 164880 248512 164892
rect 231176 164852 248512 164880
rect 231176 164840 231182 164852
rect 248506 164840 248512 164852
rect 248564 164840 248570 164892
rect 257614 164296 257620 164348
rect 257672 164336 257678 164348
rect 265066 164336 265072 164348
rect 257672 164308 265072 164336
rect 257672 164296 257678 164308
rect 265066 164296 265072 164308
rect 265124 164296 265130 164348
rect 251818 164228 251824 164280
rect 251876 164268 251882 164280
rect 264974 164268 264980 164280
rect 251876 164240 264980 164268
rect 251876 164228 251882 164240
rect 264974 164228 264980 164240
rect 265032 164228 265038 164280
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 25498 164200 25504 164212
rect 3292 164172 25504 164200
rect 3292 164160 3298 164172
rect 25498 164160 25504 164172
rect 25556 164160 25562 164212
rect 169202 164160 169208 164212
rect 169260 164200 169266 164212
rect 213914 164200 213920 164212
rect 169260 164172 213920 164200
rect 169260 164160 169266 164172
rect 213914 164160 213920 164172
rect 213972 164160 213978 164212
rect 282822 164160 282828 164212
rect 282880 164200 282886 164212
rect 303798 164200 303804 164212
rect 282880 164172 303804 164200
rect 282880 164160 282886 164172
rect 303798 164160 303804 164172
rect 303856 164160 303862 164212
rect 170582 164092 170588 164144
rect 170640 164132 170646 164144
rect 214006 164132 214012 164144
rect 170640 164104 214012 164132
rect 170640 164092 170646 164104
rect 214006 164092 214012 164104
rect 214064 164092 214070 164144
rect 282454 164092 282460 164144
rect 282512 164132 282518 164144
rect 285950 164132 285956 164144
rect 282512 164104 285956 164132
rect 282512 164092 282518 164104
rect 285950 164092 285956 164104
rect 286008 164092 286014 164144
rect 231762 163956 231768 164008
rect 231820 163996 231826 164008
rect 236086 163996 236092 164008
rect 231820 163968 236092 163996
rect 231820 163956 231826 163968
rect 236086 163956 236092 163968
rect 236144 163956 236150 164008
rect 250622 162936 250628 162988
rect 250680 162976 250686 162988
rect 264974 162976 264980 162988
rect 250680 162948 264980 162976
rect 250680 162936 250686 162948
rect 264974 162936 264980 162948
rect 265032 162936 265038 162988
rect 235534 162868 235540 162920
rect 235592 162908 235598 162920
rect 265066 162908 265072 162920
rect 235592 162880 265072 162908
rect 235592 162868 235598 162880
rect 265066 162868 265072 162880
rect 265124 162868 265130 162920
rect 173250 162800 173256 162852
rect 173308 162840 173314 162852
rect 214006 162840 214012 162852
rect 173308 162812 214012 162840
rect 173308 162800 173314 162812
rect 214006 162800 214012 162812
rect 214064 162800 214070 162852
rect 282822 162800 282828 162852
rect 282880 162840 282886 162852
rect 292758 162840 292764 162852
rect 282880 162812 292764 162840
rect 282880 162800 282886 162812
rect 292758 162800 292764 162812
rect 292816 162800 292822 162852
rect 177390 162732 177396 162784
rect 177448 162772 177454 162784
rect 213914 162772 213920 162784
rect 177448 162744 213920 162772
rect 177448 162732 177454 162744
rect 213914 162732 213920 162744
rect 213972 162732 213978 162784
rect 231302 162528 231308 162580
rect 231360 162568 231366 162580
rect 237558 162568 237564 162580
rect 231360 162540 237564 162568
rect 231360 162528 231366 162540
rect 237558 162528 237564 162540
rect 237616 162528 237622 162580
rect 236730 162120 236736 162172
rect 236788 162160 236794 162172
rect 265158 162160 265164 162172
rect 236788 162132 265164 162160
rect 236788 162120 236794 162132
rect 265158 162120 265164 162132
rect 265216 162120 265222 162172
rect 254578 161440 254584 161492
rect 254636 161480 254642 161492
rect 264974 161480 264980 161492
rect 254636 161452 264980 161480
rect 254636 161440 254642 161452
rect 264974 161440 264980 161452
rect 265032 161440 265038 161492
rect 169018 161372 169024 161424
rect 169076 161412 169082 161424
rect 214006 161412 214012 161424
rect 169076 161384 214012 161412
rect 169076 161372 169082 161384
rect 214006 161372 214012 161384
rect 214064 161372 214070 161424
rect 231762 161372 231768 161424
rect 231820 161412 231826 161424
rect 242986 161412 242992 161424
rect 231820 161384 242992 161412
rect 231820 161372 231826 161384
rect 242986 161372 242992 161384
rect 243044 161372 243050 161424
rect 195330 161304 195336 161356
rect 195388 161344 195394 161356
rect 213914 161344 213920 161356
rect 195388 161316 213920 161344
rect 195388 161304 195394 161316
rect 213914 161304 213920 161316
rect 213972 161304 213978 161356
rect 230934 160964 230940 161016
rect 230992 161004 230998 161016
rect 233234 161004 233240 161016
rect 230992 160976 233240 161004
rect 230992 160964 230998 160976
rect 233234 160964 233240 160976
rect 233292 160964 233298 161016
rect 245286 160692 245292 160744
rect 245344 160732 245350 160744
rect 262858 160732 262864 160744
rect 245344 160704 262864 160732
rect 245344 160692 245350 160704
rect 262858 160692 262864 160704
rect 262916 160692 262922 160744
rect 281534 160216 281540 160268
rect 281592 160256 281598 160268
rect 281810 160256 281816 160268
rect 281592 160228 281816 160256
rect 281592 160216 281598 160228
rect 281810 160216 281816 160228
rect 281868 160216 281874 160268
rect 282822 160148 282828 160200
rect 282880 160188 282886 160200
rect 288618 160188 288624 160200
rect 282880 160160 288624 160188
rect 282880 160148 282886 160160
rect 288618 160148 288624 160160
rect 288676 160148 288682 160200
rect 238018 160080 238024 160132
rect 238076 160120 238082 160132
rect 264974 160120 264980 160132
rect 238076 160092 264980 160120
rect 238076 160080 238082 160092
rect 264974 160080 264980 160092
rect 265032 160080 265038 160132
rect 182910 160012 182916 160064
rect 182968 160052 182974 160064
rect 213914 160052 213920 160064
rect 182968 160024 213920 160052
rect 182968 160012 182974 160024
rect 213914 160012 213920 160024
rect 213972 160012 213978 160064
rect 231762 160012 231768 160064
rect 231820 160052 231826 160064
rect 241698 160052 241704 160064
rect 231820 160024 241704 160052
rect 231820 160012 231826 160024
rect 241698 160012 241704 160024
rect 241756 160012 241762 160064
rect 281902 160012 281908 160064
rect 281960 160052 281966 160064
rect 294230 160052 294236 160064
rect 281960 160024 294236 160052
rect 281960 160012 281966 160024
rect 294230 160012 294236 160024
rect 294288 160012 294294 160064
rect 198090 159944 198096 159996
rect 198148 159984 198154 159996
rect 214006 159984 214012 159996
rect 198148 159956 214012 159984
rect 198148 159944 198154 159956
rect 214006 159944 214012 159956
rect 214064 159944 214070 159996
rect 282362 159944 282368 159996
rect 282420 159984 282426 159996
rect 290090 159984 290096 159996
rect 282420 159956 290096 159984
rect 282420 159944 282426 159956
rect 290090 159944 290096 159956
rect 290148 159944 290154 159996
rect 243906 158788 243912 158840
rect 243964 158828 243970 158840
rect 265066 158828 265072 158840
rect 243964 158800 265072 158828
rect 243964 158788 243970 158800
rect 265066 158788 265072 158800
rect 265124 158788 265130 158840
rect 233878 158720 233884 158772
rect 233936 158760 233942 158772
rect 264974 158760 264980 158772
rect 233936 158732 264980 158760
rect 233936 158720 233942 158732
rect 264974 158720 264980 158732
rect 265032 158720 265038 158772
rect 167730 158652 167736 158704
rect 167788 158692 167794 158704
rect 214006 158692 214012 158704
rect 167788 158664 214012 158692
rect 167788 158652 167794 158664
rect 214006 158652 214012 158664
rect 214064 158652 214070 158704
rect 282086 158652 282092 158704
rect 282144 158692 282150 158704
rect 300946 158692 300952 158704
rect 282144 158664 300952 158692
rect 282144 158652 282150 158664
rect 300946 158652 300952 158664
rect 301004 158652 301010 158704
rect 181530 158584 181536 158636
rect 181588 158624 181594 158636
rect 213914 158624 213920 158636
rect 181588 158596 213920 158624
rect 181588 158584 181594 158596
rect 213914 158584 213920 158596
rect 213972 158584 213978 158636
rect 231210 158584 231216 158636
rect 231268 158624 231274 158636
rect 240134 158624 240140 158636
rect 231268 158596 240140 158624
rect 231268 158584 231274 158596
rect 240134 158584 240140 158596
rect 240192 158584 240198 158636
rect 241146 157428 241152 157480
rect 241204 157468 241210 157480
rect 265066 157468 265072 157480
rect 241204 157440 265072 157468
rect 241204 157428 241210 157440
rect 265066 157428 265072 157440
rect 265124 157428 265130 157480
rect 235258 157360 235264 157412
rect 235316 157400 235322 157412
rect 264974 157400 264980 157412
rect 235316 157372 264980 157400
rect 235316 157360 235322 157372
rect 264974 157360 264980 157372
rect 265032 157360 265038 157412
rect 166350 157292 166356 157344
rect 166408 157332 166414 157344
rect 213914 157332 213920 157344
rect 166408 157304 213920 157332
rect 166408 157292 166414 157304
rect 213914 157292 213920 157304
rect 213972 157292 213978 157344
rect 180242 157224 180248 157276
rect 180300 157264 180306 157276
rect 214006 157264 214012 157276
rect 180300 157236 214012 157264
rect 180300 157224 180306 157236
rect 214006 157224 214012 157236
rect 214064 157224 214070 157276
rect 230934 156952 230940 157004
rect 230992 156992 230998 157004
rect 233418 156992 233424 157004
rect 230992 156964 233424 156992
rect 230992 156952 230998 156964
rect 233418 156952 233424 156964
rect 233476 156952 233482 157004
rect 236638 156612 236644 156664
rect 236696 156652 236702 156664
rect 265250 156652 265256 156664
rect 236696 156624 265256 156652
rect 236696 156612 236702 156624
rect 265250 156612 265256 156624
rect 265308 156612 265314 156664
rect 242434 155932 242440 155984
rect 242492 155972 242498 155984
rect 264974 155972 264980 155984
rect 242492 155944 264980 155972
rect 242492 155932 242498 155944
rect 264974 155932 264980 155944
rect 265032 155932 265038 155984
rect 178954 155864 178960 155916
rect 179012 155904 179018 155916
rect 213914 155904 213920 155916
rect 179012 155876 213920 155904
rect 179012 155864 179018 155876
rect 213914 155864 213920 155876
rect 213972 155864 213978 155916
rect 230842 155864 230848 155916
rect 230900 155904 230906 155916
rect 235994 155904 236000 155916
rect 230900 155876 236000 155904
rect 230900 155864 230906 155876
rect 235994 155864 236000 155876
rect 236052 155864 236058 155916
rect 282270 155864 282276 155916
rect 282328 155904 282334 155916
rect 310606 155904 310612 155916
rect 282328 155876 310612 155904
rect 282328 155864 282334 155876
rect 310606 155864 310612 155876
rect 310664 155864 310670 155916
rect 185762 155796 185768 155848
rect 185820 155836 185826 155848
rect 214006 155836 214012 155848
rect 185820 155808 214012 155836
rect 185820 155796 185826 155808
rect 214006 155796 214012 155808
rect 214064 155796 214070 155848
rect 246574 154640 246580 154692
rect 246632 154680 246638 154692
rect 265066 154680 265072 154692
rect 246632 154652 265072 154680
rect 246632 154640 246638 154652
rect 265066 154640 265072 154652
rect 265124 154640 265130 154692
rect 241054 154572 241060 154624
rect 241112 154612 241118 154624
rect 264974 154612 264980 154624
rect 241112 154584 264980 154612
rect 241112 154572 241118 154584
rect 264974 154572 264980 154584
rect 265032 154572 265038 154624
rect 282270 154504 282276 154556
rect 282328 154544 282334 154556
rect 302510 154544 302516 154556
rect 282328 154516 302516 154544
rect 282328 154504 282334 154516
rect 302510 154504 302516 154516
rect 302568 154504 302574 154556
rect 282822 154436 282828 154488
rect 282880 154476 282886 154488
rect 292850 154476 292856 154488
rect 282880 154448 292856 154476
rect 282880 154436 282886 154448
rect 292850 154436 292856 154448
rect 292908 154436 292914 154488
rect 231302 154368 231308 154420
rect 231360 154408 231366 154420
rect 237374 154408 237380 154420
rect 231360 154380 237380 154408
rect 231360 154368 231366 154380
rect 237374 154368 237380 154380
rect 237432 154368 237438 154420
rect 234154 153824 234160 153876
rect 234212 153864 234218 153876
rect 265710 153864 265716 153876
rect 234212 153836 265716 153864
rect 234212 153824 234218 153836
rect 265710 153824 265716 153836
rect 265768 153824 265774 153876
rect 192570 153280 192576 153332
rect 192628 153320 192634 153332
rect 213914 153320 213920 153332
rect 192628 153292 213920 153320
rect 192628 153280 192634 153292
rect 213914 153280 213920 153292
rect 213972 153280 213978 153332
rect 185670 153212 185676 153264
rect 185728 153252 185734 153264
rect 214006 153252 214012 153264
rect 185728 153224 214012 153252
rect 185728 153212 185734 153224
rect 214006 153212 214012 153224
rect 214064 153212 214070 153264
rect 262950 153212 262956 153264
rect 263008 153252 263014 153264
rect 265342 153252 265348 153264
rect 263008 153224 265348 153252
rect 263008 153212 263014 153224
rect 265342 153212 265348 153224
rect 265400 153212 265406 153264
rect 230474 153144 230480 153196
rect 230532 153184 230538 153196
rect 234614 153184 234620 153196
rect 230532 153156 234620 153184
rect 230532 153144 230538 153156
rect 234614 153144 234620 153156
rect 234672 153144 234678 153196
rect 167638 152464 167644 152516
rect 167696 152504 167702 152516
rect 194502 152504 194508 152516
rect 167696 152476 194508 152504
rect 167696 152464 167702 152476
rect 194502 152464 194508 152476
rect 194560 152464 194566 152516
rect 242158 151852 242164 151904
rect 242216 151892 242222 151904
rect 264974 151892 264980 151904
rect 242216 151864 264980 151892
rect 242216 151852 242222 151864
rect 264974 151852 264980 151864
rect 265032 151852 265038 151904
rect 206278 151784 206284 151836
rect 206336 151824 206342 151836
rect 213914 151824 213920 151836
rect 206336 151796 213920 151824
rect 206336 151784 206342 151796
rect 213914 151784 213920 151796
rect 213972 151784 213978 151836
rect 238110 151784 238116 151836
rect 238168 151824 238174 151836
rect 265066 151824 265072 151836
rect 238168 151796 265072 151824
rect 238168 151784 238174 151796
rect 265066 151784 265072 151796
rect 265124 151784 265130 151836
rect 281902 151716 281908 151768
rect 281960 151756 281966 151768
rect 307846 151756 307852 151768
rect 281960 151728 307852 151756
rect 281960 151716 281966 151728
rect 307846 151716 307852 151728
rect 307904 151716 307910 151768
rect 231578 151104 231584 151156
rect 231636 151144 231642 151156
rect 251266 151144 251272 151156
rect 231636 151116 251272 151144
rect 231636 151104 231642 151116
rect 251266 151104 251272 151116
rect 251324 151104 251330 151156
rect 232866 151036 232872 151088
rect 232924 151076 232930 151088
rect 265618 151076 265624 151088
rect 232924 151048 265624 151076
rect 232924 151036 232930 151048
rect 265618 151036 265624 151048
rect 265676 151036 265682 151088
rect 206370 150492 206376 150544
rect 206428 150532 206434 150544
rect 213914 150532 213920 150544
rect 206428 150504 213920 150532
rect 206428 150492 206434 150504
rect 213914 150492 213920 150504
rect 213972 150492 213978 150544
rect 183002 150424 183008 150476
rect 183060 150464 183066 150476
rect 214098 150464 214104 150476
rect 183060 150436 214104 150464
rect 183060 150424 183066 150436
rect 214098 150424 214104 150436
rect 214156 150424 214162 150476
rect 261478 150424 261484 150476
rect 261536 150464 261542 150476
rect 264974 150464 264980 150476
rect 261536 150436 264980 150464
rect 261536 150424 261542 150436
rect 264974 150424 264980 150436
rect 265032 150424 265038 150476
rect 194502 150356 194508 150408
rect 194560 150396 194566 150408
rect 214006 150396 214012 150408
rect 194560 150368 214012 150396
rect 194560 150356 194566 150368
rect 214006 150356 214012 150368
rect 214064 150356 214070 150408
rect 230566 150356 230572 150408
rect 230624 150396 230630 150408
rect 241514 150396 241520 150408
rect 230624 150368 241520 150396
rect 230624 150356 230630 150368
rect 241514 150356 241520 150368
rect 241572 150356 241578 150408
rect 2774 150288 2780 150340
rect 2832 150328 2838 150340
rect 4798 150328 4804 150340
rect 2832 150300 4804 150328
rect 2832 150288 2838 150300
rect 4798 150288 4804 150300
rect 4856 150288 4862 150340
rect 209038 150288 209044 150340
rect 209096 150328 209102 150340
rect 213914 150328 213920 150340
rect 209096 150300 213920 150328
rect 209096 150288 209102 150300
rect 213914 150288 213920 150300
rect 213972 150288 213978 150340
rect 249242 149676 249248 149728
rect 249300 149716 249306 149728
rect 265158 149716 265164 149728
rect 249300 149688 265164 149716
rect 249300 149676 249306 149688
rect 265158 149676 265164 149688
rect 265216 149676 265222 149728
rect 256050 149064 256056 149116
rect 256108 149104 256114 149116
rect 264974 149104 264980 149116
rect 256108 149076 264980 149104
rect 256108 149064 256114 149076
rect 264974 149064 264980 149076
rect 265032 149064 265038 149116
rect 231762 148996 231768 149048
rect 231820 149036 231826 149048
rect 247218 149036 247224 149048
rect 231820 149008 247224 149036
rect 231820 148996 231826 149008
rect 247218 148996 247224 149008
rect 247276 148996 247282 149048
rect 282822 148996 282828 149048
rect 282880 149036 282886 149048
rect 306558 149036 306564 149048
rect 282880 149008 306564 149036
rect 282880 148996 282886 149008
rect 306558 148996 306564 149008
rect 306616 148996 306622 149048
rect 234062 148316 234068 148368
rect 234120 148356 234126 148368
rect 265250 148356 265256 148368
rect 234120 148328 265256 148356
rect 234120 148316 234126 148328
rect 265250 148316 265256 148328
rect 265308 148316 265314 148368
rect 282638 147840 282644 147892
rect 282696 147880 282702 147892
rect 287238 147880 287244 147892
rect 282696 147852 287244 147880
rect 282696 147840 282702 147852
rect 287238 147840 287244 147852
rect 287296 147840 287302 147892
rect 166350 147636 166356 147688
rect 166408 147676 166414 147688
rect 213914 147676 213920 147688
rect 166408 147648 213920 147676
rect 166408 147636 166414 147648
rect 213914 147636 213920 147648
rect 213972 147636 213978 147688
rect 259086 147636 259092 147688
rect 259144 147676 259150 147688
rect 264974 147676 264980 147688
rect 259144 147648 264980 147676
rect 259144 147636 259150 147648
rect 264974 147636 264980 147648
rect 265032 147636 265038 147688
rect 282822 147568 282828 147620
rect 282880 147608 282886 147620
rect 305178 147608 305184 147620
rect 282880 147580 305184 147608
rect 282880 147568 282886 147580
rect 305178 147568 305184 147580
rect 305236 147568 305242 147620
rect 282270 147500 282276 147552
rect 282328 147540 282334 147552
rect 298278 147540 298284 147552
rect 282328 147512 298284 147540
rect 282328 147500 282334 147512
rect 298278 147500 298284 147512
rect 298336 147500 298342 147552
rect 239674 146888 239680 146940
rect 239732 146928 239738 146940
rect 265066 146928 265072 146940
rect 239732 146900 265072 146928
rect 239732 146888 239738 146900
rect 265066 146888 265072 146900
rect 265124 146888 265130 146940
rect 231118 146820 231124 146872
rect 231176 146860 231182 146872
rect 236822 146860 236828 146872
rect 231176 146832 236828 146860
rect 231176 146820 231182 146832
rect 236822 146820 236828 146832
rect 236880 146820 236886 146872
rect 231302 146548 231308 146600
rect 231360 146588 231366 146600
rect 238202 146588 238208 146600
rect 231360 146560 238208 146588
rect 231360 146548 231366 146560
rect 238202 146548 238208 146560
rect 238260 146548 238266 146600
rect 184382 146276 184388 146328
rect 184440 146316 184446 146328
rect 213914 146316 213920 146328
rect 184440 146288 213920 146316
rect 184440 146276 184446 146288
rect 213914 146276 213920 146288
rect 213972 146276 213978 146328
rect 247954 146276 247960 146328
rect 248012 146316 248018 146328
rect 264974 146316 264980 146328
rect 248012 146288 264980 146316
rect 248012 146276 248018 146288
rect 264974 146276 264980 146288
rect 265032 146276 265038 146328
rect 282822 146208 282828 146260
rect 282880 146248 282886 146260
rect 313274 146248 313280 146260
rect 282880 146220 313280 146248
rect 282880 146208 282886 146220
rect 313274 146208 313280 146220
rect 313332 146208 313338 146260
rect 282730 146140 282736 146192
rect 282788 146180 282794 146192
rect 294138 146180 294144 146192
rect 282788 146152 294144 146180
rect 282788 146140 282794 146152
rect 294138 146140 294144 146152
rect 294196 146140 294202 146192
rect 231210 145528 231216 145580
rect 231268 145568 231274 145580
rect 240778 145568 240784 145580
rect 231268 145540 240784 145568
rect 231268 145528 231274 145540
rect 240778 145528 240784 145540
rect 240836 145528 240842 145580
rect 198182 144984 198188 145036
rect 198240 145024 198246 145036
rect 214006 145024 214012 145036
rect 198240 144996 214012 145024
rect 198240 144984 198246 144996
rect 214006 144984 214012 144996
rect 214064 144984 214070 145036
rect 240962 144984 240968 145036
rect 241020 145024 241026 145036
rect 264974 145024 264980 145036
rect 241020 144996 264980 145024
rect 241020 144984 241026 144996
rect 264974 144984 264980 144996
rect 265032 144984 265038 145036
rect 169018 144916 169024 144968
rect 169076 144956 169082 144968
rect 213914 144956 213920 144968
rect 169076 144928 213920 144956
rect 169076 144916 169082 144928
rect 213914 144916 213920 144928
rect 213972 144916 213978 144968
rect 235350 144916 235356 144968
rect 235408 144956 235414 144968
rect 265066 144956 265072 144968
rect 235408 144928 265072 144956
rect 235408 144916 235414 144928
rect 265066 144916 265072 144928
rect 265124 144916 265130 144968
rect 282822 144848 282828 144900
rect 282880 144888 282886 144900
rect 299750 144888 299756 144900
rect 282880 144860 299756 144888
rect 282880 144848 282886 144860
rect 299750 144848 299756 144860
rect 299808 144848 299814 144900
rect 173158 144168 173164 144220
rect 173216 144208 173222 144220
rect 184290 144208 184296 144220
rect 173216 144180 184296 144208
rect 173216 144168 173222 144180
rect 184290 144168 184296 144180
rect 184348 144168 184354 144220
rect 230566 144168 230572 144220
rect 230624 144208 230630 144220
rect 249058 144208 249064 144220
rect 230624 144180 249064 144208
rect 230624 144168 230630 144180
rect 249058 144168 249064 144180
rect 249116 144168 249122 144220
rect 231762 144032 231768 144084
rect 231820 144072 231826 144084
rect 238386 144072 238392 144084
rect 231820 144044 238392 144072
rect 231820 144032 231826 144044
rect 238386 144032 238392 144044
rect 238444 144032 238450 144084
rect 202230 143624 202236 143676
rect 202288 143664 202294 143676
rect 214006 143664 214012 143676
rect 202288 143636 214012 143664
rect 202288 143624 202294 143636
rect 214006 143624 214012 143636
rect 214064 143624 214070 143676
rect 250806 143624 250812 143676
rect 250864 143664 250870 143676
rect 265066 143664 265072 143676
rect 250864 143636 265072 143664
rect 250864 143624 250870 143636
rect 265066 143624 265072 143636
rect 265124 143624 265130 143676
rect 189810 143556 189816 143608
rect 189868 143596 189874 143608
rect 213914 143596 213920 143608
rect 189868 143568 213920 143596
rect 189868 143556 189874 143568
rect 213914 143556 213920 143568
rect 213972 143556 213978 143608
rect 242342 143556 242348 143608
rect 242400 143596 242406 143608
rect 264974 143596 264980 143608
rect 242400 143568 264980 143596
rect 242400 143556 242406 143568
rect 264974 143556 264980 143568
rect 265032 143556 265038 143608
rect 231762 143488 231768 143540
rect 231820 143528 231826 143540
rect 243814 143528 243820 143540
rect 231820 143500 243820 143528
rect 231820 143488 231826 143500
rect 243814 143488 243820 143500
rect 243872 143488 243878 143540
rect 282822 143488 282828 143540
rect 282880 143528 282886 143540
rect 295334 143528 295340 143540
rect 282880 143500 295340 143528
rect 282880 143488 282886 143500
rect 295334 143488 295340 143500
rect 295392 143488 295398 143540
rect 171778 142808 171784 142860
rect 171836 142848 171842 142860
rect 193858 142848 193864 142860
rect 171836 142820 193864 142848
rect 171836 142808 171842 142820
rect 193858 142808 193864 142820
rect 193916 142808 193922 142860
rect 209222 142196 209228 142248
rect 209280 142236 209286 142248
rect 213914 142236 213920 142248
rect 209280 142208 213920 142236
rect 209280 142196 209286 142208
rect 213914 142196 213920 142208
rect 213972 142196 213978 142248
rect 254762 142196 254768 142248
rect 254820 142236 254826 142248
rect 265066 142236 265072 142248
rect 254820 142208 265072 142236
rect 254820 142196 254826 142208
rect 265066 142196 265072 142208
rect 265124 142196 265130 142248
rect 180334 142128 180340 142180
rect 180392 142168 180398 142180
rect 214006 142168 214012 142180
rect 180392 142140 214012 142168
rect 180392 142128 180398 142140
rect 214006 142128 214012 142140
rect 214064 142128 214070 142180
rect 238202 142128 238208 142180
rect 238260 142168 238266 142180
rect 264974 142168 264980 142180
rect 238260 142140 264980 142168
rect 238260 142128 238266 142140
rect 264974 142128 264980 142140
rect 265032 142128 265038 142180
rect 282546 142060 282552 142112
rect 282604 142100 282610 142112
rect 285858 142100 285864 142112
rect 282604 142072 285864 142100
rect 282604 142060 282610 142072
rect 285858 142060 285864 142072
rect 285916 142060 285922 142112
rect 169110 141380 169116 141432
rect 169168 141420 169174 141432
rect 209038 141420 209044 141432
rect 169168 141392 209044 141420
rect 169168 141380 169174 141392
rect 209038 141380 209044 141392
rect 209096 141380 209102 141432
rect 230934 141380 230940 141432
rect 230992 141420 230998 141432
rect 263134 141420 263140 141432
rect 230992 141392 263140 141420
rect 230992 141380 230998 141392
rect 263134 141380 263140 141392
rect 263192 141380 263198 141432
rect 282822 141312 282828 141364
rect 282880 141352 282886 141364
rect 288434 141352 288440 141364
rect 282880 141324 288440 141352
rect 282880 141312 282886 141324
rect 288434 141312 288440 141324
rect 288492 141312 288498 141364
rect 263042 140836 263048 140888
rect 263100 140876 263106 140888
rect 265250 140876 265256 140888
rect 263100 140848 265256 140876
rect 263100 140836 263106 140848
rect 265250 140836 265256 140848
rect 265308 140836 265314 140888
rect 180242 140768 180248 140820
rect 180300 140808 180306 140820
rect 213914 140808 213920 140820
rect 180300 140780 213920 140808
rect 180300 140768 180306 140780
rect 213914 140768 213920 140780
rect 213972 140768 213978 140820
rect 236822 140768 236828 140820
rect 236880 140808 236886 140820
rect 264974 140808 264980 140820
rect 236880 140780 264980 140808
rect 236880 140768 236886 140780
rect 264974 140768 264980 140780
rect 265032 140768 265038 140820
rect 231762 140700 231768 140752
rect 231820 140740 231826 140752
rect 245746 140740 245752 140752
rect 231820 140712 245752 140740
rect 231820 140700 231826 140712
rect 245746 140700 245752 140712
rect 245804 140700 245810 140752
rect 282822 140700 282828 140752
rect 282880 140740 282886 140752
rect 291470 140740 291476 140752
rect 282880 140712 291476 140740
rect 282880 140700 282886 140712
rect 291470 140700 291476 140712
rect 291528 140700 291534 140752
rect 180150 140020 180156 140072
rect 180208 140060 180214 140072
rect 199378 140060 199384 140072
rect 180208 140032 199384 140060
rect 180208 140020 180214 140032
rect 199378 140020 199384 140032
rect 199436 140020 199442 140072
rect 240778 140020 240784 140072
rect 240836 140060 240842 140072
rect 263226 140060 263232 140072
rect 240836 140032 263232 140060
rect 240836 140020 240842 140032
rect 263226 140020 263232 140032
rect 263284 140020 263290 140072
rect 210602 139476 210608 139528
rect 210660 139516 210666 139528
rect 214098 139516 214104 139528
rect 210660 139488 214104 139516
rect 210660 139476 210666 139488
rect 214098 139476 214104 139488
rect 214156 139476 214162 139528
rect 258994 139476 259000 139528
rect 259052 139516 259058 139528
rect 265158 139516 265164 139528
rect 259052 139488 265164 139516
rect 259052 139476 259058 139488
rect 265158 139476 265164 139488
rect 265216 139476 265222 139528
rect 211798 139408 211804 139460
rect 211856 139448 211862 139460
rect 213914 139448 213920 139460
rect 211856 139420 213920 139448
rect 211856 139408 211862 139420
rect 213914 139408 213920 139420
rect 213972 139408 213978 139460
rect 263134 139408 263140 139460
rect 263192 139448 263198 139460
rect 264974 139448 264980 139460
rect 263192 139420 264980 139448
rect 263192 139408 263198 139420
rect 264974 139408 264980 139420
rect 265032 139408 265038 139460
rect 177298 138660 177304 138712
rect 177356 138700 177362 138712
rect 200850 138700 200856 138712
rect 177356 138672 200856 138700
rect 177356 138660 177362 138672
rect 200850 138660 200856 138672
rect 200908 138660 200914 138712
rect 229922 138660 229928 138712
rect 229980 138700 229986 138712
rect 264974 138700 264980 138712
rect 229980 138672 264980 138700
rect 229980 138660 229986 138672
rect 264974 138660 264980 138672
rect 265032 138660 265038 138712
rect 281534 138320 281540 138372
rect 281592 138360 281598 138372
rect 284478 138360 284484 138372
rect 281592 138332 284484 138360
rect 281592 138320 281598 138332
rect 284478 138320 284484 138332
rect 284536 138320 284542 138372
rect 192478 137980 192484 138032
rect 192536 138020 192542 138032
rect 213914 138020 213920 138032
rect 192536 137992 213920 138020
rect 192536 137980 192542 137992
rect 213914 137980 213920 137992
rect 213972 137980 213978 138032
rect 231486 137912 231492 137964
rect 231544 137952 231550 137964
rect 254026 137952 254032 137964
rect 231544 137924 254032 137952
rect 231544 137912 231550 137924
rect 254026 137912 254032 137924
rect 254084 137912 254090 137964
rect 231762 137844 231768 137896
rect 231820 137884 231826 137896
rect 242894 137884 242900 137896
rect 231820 137856 242900 137884
rect 231820 137844 231826 137856
rect 242894 137844 242900 137856
rect 242952 137844 242958 137896
rect 282822 137436 282828 137488
rect 282880 137476 282886 137488
rect 287054 137476 287060 137488
rect 282880 137448 287060 137476
rect 282880 137436 282886 137448
rect 287054 137436 287060 137448
rect 287112 137436 287118 137488
rect 181530 137232 181536 137284
rect 181588 137272 181594 137284
rect 214006 137272 214012 137284
rect 181588 137244 214012 137272
rect 181588 137232 181594 137244
rect 214006 137232 214012 137244
rect 214064 137232 214070 137284
rect 3510 136892 3516 136944
rect 3568 136932 3574 136944
rect 7558 136932 7564 136944
rect 3568 136904 7564 136932
rect 3568 136892 3574 136904
rect 7558 136892 7564 136904
rect 7616 136892 7622 136944
rect 257522 136688 257528 136740
rect 257580 136728 257586 136740
rect 264974 136728 264980 136740
rect 257580 136700 264980 136728
rect 257580 136688 257586 136700
rect 264974 136688 264980 136700
rect 265032 136688 265038 136740
rect 171778 136620 171784 136672
rect 171836 136660 171842 136672
rect 213914 136660 213920 136672
rect 171836 136632 213920 136660
rect 171836 136620 171842 136632
rect 213914 136620 213920 136632
rect 213972 136620 213978 136672
rect 243722 136620 243728 136672
rect 243780 136660 243786 136672
rect 265066 136660 265072 136672
rect 243780 136632 265072 136660
rect 243780 136620 243786 136632
rect 265066 136620 265072 136632
rect 265124 136620 265130 136672
rect 231762 136552 231768 136604
rect 231820 136592 231826 136604
rect 256694 136592 256700 136604
rect 231820 136564 256700 136592
rect 231820 136552 231826 136564
rect 256694 136552 256700 136564
rect 256752 136552 256758 136604
rect 282822 136552 282828 136604
rect 282880 136592 282886 136604
rect 296898 136592 296904 136604
rect 282880 136564 296904 136592
rect 282880 136552 282886 136564
rect 296898 136552 296904 136564
rect 296956 136552 296962 136604
rect 231670 136484 231676 136536
rect 231728 136524 231734 136536
rect 245010 136524 245016 136536
rect 231728 136496 245016 136524
rect 231728 136484 231734 136496
rect 245010 136484 245016 136496
rect 245068 136484 245074 136536
rect 170398 135872 170404 135924
rect 170456 135912 170462 135924
rect 209130 135912 209136 135924
rect 170456 135884 209136 135912
rect 170456 135872 170462 135884
rect 209130 135872 209136 135884
rect 209188 135872 209194 135924
rect 187050 135260 187056 135312
rect 187108 135300 187114 135312
rect 213914 135300 213920 135312
rect 187108 135272 213920 135300
rect 187108 135260 187114 135272
rect 213914 135260 213920 135272
rect 213972 135260 213978 135312
rect 256234 135260 256240 135312
rect 256292 135300 256298 135312
rect 264974 135300 264980 135312
rect 256292 135272 264980 135300
rect 256292 135260 256298 135272
rect 264974 135260 264980 135272
rect 265032 135260 265038 135312
rect 231762 135192 231768 135244
rect 231820 135232 231826 135244
rect 256142 135232 256148 135244
rect 231820 135204 256148 135232
rect 231820 135192 231826 135204
rect 256142 135192 256148 135204
rect 256200 135192 256206 135244
rect 231670 135124 231676 135176
rect 231728 135164 231734 135176
rect 249150 135164 249156 135176
rect 231728 135136 249156 135164
rect 231728 135124 231734 135136
rect 249150 135124 249156 135136
rect 249208 135124 249214 135176
rect 166258 134580 166264 134632
rect 166316 134620 166322 134632
rect 185578 134620 185584 134632
rect 166316 134592 185584 134620
rect 166316 134580 166322 134592
rect 185578 134580 185584 134592
rect 185636 134580 185642 134632
rect 178862 134512 178868 134564
rect 178920 134552 178926 134564
rect 214006 134552 214012 134564
rect 178920 134524 214012 134552
rect 178920 134512 178926 134524
rect 214006 134512 214012 134524
rect 214064 134512 214070 134564
rect 261754 133968 261760 134020
rect 261812 134008 261818 134020
rect 265066 134008 265072 134020
rect 261812 133980 265072 134008
rect 261812 133968 261818 133980
rect 265066 133968 265072 133980
rect 265124 133968 265130 134020
rect 204990 133900 204996 133952
rect 205048 133940 205054 133952
rect 213914 133940 213920 133952
rect 205048 133912 213920 133940
rect 205048 133900 205054 133912
rect 213914 133900 213920 133912
rect 213972 133900 213978 133952
rect 257430 133900 257436 133952
rect 257488 133940 257494 133952
rect 264974 133940 264980 133952
rect 257488 133912 264980 133940
rect 257488 133900 257494 133912
rect 264974 133900 264980 133912
rect 265032 133900 265038 133952
rect 231486 133832 231492 133884
rect 231544 133872 231550 133884
rect 250530 133872 250536 133884
rect 231544 133844 250536 133872
rect 231544 133832 231550 133844
rect 250530 133832 250536 133844
rect 250588 133832 250594 133884
rect 282822 133832 282828 133884
rect 282880 133872 282886 133884
rect 309318 133872 309324 133884
rect 282880 133844 309324 133872
rect 282880 133832 282886 133844
rect 309318 133832 309324 133844
rect 309376 133832 309382 133884
rect 230750 133152 230756 133204
rect 230808 133192 230814 133204
rect 239490 133192 239496 133204
rect 230808 133164 239496 133192
rect 230808 133152 230814 133164
rect 239490 133152 239496 133164
rect 239548 133152 239554 133204
rect 202414 132540 202420 132592
rect 202472 132580 202478 132592
rect 213914 132580 213920 132592
rect 202472 132552 213920 132580
rect 202472 132540 202478 132552
rect 213914 132540 213920 132552
rect 213972 132540 213978 132592
rect 173158 132472 173164 132524
rect 173216 132512 173222 132524
rect 214006 132512 214012 132524
rect 173216 132484 214012 132512
rect 173216 132472 173222 132484
rect 214006 132472 214012 132484
rect 214064 132472 214070 132524
rect 230934 132404 230940 132456
rect 230992 132444 230998 132456
rect 244918 132444 244924 132456
rect 230992 132416 244924 132444
rect 230992 132404 230998 132416
rect 244918 132404 244924 132416
rect 244976 132404 244982 132456
rect 282822 132404 282828 132456
rect 282880 132444 282886 132456
rect 311894 132444 311900 132456
rect 282880 132416 311900 132444
rect 282880 132404 282886 132416
rect 311894 132404 311900 132416
rect 311952 132404 311958 132456
rect 181438 131724 181444 131776
rect 181496 131764 181502 131776
rect 209222 131764 209228 131776
rect 181496 131736 209228 131764
rect 181496 131724 181502 131736
rect 209222 131724 209228 131736
rect 209280 131724 209286 131776
rect 264238 131588 264244 131640
rect 264296 131628 264302 131640
rect 267182 131628 267188 131640
rect 264296 131600 267188 131628
rect 264296 131588 264302 131600
rect 267182 131588 267188 131600
rect 267240 131588 267246 131640
rect 230474 131316 230480 131368
rect 230532 131356 230538 131368
rect 233970 131356 233976 131368
rect 230532 131328 233976 131356
rect 230532 131316 230538 131328
rect 233970 131316 233976 131328
rect 234028 131316 234034 131368
rect 209314 131180 209320 131232
rect 209372 131220 209378 131232
rect 213914 131220 213920 131232
rect 209372 131192 213920 131220
rect 209372 131180 209378 131192
rect 213914 131180 213920 131192
rect 213972 131180 213978 131232
rect 205082 131112 205088 131164
rect 205140 131152 205146 131164
rect 214006 131152 214012 131164
rect 205140 131124 214012 131152
rect 205140 131112 205146 131124
rect 214006 131112 214012 131124
rect 214064 131112 214070 131164
rect 245194 131112 245200 131164
rect 245252 131152 245258 131164
rect 264974 131152 264980 131164
rect 245252 131124 264980 131152
rect 245252 131112 245258 131124
rect 264974 131112 264980 131124
rect 265032 131112 265038 131164
rect 231762 131044 231768 131096
rect 231820 131084 231826 131096
rect 260282 131084 260288 131096
rect 231820 131056 260288 131084
rect 231820 131044 231826 131056
rect 260282 131044 260288 131056
rect 260340 131044 260346 131096
rect 231486 130976 231492 131028
rect 231544 131016 231550 131028
rect 242250 131016 242256 131028
rect 231544 130988 242256 131016
rect 231544 130976 231550 130988
rect 242250 130976 242256 130988
rect 242308 130976 242314 131028
rect 282270 130976 282276 131028
rect 282328 131016 282334 131028
rect 285674 131016 285680 131028
rect 282328 130988 285680 131016
rect 282328 130976 282334 130988
rect 285674 130976 285680 130988
rect 285732 130976 285738 131028
rect 207658 129820 207664 129872
rect 207716 129860 207722 129872
rect 213914 129860 213920 129872
rect 207716 129832 213920 129860
rect 207716 129820 207722 129832
rect 213914 129820 213920 129832
rect 213972 129820 213978 129872
rect 164878 129752 164884 129804
rect 164936 129792 164942 129804
rect 214006 129792 214012 129804
rect 164936 129764 214012 129792
rect 164936 129752 164942 129764
rect 214006 129752 214012 129764
rect 214064 129752 214070 129804
rect 253382 129752 253388 129804
rect 253440 129792 253446 129804
rect 264974 129792 264980 129804
rect 253440 129764 264980 129792
rect 253440 129752 253446 129764
rect 264974 129752 264980 129764
rect 265032 129752 265038 129804
rect 231762 129684 231768 129736
rect 231820 129724 231826 129736
rect 247770 129724 247776 129736
rect 231820 129696 247776 129724
rect 231820 129684 231826 129696
rect 247770 129684 247776 129696
rect 247828 129684 247834 129736
rect 282086 129684 282092 129736
rect 282144 129724 282150 129736
rect 301038 129724 301044 129736
rect 282144 129696 301044 129724
rect 282144 129684 282150 129696
rect 301038 129684 301044 129696
rect 301096 129684 301102 129736
rect 231486 129548 231492 129600
rect 231544 129588 231550 129600
rect 236730 129588 236736 129600
rect 231544 129560 236736 129588
rect 231544 129548 231550 129560
rect 236730 129548 236736 129560
rect 236788 129548 236794 129600
rect 167822 129004 167828 129056
rect 167880 129044 167886 129056
rect 206370 129044 206376 129056
rect 167880 129016 206376 129044
rect 167880 129004 167886 129016
rect 206370 129004 206376 129016
rect 206428 129004 206434 129056
rect 210418 128392 210424 128444
rect 210476 128432 210482 128444
rect 214006 128432 214012 128444
rect 210476 128404 214012 128432
rect 210476 128392 210482 128404
rect 214006 128392 214012 128404
rect 214064 128392 214070 128444
rect 261570 128392 261576 128444
rect 261628 128432 261634 128444
rect 265158 128432 265164 128444
rect 261628 128404 265164 128432
rect 261628 128392 261634 128404
rect 265158 128392 265164 128404
rect 265216 128392 265222 128444
rect 196802 128324 196808 128376
rect 196860 128364 196866 128376
rect 213914 128364 213920 128376
rect 196860 128336 213920 128364
rect 196860 128324 196866 128336
rect 213914 128324 213920 128336
rect 213972 128324 213978 128376
rect 244918 128324 244924 128376
rect 244976 128364 244982 128376
rect 264974 128364 264980 128376
rect 244976 128336 264980 128364
rect 244976 128324 244982 128336
rect 264974 128324 264980 128336
rect 265032 128324 265038 128376
rect 231762 128256 231768 128308
rect 231820 128296 231826 128308
rect 253290 128296 253296 128308
rect 231820 128268 253296 128296
rect 231820 128256 231826 128268
rect 253290 128256 253296 128268
rect 253348 128256 253354 128308
rect 281994 128256 282000 128308
rect 282052 128296 282058 128308
rect 311986 128296 311992 128308
rect 282052 128268 311992 128296
rect 282052 128256 282058 128268
rect 311986 128256 311992 128268
rect 312044 128256 312050 128308
rect 231670 128188 231676 128240
rect 231728 128228 231734 128240
rect 248046 128228 248052 128240
rect 231728 128200 248052 128228
rect 231728 128188 231734 128200
rect 248046 128188 248052 128200
rect 248104 128188 248110 128240
rect 282822 128188 282828 128240
rect 282880 128228 282886 128240
rect 306650 128228 306656 128240
rect 282880 128200 306656 128228
rect 282880 128188 282886 128200
rect 306650 128188 306656 128200
rect 306708 128188 306714 128240
rect 174630 127576 174636 127628
rect 174688 127616 174694 127628
rect 211798 127616 211804 127628
rect 174688 127588 211804 127616
rect 174688 127576 174694 127588
rect 211798 127576 211804 127588
rect 211856 127576 211862 127628
rect 247862 127576 247868 127628
rect 247920 127616 247926 127628
rect 265066 127616 265072 127628
rect 247920 127588 265072 127616
rect 247920 127576 247926 127588
rect 265066 127576 265072 127588
rect 265124 127576 265130 127628
rect 59170 126964 59176 127016
rect 59228 127004 59234 127016
rect 65518 127004 65524 127016
rect 59228 126976 65524 127004
rect 59228 126964 59234 126976
rect 65518 126964 65524 126976
rect 65576 126964 65582 127016
rect 195330 126964 195336 127016
rect 195388 127004 195394 127016
rect 213914 127004 213920 127016
rect 195388 126976 213920 127004
rect 195388 126964 195394 126976
rect 213914 126964 213920 126976
rect 213972 126964 213978 127016
rect 231762 126896 231768 126948
rect 231820 126936 231826 126948
rect 245286 126936 245292 126948
rect 231820 126908 245292 126936
rect 231820 126896 231826 126908
rect 245286 126896 245292 126908
rect 245344 126896 245350 126948
rect 282270 126896 282276 126948
rect 282328 126936 282334 126948
rect 296714 126936 296720 126948
rect 282328 126908 296720 126936
rect 282328 126896 282334 126908
rect 296714 126896 296720 126908
rect 296772 126896 296778 126948
rect 173250 126216 173256 126268
rect 173308 126256 173314 126268
rect 214558 126256 214564 126268
rect 173308 126228 214564 126256
rect 173308 126216 173314 126228
rect 214558 126216 214564 126228
rect 214616 126216 214622 126268
rect 231118 126216 231124 126268
rect 231176 126256 231182 126268
rect 246574 126256 246580 126268
rect 231176 126228 246580 126256
rect 231176 126216 231182 126228
rect 246574 126216 246580 126228
rect 246632 126216 246638 126268
rect 253290 125672 253296 125724
rect 253348 125712 253354 125724
rect 265066 125712 265072 125724
rect 253348 125684 265072 125712
rect 253348 125672 253354 125684
rect 265066 125672 265072 125684
rect 265124 125672 265130 125724
rect 206370 125604 206376 125656
rect 206428 125644 206434 125656
rect 213914 125644 213920 125656
rect 206428 125616 213920 125644
rect 206428 125604 206434 125616
rect 213914 125604 213920 125616
rect 213972 125604 213978 125656
rect 249150 125604 249156 125656
rect 249208 125644 249214 125656
rect 264974 125644 264980 125656
rect 249208 125616 264980 125644
rect 249208 125604 249214 125616
rect 264974 125604 264980 125616
rect 265032 125604 265038 125656
rect 282822 125536 282828 125588
rect 282880 125576 282886 125588
rect 317414 125576 317420 125588
rect 282880 125548 317420 125576
rect 282880 125536 282886 125548
rect 317414 125536 317420 125548
rect 317472 125536 317478 125588
rect 282730 125468 282736 125520
rect 282788 125508 282794 125520
rect 314654 125508 314660 125520
rect 282788 125480 314660 125508
rect 282788 125468 282794 125480
rect 314654 125468 314660 125480
rect 314712 125468 314718 125520
rect 230842 124924 230848 124976
rect 230900 124964 230906 124976
rect 242434 124964 242440 124976
rect 230900 124936 242440 124964
rect 230900 124924 230906 124936
rect 242434 124924 242440 124936
rect 242492 124924 242498 124976
rect 171870 124856 171876 124908
rect 171928 124896 171934 124908
rect 206278 124896 206284 124908
rect 171928 124868 206284 124896
rect 171928 124856 171934 124868
rect 206278 124856 206284 124868
rect 206336 124856 206342 124908
rect 230934 124856 230940 124908
rect 230992 124896 230998 124908
rect 250622 124896 250628 124908
rect 230992 124868 250628 124896
rect 230992 124856 230998 124868
rect 250622 124856 250628 124868
rect 250680 124856 250686 124908
rect 252002 124244 252008 124296
rect 252060 124284 252066 124296
rect 265066 124284 265072 124296
rect 252060 124256 265072 124284
rect 252060 124244 252066 124256
rect 265066 124244 265072 124256
rect 265124 124244 265130 124296
rect 191098 124176 191104 124228
rect 191156 124216 191162 124228
rect 213914 124216 213920 124228
rect 191156 124188 213920 124216
rect 191156 124176 191162 124188
rect 213914 124176 213920 124188
rect 213972 124176 213978 124228
rect 243538 124176 243544 124228
rect 243596 124216 243602 124228
rect 264974 124216 264980 124228
rect 243596 124188 264980 124216
rect 243596 124176 243602 124188
rect 264974 124176 264980 124188
rect 265032 124176 265038 124228
rect 282270 124108 282276 124160
rect 282328 124148 282334 124160
rect 296806 124148 296812 124160
rect 282328 124120 296812 124148
rect 282328 124108 282334 124120
rect 296806 124108 296812 124120
rect 296864 124108 296870 124160
rect 282822 124040 282828 124092
rect 282880 124080 282886 124092
rect 294046 124080 294052 124092
rect 282880 124052 294052 124080
rect 282880 124040 282886 124052
rect 294046 124040 294052 124052
rect 294104 124040 294110 124092
rect 231762 123836 231768 123888
rect 231820 123876 231826 123888
rect 235534 123876 235540 123888
rect 231820 123848 235540 123876
rect 231820 123836 231826 123848
rect 235534 123836 235540 123848
rect 235592 123836 235598 123888
rect 230658 123428 230664 123480
rect 230716 123468 230722 123480
rect 243906 123468 243912 123480
rect 230716 123440 243912 123468
rect 230716 123428 230722 123440
rect 243906 123428 243912 123440
rect 243964 123428 243970 123480
rect 250714 123428 250720 123480
rect 250772 123468 250778 123480
rect 263134 123468 263140 123480
rect 250772 123440 263140 123468
rect 250772 123428 250778 123440
rect 263134 123428 263140 123440
rect 263192 123428 263198 123480
rect 187142 122884 187148 122936
rect 187200 122924 187206 122936
rect 214006 122924 214012 122936
rect 187200 122896 214012 122924
rect 187200 122884 187206 122896
rect 214006 122884 214012 122896
rect 214064 122884 214070 122936
rect 166258 122816 166264 122868
rect 166316 122856 166322 122868
rect 213914 122856 213920 122868
rect 166316 122828 213920 122856
rect 166316 122816 166322 122828
rect 213914 122816 213920 122828
rect 213972 122816 213978 122868
rect 240870 122816 240876 122868
rect 240928 122856 240934 122868
rect 264974 122856 264980 122868
rect 240928 122828 264980 122856
rect 240928 122816 240934 122828
rect 264974 122816 264980 122828
rect 265032 122816 265038 122868
rect 282822 122748 282828 122800
rect 282880 122788 282886 122800
rect 307938 122788 307944 122800
rect 282880 122760 307944 122788
rect 282880 122748 282886 122760
rect 307938 122748 307944 122760
rect 307996 122748 308002 122800
rect 231578 122680 231584 122732
rect 231636 122720 231642 122732
rect 254578 122720 254584 122732
rect 231636 122692 254584 122720
rect 231636 122680 231642 122692
rect 254578 122680 254584 122692
rect 254636 122680 254642 122732
rect 230750 122476 230756 122528
rect 230808 122516 230814 122528
rect 232590 122516 232596 122528
rect 230808 122488 232596 122516
rect 230808 122476 230814 122488
rect 232590 122476 232596 122488
rect 232648 122476 232654 122528
rect 169110 122068 169116 122120
rect 169168 122108 169174 122120
rect 214558 122108 214564 122120
rect 169168 122080 214564 122108
rect 169168 122068 169174 122080
rect 214558 122068 214564 122080
rect 214616 122068 214622 122120
rect 203610 121456 203616 121508
rect 203668 121496 203674 121508
rect 213914 121496 213920 121508
rect 203668 121468 213920 121496
rect 203668 121456 203674 121468
rect 213914 121456 213920 121468
rect 213972 121456 213978 121508
rect 253474 121456 253480 121508
rect 253532 121496 253538 121508
rect 264974 121496 264980 121508
rect 253532 121468 264980 121496
rect 253532 121456 253538 121468
rect 264974 121456 264980 121468
rect 265032 121456 265038 121508
rect 231762 121388 231768 121440
rect 231820 121428 231826 121440
rect 255958 121428 255964 121440
rect 231820 121400 255964 121428
rect 231820 121388 231826 121400
rect 255958 121388 255964 121400
rect 256016 121388 256022 121440
rect 282822 121388 282828 121440
rect 282880 121428 282886 121440
rect 302418 121428 302424 121440
rect 282880 121400 302424 121428
rect 282880 121388 282886 121400
rect 302418 121388 302424 121400
rect 302476 121388 302482 121440
rect 231670 120912 231676 120964
rect 231728 120952 231734 120964
rect 238018 120952 238024 120964
rect 231728 120924 238024 120952
rect 231728 120912 231734 120924
rect 238018 120912 238024 120924
rect 238076 120912 238082 120964
rect 193950 120164 193956 120216
rect 194008 120204 194014 120216
rect 213914 120204 213920 120216
rect 194008 120176 213920 120204
rect 194008 120164 194014 120176
rect 213914 120164 213920 120176
rect 213972 120164 213978 120216
rect 177574 120096 177580 120148
rect 177632 120136 177638 120148
rect 214006 120136 214012 120148
rect 177632 120108 214012 120136
rect 177632 120096 177638 120108
rect 214006 120096 214012 120108
rect 214064 120096 214070 120148
rect 260282 120096 260288 120148
rect 260340 120136 260346 120148
rect 264974 120136 264980 120148
rect 260340 120108 264980 120136
rect 260340 120096 260346 120108
rect 264974 120096 264980 120108
rect 265032 120096 265038 120148
rect 231762 120028 231768 120080
rect 231820 120068 231826 120080
rect 258718 120068 258724 120080
rect 231820 120040 258724 120068
rect 231820 120028 231826 120040
rect 258718 120028 258724 120040
rect 258776 120028 258782 120080
rect 282822 120028 282828 120080
rect 282880 120068 282886 120080
rect 302234 120068 302240 120080
rect 282880 120040 302240 120068
rect 282880 120028 282886 120040
rect 302234 120028 302240 120040
rect 302292 120028 302298 120080
rect 282730 119960 282736 120012
rect 282788 120000 282794 120012
rect 288526 120000 288532 120012
rect 282788 119972 288532 120000
rect 282788 119960 282794 119972
rect 288526 119960 288532 119972
rect 288584 119960 288590 120012
rect 211798 118736 211804 118788
rect 211856 118776 211862 118788
rect 214006 118776 214012 118788
rect 211856 118748 214012 118776
rect 211856 118736 211862 118748
rect 214006 118736 214012 118748
rect 214064 118736 214070 118788
rect 263134 118736 263140 118788
rect 263192 118776 263198 118788
rect 265434 118776 265440 118788
rect 263192 118748 265440 118776
rect 263192 118736 263198 118748
rect 265434 118736 265440 118748
rect 265492 118736 265498 118788
rect 176102 118668 176108 118720
rect 176160 118708 176166 118720
rect 213914 118708 213920 118720
rect 176160 118680 213920 118708
rect 176160 118668 176166 118680
rect 213914 118668 213920 118680
rect 213972 118668 213978 118720
rect 231210 118668 231216 118720
rect 231268 118708 231274 118720
rect 238110 118708 238116 118720
rect 231268 118680 238116 118708
rect 231268 118668 231274 118680
rect 238110 118668 238116 118680
rect 238168 118668 238174 118720
rect 255958 118668 255964 118720
rect 256016 118708 256022 118720
rect 264974 118708 264980 118720
rect 256016 118680 264980 118708
rect 256016 118668 256022 118680
rect 264974 118668 264980 118680
rect 265032 118668 265038 118720
rect 231394 118600 231400 118652
rect 231452 118640 231458 118652
rect 251910 118640 251916 118652
rect 231452 118612 251916 118640
rect 231452 118600 231458 118612
rect 251910 118600 251916 118612
rect 251968 118600 251974 118652
rect 282822 118600 282828 118652
rect 282880 118640 282886 118652
rect 309226 118640 309232 118652
rect 282880 118612 309232 118640
rect 282880 118600 282886 118612
rect 309226 118600 309232 118612
rect 309284 118600 309290 118652
rect 282270 118532 282276 118584
rect 282328 118572 282334 118584
rect 292666 118572 292672 118584
rect 282328 118544 292672 118572
rect 282328 118532 282334 118544
rect 292666 118532 292672 118544
rect 292724 118532 292730 118584
rect 238386 117920 238392 117972
rect 238444 117960 238450 117972
rect 249150 117960 249156 117972
rect 238444 117932 249156 117960
rect 238444 117920 238450 117932
rect 249150 117920 249156 117932
rect 249208 117920 249214 117972
rect 231486 117648 231492 117700
rect 231544 117688 231550 117700
rect 236638 117688 236644 117700
rect 231544 117660 236644 117688
rect 231544 117648 231550 117660
rect 236638 117648 236644 117660
rect 236696 117648 236702 117700
rect 206462 117376 206468 117428
rect 206520 117416 206526 117428
rect 213914 117416 213920 117428
rect 206520 117388 213920 117416
rect 206520 117376 206526 117388
rect 213914 117376 213920 117388
rect 213972 117376 213978 117428
rect 254578 117376 254584 117428
rect 254636 117416 254642 117428
rect 264974 117416 264980 117428
rect 254636 117388 264980 117416
rect 254636 117376 254642 117388
rect 264974 117376 264980 117388
rect 265032 117376 265038 117428
rect 170398 117308 170404 117360
rect 170456 117348 170462 117360
rect 214006 117348 214012 117360
rect 170456 117320 214012 117348
rect 170456 117308 170462 117320
rect 214006 117308 214012 117320
rect 214064 117308 214070 117360
rect 249058 117308 249064 117360
rect 249116 117348 249122 117360
rect 265066 117348 265072 117360
rect 249116 117320 265072 117348
rect 249116 117308 249122 117320
rect 265066 117308 265072 117320
rect 265124 117308 265130 117360
rect 231762 117240 231768 117292
rect 231820 117280 231826 117292
rect 241146 117280 241152 117292
rect 231820 117252 241152 117280
rect 231820 117240 231826 117252
rect 241146 117240 241152 117252
rect 241204 117240 241210 117292
rect 282822 117240 282828 117292
rect 282880 117280 282886 117292
rect 303706 117280 303712 117292
rect 282880 117252 303712 117280
rect 282880 117240 282886 117252
rect 303706 117240 303712 117252
rect 303764 117240 303770 117292
rect 231670 116832 231676 116884
rect 231728 116872 231734 116884
rect 235258 116872 235264 116884
rect 231728 116844 235264 116872
rect 231728 116832 231734 116844
rect 235258 116832 235264 116844
rect 235316 116832 235322 116884
rect 199470 116016 199476 116068
rect 199528 116056 199534 116068
rect 213914 116056 213920 116068
rect 199528 116028 213920 116056
rect 199528 116016 199534 116028
rect 213914 116016 213920 116028
rect 213972 116016 213978 116068
rect 240778 116016 240784 116068
rect 240836 116056 240842 116068
rect 265066 116056 265072 116068
rect 240836 116028 265072 116056
rect 240836 116016 240842 116028
rect 265066 116016 265072 116028
rect 265124 116016 265130 116068
rect 177298 115948 177304 116000
rect 177356 115988 177362 116000
rect 214006 115988 214012 116000
rect 177356 115960 214012 115988
rect 177356 115948 177362 115960
rect 214006 115948 214012 115960
rect 214064 115948 214070 116000
rect 236638 115948 236644 116000
rect 236696 115988 236702 116000
rect 264974 115988 264980 116000
rect 236696 115960 264980 115988
rect 236696 115948 236702 115960
rect 264974 115948 264980 115960
rect 265032 115948 265038 116000
rect 231486 115880 231492 115932
rect 231544 115920 231550 115932
rect 264330 115920 264336 115932
rect 231544 115892 264336 115920
rect 231544 115880 231550 115892
rect 264330 115880 264336 115892
rect 264388 115880 264394 115932
rect 282362 115880 282368 115932
rect 282420 115920 282426 115932
rect 305086 115920 305092 115932
rect 282420 115892 305092 115920
rect 282420 115880 282426 115892
rect 305086 115880 305092 115892
rect 305144 115880 305150 115932
rect 282822 115812 282828 115864
rect 282880 115852 282886 115864
rect 303890 115852 303896 115864
rect 282880 115824 303896 115852
rect 282880 115812 282886 115824
rect 303890 115812 303896 115824
rect 303948 115812 303954 115864
rect 168282 115200 168288 115252
rect 168340 115240 168346 115252
rect 183002 115240 183008 115252
rect 168340 115212 183008 115240
rect 168340 115200 168346 115212
rect 183002 115200 183008 115212
rect 183060 115200 183066 115252
rect 203518 114588 203524 114640
rect 203576 114628 203582 114640
rect 214006 114628 214012 114640
rect 203576 114600 214012 114628
rect 203576 114588 203582 114600
rect 214006 114588 214012 114600
rect 214064 114588 214070 114640
rect 230566 114588 230572 114640
rect 230624 114628 230630 114640
rect 232682 114628 232688 114640
rect 230624 114600 232688 114628
rect 230624 114588 230630 114600
rect 232682 114588 232688 114600
rect 232740 114588 232746 114640
rect 183094 114520 183100 114572
rect 183152 114560 183158 114572
rect 213914 114560 213920 114572
rect 183152 114532 213920 114560
rect 183152 114520 183158 114532
rect 213914 114520 213920 114532
rect 213972 114520 213978 114572
rect 249150 114520 249156 114572
rect 249208 114560 249214 114572
rect 264974 114560 264980 114572
rect 249208 114532 264980 114560
rect 249208 114520 249214 114532
rect 264974 114520 264980 114532
rect 265032 114520 265038 114572
rect 231762 114452 231768 114504
rect 231820 114492 231826 114504
rect 267090 114492 267096 114504
rect 231820 114464 267096 114492
rect 231820 114452 231826 114464
rect 267090 114452 267096 114464
rect 267148 114452 267154 114504
rect 282086 114452 282092 114504
rect 282144 114492 282150 114504
rect 307754 114492 307760 114504
rect 282144 114464 307760 114492
rect 282144 114452 282150 114464
rect 307754 114452 307760 114464
rect 307812 114452 307818 114504
rect 231486 114384 231492 114436
rect 231544 114424 231550 114436
rect 241054 114424 241060 114436
rect 231544 114396 241060 114424
rect 231544 114384 231550 114396
rect 241054 114384 241060 114396
rect 241112 114384 241118 114436
rect 167730 113772 167736 113824
rect 167788 113812 167794 113824
rect 184382 113812 184388 113824
rect 167788 113784 184388 113812
rect 167788 113772 167794 113784
rect 184382 113772 184388 113784
rect 184440 113772 184446 113824
rect 261662 113568 261668 113620
rect 261720 113608 261726 113620
rect 264974 113608 264980 113620
rect 261720 113580 264980 113608
rect 261720 113568 261726 113580
rect 264974 113568 264980 113580
rect 265032 113568 265038 113620
rect 211982 113296 211988 113348
rect 212040 113336 212046 113348
rect 214282 113336 214288 113348
rect 212040 113308 214288 113336
rect 212040 113296 212046 113308
rect 214282 113296 214288 113308
rect 214340 113296 214346 113348
rect 184474 113160 184480 113212
rect 184532 113200 184538 113212
rect 213914 113200 213920 113212
rect 184532 113172 213920 113200
rect 184532 113160 184538 113172
rect 213914 113160 213920 113172
rect 213972 113160 213978 113212
rect 231762 113092 231768 113144
rect 231820 113132 231826 113144
rect 262950 113132 262956 113144
rect 231820 113104 262956 113132
rect 231820 113092 231826 113104
rect 262950 113092 262956 113104
rect 263008 113092 263014 113144
rect 282822 113092 282828 113144
rect 282880 113132 282886 113144
rect 291194 113132 291200 113144
rect 282880 113104 291200 113132
rect 282880 113092 282886 113104
rect 291194 113092 291200 113104
rect 291252 113092 291258 113144
rect 231394 113024 231400 113076
rect 231452 113064 231458 113076
rect 249242 113064 249248 113076
rect 231452 113036 249248 113064
rect 231452 113024 231458 113036
rect 249242 113024 249248 113036
rect 249300 113024 249306 113076
rect 282454 113024 282460 113076
rect 282512 113064 282518 113076
rect 285766 113064 285772 113076
rect 282512 113036 285772 113064
rect 282512 113024 282518 113036
rect 285766 113024 285772 113036
rect 285824 113024 285830 113076
rect 202506 112412 202512 112464
rect 202564 112452 202570 112464
rect 214742 112452 214748 112464
rect 202564 112424 214748 112452
rect 202564 112412 202570 112424
rect 214742 112412 214748 112424
rect 214800 112412 214806 112464
rect 210510 111800 210516 111852
rect 210568 111840 210574 111852
rect 213914 111840 213920 111852
rect 210568 111812 213920 111840
rect 210568 111800 210574 111812
rect 213914 111800 213920 111812
rect 213972 111800 213978 111852
rect 260374 111800 260380 111852
rect 260432 111840 260438 111852
rect 264974 111840 264980 111852
rect 260432 111812 264980 111840
rect 260432 111800 260438 111812
rect 264974 111800 264980 111812
rect 265032 111800 265038 111852
rect 230750 111732 230756 111784
rect 230808 111772 230814 111784
rect 234062 111772 234068 111784
rect 230808 111744 234068 111772
rect 230808 111732 230814 111744
rect 234062 111732 234068 111744
rect 234120 111732 234126 111784
rect 282822 111732 282828 111784
rect 282880 111772 282886 111784
rect 289814 111772 289820 111784
rect 282880 111744 289820 111772
rect 282880 111732 282886 111744
rect 289814 111732 289820 111744
rect 289872 111732 289878 111784
rect 281718 111596 281724 111648
rect 281776 111636 281782 111648
rect 284294 111636 284300 111648
rect 281776 111608 284300 111636
rect 281776 111596 281782 111608
rect 284294 111596 284300 111608
rect 284352 111596 284358 111648
rect 231578 111052 231584 111104
rect 231636 111092 231642 111104
rect 250806 111092 250812 111104
rect 231636 111064 250812 111092
rect 231636 111052 231642 111064
rect 250806 111052 250812 111064
rect 250864 111052 250870 111104
rect 177482 110508 177488 110560
rect 177540 110548 177546 110560
rect 213914 110548 213920 110560
rect 177540 110520 213920 110548
rect 177540 110508 177546 110520
rect 213914 110508 213920 110520
rect 213972 110508 213978 110560
rect 261478 110508 261484 110560
rect 261536 110548 261542 110560
rect 265066 110548 265072 110560
rect 261536 110520 265072 110548
rect 261536 110508 261542 110520
rect 265066 110508 265072 110520
rect 265124 110508 265130 110560
rect 167638 110440 167644 110492
rect 167696 110480 167702 110492
rect 214006 110480 214012 110492
rect 167696 110452 214012 110480
rect 167696 110440 167702 110452
rect 214006 110440 214012 110452
rect 214064 110440 214070 110492
rect 247770 110440 247776 110492
rect 247828 110480 247834 110492
rect 264974 110480 264980 110492
rect 247828 110452 264980 110480
rect 247828 110440 247834 110452
rect 264974 110440 264980 110452
rect 265032 110440 265038 110492
rect 231762 110372 231768 110424
rect 231820 110412 231826 110424
rect 242158 110412 242164 110424
rect 231820 110384 242164 110412
rect 231820 110372 231826 110384
rect 242158 110372 242164 110384
rect 242216 110372 242222 110424
rect 282270 110372 282276 110424
rect 282328 110412 282334 110424
rect 299566 110412 299572 110424
rect 282328 110384 299572 110412
rect 282328 110372 282334 110384
rect 299566 110372 299572 110384
rect 299624 110372 299630 110424
rect 282822 110304 282828 110356
rect 282880 110344 282886 110356
rect 298094 110344 298100 110356
rect 282880 110316 298100 110344
rect 282880 110304 282886 110316
rect 298094 110304 298100 110316
rect 298152 110304 298158 110356
rect 231394 109692 231400 109744
rect 231452 109732 231458 109744
rect 249334 109732 249340 109744
rect 231452 109704 249340 109732
rect 231452 109692 231458 109704
rect 249334 109692 249340 109704
rect 249392 109692 249398 109744
rect 173342 109080 173348 109132
rect 173400 109120 173406 109132
rect 213914 109120 213920 109132
rect 173400 109092 213920 109120
rect 173400 109080 173406 109092
rect 213914 109080 213920 109092
rect 213972 109080 213978 109132
rect 251818 109080 251824 109132
rect 251876 109120 251882 109132
rect 265066 109120 265072 109132
rect 251876 109092 265072 109120
rect 251876 109080 251882 109092
rect 265066 109080 265072 109092
rect 265124 109080 265130 109132
rect 171962 109012 171968 109064
rect 172020 109052 172026 109064
rect 214006 109052 214012 109064
rect 172020 109024 214012 109052
rect 172020 109012 172026 109024
rect 214006 109012 214012 109024
rect 214064 109012 214070 109064
rect 242250 109012 242256 109064
rect 242308 109052 242314 109064
rect 264974 109052 264980 109064
rect 242308 109024 264980 109052
rect 242308 109012 242314 109024
rect 264974 109012 264980 109024
rect 265032 109012 265038 109064
rect 168006 108944 168012 108996
rect 168064 108984 168070 108996
rect 169202 108984 169208 108996
rect 168064 108956 169208 108984
rect 168064 108944 168070 108956
rect 169202 108944 169208 108956
rect 169260 108944 169266 108996
rect 231578 108944 231584 108996
rect 231636 108984 231642 108996
rect 256050 108984 256056 108996
rect 231636 108956 256056 108984
rect 231636 108944 231642 108956
rect 256050 108944 256056 108956
rect 256108 108944 256114 108996
rect 282362 108944 282368 108996
rect 282420 108984 282426 108996
rect 295518 108984 295524 108996
rect 282420 108956 295524 108984
rect 282420 108944 282426 108956
rect 295518 108944 295524 108956
rect 295576 108944 295582 108996
rect 231762 108536 231768 108588
rect 231820 108576 231826 108588
rect 236914 108576 236920 108588
rect 231820 108548 236920 108576
rect 231820 108536 231826 108548
rect 236914 108536 236920 108548
rect 236972 108536 236978 108588
rect 192662 108264 192668 108316
rect 192720 108304 192726 108316
rect 202414 108304 202420 108316
rect 192720 108276 202420 108304
rect 192720 108264 192726 108276
rect 202414 108264 202420 108276
rect 202472 108264 202478 108316
rect 236730 108264 236736 108316
rect 236788 108304 236794 108316
rect 246390 108304 246396 108316
rect 236788 108276 246396 108304
rect 236788 108264 236794 108276
rect 246390 108264 246396 108276
rect 246448 108264 246454 108316
rect 282822 107924 282828 107976
rect 282880 107964 282886 107976
rect 287146 107964 287152 107976
rect 282880 107936 287152 107964
rect 282880 107924 282886 107936
rect 287146 107924 287152 107936
rect 287204 107924 287210 107976
rect 202322 107720 202328 107772
rect 202380 107760 202386 107772
rect 213914 107760 213920 107772
rect 202380 107732 213920 107760
rect 202380 107720 202386 107732
rect 213914 107720 213920 107732
rect 213972 107720 213978 107772
rect 258718 107720 258724 107772
rect 258776 107760 258782 107772
rect 265066 107760 265072 107772
rect 258776 107732 265072 107760
rect 258776 107720 258782 107732
rect 265066 107720 265072 107732
rect 265124 107720 265130 107772
rect 165062 107652 165068 107704
rect 165120 107692 165126 107704
rect 214006 107692 214012 107704
rect 165120 107664 214012 107692
rect 165120 107652 165126 107664
rect 214006 107652 214012 107664
rect 214064 107652 214070 107704
rect 250530 107652 250536 107704
rect 250588 107692 250594 107704
rect 264974 107692 264980 107704
rect 250588 107664 264980 107692
rect 250588 107652 250594 107664
rect 264974 107652 264980 107664
rect 265032 107652 265038 107704
rect 231302 107584 231308 107636
rect 231360 107624 231366 107636
rect 259086 107624 259092 107636
rect 231360 107596 259092 107624
rect 231360 107584 231366 107596
rect 259086 107584 259092 107596
rect 259144 107584 259150 107636
rect 231762 107516 231768 107568
rect 231820 107556 231826 107568
rect 239674 107556 239680 107568
rect 231820 107528 239680 107556
rect 231820 107516 231826 107528
rect 239674 107516 239680 107528
rect 239732 107516 239738 107568
rect 209222 106360 209228 106412
rect 209280 106400 209286 106412
rect 214006 106400 214012 106412
rect 209280 106372 214012 106400
rect 209280 106360 209286 106372
rect 214006 106360 214012 106372
rect 214064 106360 214070 106412
rect 258902 106360 258908 106412
rect 258960 106400 258966 106412
rect 265066 106400 265072 106412
rect 258960 106372 265072 106400
rect 258960 106360 258966 106372
rect 265066 106360 265072 106372
rect 265124 106360 265130 106412
rect 181622 106292 181628 106344
rect 181680 106332 181686 106344
rect 213914 106332 213920 106344
rect 181680 106304 213920 106332
rect 181680 106292 181686 106304
rect 213914 106292 213920 106304
rect 213972 106292 213978 106344
rect 252094 106292 252100 106344
rect 252152 106332 252158 106344
rect 264974 106332 264980 106344
rect 252152 106304 264980 106332
rect 252152 106292 252158 106304
rect 264974 106292 264980 106304
rect 265032 106292 265038 106344
rect 231394 106224 231400 106276
rect 231452 106264 231458 106276
rect 262858 106264 262864 106276
rect 231452 106236 262864 106264
rect 231452 106224 231458 106236
rect 262858 106224 262864 106236
rect 262916 106224 262922 106276
rect 282822 106224 282828 106276
rect 282880 106264 282886 106276
rect 291286 106264 291292 106276
rect 282880 106236 291292 106264
rect 282880 106224 282886 106236
rect 291286 106224 291292 106236
rect 291344 106224 291350 106276
rect 231762 106156 231768 106208
rect 231820 106196 231826 106208
rect 247954 106196 247960 106208
rect 231820 106168 247960 106196
rect 231820 106156 231826 106168
rect 247954 106156 247960 106168
rect 248012 106156 248018 106208
rect 166534 105544 166540 105596
rect 166592 105584 166598 105596
rect 203610 105584 203616 105596
rect 166592 105556 203616 105584
rect 166592 105544 166598 105556
rect 203610 105544 203616 105556
rect 203668 105544 203674 105596
rect 205174 104932 205180 104984
rect 205232 104972 205238 104984
rect 213914 104972 213920 104984
rect 205232 104944 213920 104972
rect 205232 104932 205238 104944
rect 213914 104932 213920 104944
rect 213972 104932 213978 104984
rect 262950 104932 262956 104984
rect 263008 104972 263014 104984
rect 265066 104972 265072 104984
rect 263008 104944 265072 104972
rect 263008 104932 263014 104944
rect 265066 104932 265072 104944
rect 265124 104932 265130 104984
rect 176010 104864 176016 104916
rect 176068 104904 176074 104916
rect 214006 104904 214012 104916
rect 176068 104876 214012 104904
rect 176068 104864 176074 104876
rect 214006 104864 214012 104876
rect 214064 104864 214070 104916
rect 253566 104864 253572 104916
rect 253624 104904 253630 104916
rect 264974 104904 264980 104916
rect 253624 104876 264980 104904
rect 253624 104864 253630 104876
rect 264974 104864 264980 104876
rect 265032 104864 265038 104916
rect 282822 104796 282828 104848
rect 282880 104836 282886 104848
rect 292574 104836 292580 104848
rect 282880 104808 292580 104836
rect 282880 104796 282886 104808
rect 292574 104796 292580 104808
rect 292632 104796 292638 104848
rect 231762 104728 231768 104780
rect 231820 104768 231826 104780
rect 238294 104768 238300 104780
rect 231820 104740 238300 104768
rect 231820 104728 231826 104740
rect 238294 104728 238300 104740
rect 238352 104728 238358 104780
rect 231118 104320 231124 104372
rect 231176 104360 231182 104372
rect 235350 104360 235356 104372
rect 231176 104332 235356 104360
rect 231176 104320 231182 104332
rect 235350 104320 235356 104332
rect 235408 104320 235414 104372
rect 181530 103572 181536 103624
rect 181588 103612 181594 103624
rect 214006 103612 214012 103624
rect 181588 103584 214012 103612
rect 181588 103572 181594 103584
rect 214006 103572 214012 103584
rect 214064 103572 214070 103624
rect 170490 103504 170496 103556
rect 170548 103544 170554 103556
rect 213914 103544 213920 103556
rect 170548 103516 213920 103544
rect 170548 103504 170554 103516
rect 213914 103504 213920 103516
rect 213972 103504 213978 103556
rect 238110 103504 238116 103556
rect 238168 103544 238174 103556
rect 264974 103544 264980 103556
rect 238168 103516 264980 103544
rect 238168 103504 238174 103516
rect 264974 103504 264980 103516
rect 265032 103504 265038 103556
rect 231762 103436 231768 103488
rect 231820 103476 231826 103488
rect 240962 103476 240968 103488
rect 231820 103448 240968 103476
rect 231820 103436 231826 103448
rect 240962 103436 240968 103448
rect 241020 103436 241026 103488
rect 282822 103436 282828 103488
rect 282880 103476 282886 103488
rect 289998 103476 290004 103488
rect 282880 103448 290004 103476
rect 282880 103436 282886 103448
rect 289998 103436 290004 103448
rect 290056 103436 290062 103488
rect 241054 102824 241060 102876
rect 241112 102864 241118 102876
rect 263134 102864 263140 102876
rect 241112 102836 263140 102864
rect 241112 102824 241118 102836
rect 263134 102824 263140 102836
rect 263192 102824 263198 102876
rect 169202 102756 169208 102808
rect 169260 102796 169266 102808
rect 213178 102796 213184 102808
rect 169260 102768 213184 102796
rect 169260 102756 169266 102768
rect 213178 102756 213184 102768
rect 213236 102756 213242 102808
rect 231026 102756 231032 102808
rect 231084 102796 231090 102808
rect 256326 102796 256332 102808
rect 231084 102768 256332 102796
rect 231084 102756 231090 102768
rect 256326 102756 256332 102768
rect 256384 102756 256390 102808
rect 262766 102212 262772 102264
rect 262824 102252 262830 102264
rect 265158 102252 265164 102264
rect 262824 102224 265164 102252
rect 262824 102212 262830 102224
rect 265158 102212 265164 102224
rect 265216 102212 265222 102264
rect 256142 102144 256148 102196
rect 256200 102184 256206 102196
rect 264974 102184 264980 102196
rect 256200 102156 264980 102184
rect 256200 102144 256206 102156
rect 264974 102144 264980 102156
rect 265032 102144 265038 102196
rect 231670 102076 231676 102128
rect 231728 102116 231734 102128
rect 254762 102116 254768 102128
rect 231728 102088 254768 102116
rect 231728 102076 231734 102088
rect 254762 102076 254768 102088
rect 254820 102076 254826 102128
rect 230566 102008 230572 102060
rect 230624 102048 230630 102060
rect 242342 102048 242348 102060
rect 230624 102020 242348 102048
rect 230624 102008 230630 102020
rect 242342 102008 242348 102020
rect 242400 102008 242406 102060
rect 281718 102008 281724 102060
rect 281776 102048 281782 102060
rect 284386 102048 284392 102060
rect 281776 102020 284392 102048
rect 281776 102008 281782 102020
rect 284386 102008 284392 102020
rect 284444 102008 284450 102060
rect 173434 101396 173440 101448
rect 173492 101436 173498 101448
rect 189810 101436 189816 101448
rect 173492 101408 189816 101436
rect 173492 101396 173498 101408
rect 189810 101396 189816 101408
rect 189868 101396 189874 101448
rect 169294 100716 169300 100768
rect 169352 100756 169358 100768
rect 213914 100756 213920 100768
rect 169352 100728 213920 100756
rect 169352 100716 169358 100728
rect 213914 100716 213920 100728
rect 213972 100716 213978 100768
rect 246390 100716 246396 100768
rect 246448 100756 246454 100768
rect 264974 100756 264980 100768
rect 246448 100728 264980 100756
rect 246448 100716 246454 100728
rect 264974 100716 264980 100728
rect 265032 100716 265038 100768
rect 230566 100648 230572 100700
rect 230624 100688 230630 100700
rect 263042 100688 263048 100700
rect 230624 100660 263048 100688
rect 230624 100648 230630 100660
rect 263042 100648 263048 100660
rect 263100 100648 263106 100700
rect 281718 100648 281724 100700
rect 281776 100688 281782 100700
rect 302326 100688 302332 100700
rect 281776 100660 302332 100688
rect 281776 100648 281782 100660
rect 302326 100648 302332 100660
rect 302384 100648 302390 100700
rect 231118 100580 231124 100632
rect 231176 100620 231182 100632
rect 238202 100620 238208 100632
rect 231176 100592 238208 100620
rect 231176 100580 231182 100592
rect 238202 100580 238208 100592
rect 238260 100580 238266 100632
rect 211890 99424 211896 99476
rect 211948 99464 211954 99476
rect 214006 99464 214012 99476
rect 211948 99436 214012 99464
rect 211948 99424 211954 99436
rect 214006 99424 214012 99436
rect 214064 99424 214070 99476
rect 263134 99424 263140 99476
rect 263192 99464 263198 99476
rect 265066 99464 265072 99476
rect 263192 99436 265072 99464
rect 263192 99424 263198 99436
rect 265066 99424 265072 99436
rect 265124 99424 265130 99476
rect 170674 99356 170680 99408
rect 170732 99396 170738 99408
rect 213914 99396 213920 99408
rect 170732 99368 213920 99396
rect 170732 99356 170738 99368
rect 213914 99356 213920 99368
rect 213972 99356 213978 99408
rect 257614 99356 257620 99408
rect 257672 99396 257678 99408
rect 264974 99396 264980 99408
rect 257672 99368 264980 99396
rect 257672 99356 257678 99368
rect 264974 99356 264980 99368
rect 265032 99356 265038 99408
rect 231118 99288 231124 99340
rect 231176 99328 231182 99340
rect 236822 99328 236828 99340
rect 231176 99300 236828 99328
rect 231176 99288 231182 99300
rect 236822 99288 236828 99300
rect 236880 99288 236886 99340
rect 282822 99288 282828 99340
rect 282880 99328 282886 99340
rect 310514 99328 310520 99340
rect 282880 99300 310520 99328
rect 282880 99288 282886 99300
rect 310514 99288 310520 99300
rect 310572 99288 310578 99340
rect 231670 98608 231676 98660
rect 231728 98648 231734 98660
rect 246298 98648 246304 98660
rect 231728 98620 246304 98648
rect 231728 98608 231734 98620
rect 246298 98608 246304 98620
rect 246356 98608 246362 98660
rect 253382 98064 253388 98116
rect 253440 98104 253446 98116
rect 265066 98104 265072 98116
rect 253440 98076 265072 98104
rect 253440 98064 253446 98076
rect 265066 98064 265072 98076
rect 265124 98064 265130 98116
rect 167822 97996 167828 98048
rect 167880 98036 167886 98048
rect 213914 98036 213920 98048
rect 167880 98008 213920 98036
rect 167880 97996 167886 98008
rect 213914 97996 213920 98008
rect 213972 97996 213978 98048
rect 246574 97996 246580 98048
rect 246632 98036 246638 98048
rect 264974 98036 264980 98048
rect 246632 98008 264980 98036
rect 246632 97996 246638 98008
rect 264974 97996 264980 98008
rect 265032 97996 265038 98048
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 17218 97968 17224 97980
rect 3476 97940 17224 97968
rect 3476 97928 3482 97940
rect 17218 97928 17224 97940
rect 17276 97928 17282 97980
rect 231762 97928 231768 97980
rect 231820 97968 231826 97980
rect 258994 97968 259000 97980
rect 231820 97940 259000 97968
rect 231820 97928 231826 97940
rect 258994 97928 259000 97940
rect 259052 97928 259058 97980
rect 282178 97928 282184 97980
rect 282236 97968 282242 97980
rect 298370 97968 298376 97980
rect 282236 97940 298376 97968
rect 282236 97928 282242 97940
rect 298370 97928 298376 97940
rect 298428 97928 298434 97980
rect 282822 97860 282828 97912
rect 282880 97900 282886 97912
rect 295426 97900 295432 97912
rect 282880 97872 295432 97900
rect 282880 97860 282886 97872
rect 295426 97860 295432 97872
rect 295484 97860 295490 97912
rect 177390 97248 177396 97300
rect 177448 97288 177454 97300
rect 214834 97288 214840 97300
rect 177448 97260 214840 97288
rect 177448 97248 177454 97260
rect 214834 97248 214840 97260
rect 214892 97248 214898 97300
rect 264974 97288 264980 97300
rect 229066 97260 264980 97288
rect 206278 96636 206284 96688
rect 206336 96676 206342 96688
rect 213914 96676 213920 96688
rect 206336 96648 213920 96676
rect 206336 96636 206342 96648
rect 213914 96636 213920 96648
rect 213972 96636 213978 96688
rect 214466 96636 214472 96688
rect 214524 96676 214530 96688
rect 229066 96676 229094 97260
rect 264974 97248 264980 97260
rect 265032 97248 265038 97300
rect 214524 96648 219204 96676
rect 214524 96636 214530 96648
rect 219176 96076 219204 96648
rect 220832 96648 229094 96676
rect 219158 96024 219164 96076
rect 219216 96024 219222 96076
rect 219250 96024 219256 96076
rect 219308 96064 219314 96076
rect 220832 96064 220860 96648
rect 259086 96636 259092 96688
rect 259144 96676 259150 96688
rect 265066 96676 265072 96688
rect 259144 96648 265072 96676
rect 259144 96636 259150 96648
rect 265066 96636 265072 96648
rect 265124 96636 265130 96688
rect 219308 96036 220860 96064
rect 219308 96024 219314 96036
rect 209130 95956 209136 96008
rect 209188 95996 209194 96008
rect 220078 95996 220084 96008
rect 209188 95968 220084 95996
rect 209188 95956 209194 95968
rect 220078 95956 220084 95968
rect 220136 95956 220142 96008
rect 164970 95888 164976 95940
rect 165028 95928 165034 95940
rect 214098 95928 214104 95940
rect 165028 95900 214104 95928
rect 165028 95888 165034 95900
rect 214098 95888 214104 95900
rect 214156 95888 214162 95940
rect 230566 95820 230572 95872
rect 230624 95860 230630 95872
rect 232590 95860 232596 95872
rect 230624 95832 232596 95860
rect 230624 95820 230630 95832
rect 232590 95820 232596 95832
rect 232648 95820 232654 95872
rect 224402 95208 224408 95260
rect 224460 95248 224466 95260
rect 227714 95248 227720 95260
rect 224460 95220 227720 95248
rect 224460 95208 224466 95220
rect 227714 95208 227720 95220
rect 227772 95208 227778 95260
rect 230566 95208 230572 95260
rect 230624 95248 230630 95260
rect 240134 95248 240140 95260
rect 230624 95220 240140 95248
rect 230624 95208 230630 95220
rect 240134 95208 240140 95220
rect 240192 95208 240198 95260
rect 260098 95140 260104 95192
rect 260156 95180 260162 95192
rect 278774 95180 278780 95192
rect 260156 95152 278780 95180
rect 260156 95140 260162 95152
rect 278774 95140 278780 95152
rect 278832 95140 278838 95192
rect 67358 94460 67364 94512
rect 67416 94500 67422 94512
rect 124858 94500 124864 94512
rect 67416 94472 124864 94500
rect 67416 94460 67422 94472
rect 124858 94460 124864 94472
rect 124916 94460 124922 94512
rect 135806 94460 135812 94512
rect 135864 94500 135870 94512
rect 167730 94500 167736 94512
rect 135864 94472 167736 94500
rect 135864 94460 135870 94472
rect 167730 94460 167736 94472
rect 167788 94460 167794 94512
rect 191282 94460 191288 94512
rect 191340 94500 191346 94512
rect 213362 94500 213368 94512
rect 191340 94472 213368 94500
rect 191340 94460 191346 94472
rect 213362 94460 213368 94472
rect 213420 94460 213426 94512
rect 217318 94460 217324 94512
rect 217376 94500 217382 94512
rect 253474 94500 253480 94512
rect 217376 94472 253480 94500
rect 217376 94460 217382 94472
rect 253474 94460 253480 94472
rect 253532 94460 253538 94512
rect 267642 94460 267648 94512
rect 267700 94500 267706 94512
rect 269114 94500 269120 94512
rect 267700 94472 269120 94500
rect 267700 94460 267706 94472
rect 269114 94460 269120 94472
rect 269172 94460 269178 94512
rect 100662 93848 100668 93900
rect 100720 93888 100726 93900
rect 166442 93888 166448 93900
rect 100720 93860 166448 93888
rect 100720 93848 100726 93860
rect 166442 93848 166448 93860
rect 166500 93848 166506 93900
rect 228358 93848 228364 93900
rect 228416 93888 228422 93900
rect 229830 93888 229836 93900
rect 228416 93860 229836 93888
rect 228416 93848 228422 93860
rect 229830 93848 229836 93860
rect 229888 93848 229894 93900
rect 213270 93780 213276 93832
rect 213328 93820 213334 93832
rect 281626 93820 281632 93832
rect 213328 93792 281632 93820
rect 213328 93780 213334 93792
rect 281626 93780 281632 93792
rect 281684 93780 281690 93832
rect 217226 93712 217232 93764
rect 217284 93752 217290 93764
rect 230474 93752 230480 93764
rect 217284 93724 230480 93752
rect 217284 93712 217290 93724
rect 230474 93712 230480 93724
rect 230532 93712 230538 93764
rect 240134 93712 240140 93764
rect 240192 93752 240198 93764
rect 273990 93752 273996 93764
rect 240192 93724 273996 93752
rect 240192 93712 240198 93724
rect 273990 93712 273996 93724
rect 274048 93712 274054 93764
rect 67542 93168 67548 93220
rect 67600 93208 67606 93220
rect 97258 93208 97264 93220
rect 67600 93180 97264 93208
rect 67600 93168 67606 93180
rect 97258 93168 97264 93180
rect 97316 93168 97322 93220
rect 117130 93168 117136 93220
rect 117188 93208 117194 93220
rect 177574 93208 177580 93220
rect 117188 93180 177580 93208
rect 117188 93168 117194 93180
rect 177574 93168 177580 93180
rect 177632 93168 177638 93220
rect 185762 93168 185768 93220
rect 185820 93208 185826 93220
rect 202506 93208 202512 93220
rect 185820 93180 202512 93208
rect 185820 93168 185826 93180
rect 202506 93168 202512 93180
rect 202564 93168 202570 93220
rect 65978 93100 65984 93152
rect 66036 93140 66042 93152
rect 106918 93140 106924 93152
rect 66036 93112 106924 93140
rect 66036 93100 66042 93112
rect 106918 93100 106924 93112
rect 106976 93100 106982 93152
rect 121730 93100 121736 93152
rect 121788 93140 121794 93152
rect 187142 93140 187148 93152
rect 121788 93112 187148 93140
rect 121788 93100 121794 93112
rect 187142 93100 187148 93112
rect 187200 93100 187206 93152
rect 106826 92556 106832 92608
rect 106884 92596 106890 92608
rect 116578 92596 116584 92608
rect 106884 92568 116584 92596
rect 106884 92556 106890 92568
rect 116578 92556 116584 92568
rect 116636 92556 116642 92608
rect 99098 92488 99104 92540
rect 99156 92528 99162 92540
rect 112438 92528 112444 92540
rect 99156 92500 112444 92528
rect 99156 92488 99162 92500
rect 112438 92488 112444 92500
rect 112496 92488 112502 92540
rect 110690 92420 110696 92472
rect 110748 92460 110754 92472
rect 133874 92460 133880 92472
rect 110748 92432 133880 92460
rect 110748 92420 110754 92432
rect 133874 92420 133880 92432
rect 133932 92420 133938 92472
rect 136082 92420 136088 92472
rect 136140 92460 136146 92472
rect 166350 92460 166356 92472
rect 136140 92432 166356 92460
rect 136140 92420 136146 92432
rect 166350 92420 166356 92432
rect 166408 92420 166414 92472
rect 267182 92420 267188 92472
rect 267240 92460 267246 92472
rect 281534 92460 281540 92472
rect 267240 92432 281540 92460
rect 267240 92420 267246 92432
rect 281534 92420 281540 92432
rect 281592 92420 281598 92472
rect 159358 91808 159364 91860
rect 159416 91848 159422 91860
rect 181438 91848 181444 91860
rect 159416 91820 181444 91848
rect 159416 91808 159422 91820
rect 181438 91808 181444 91820
rect 181496 91808 181502 91860
rect 214650 91808 214656 91860
rect 214708 91848 214714 91860
rect 265802 91848 265808 91860
rect 214708 91820 265808 91848
rect 214708 91808 214714 91820
rect 265802 91808 265808 91820
rect 265860 91808 265866 91860
rect 59170 91740 59176 91792
rect 59228 91780 59234 91792
rect 88978 91780 88984 91792
rect 59228 91752 88984 91780
rect 59228 91740 59234 91752
rect 88978 91740 88984 91752
rect 89036 91740 89042 91792
rect 180150 91740 180156 91792
rect 180208 91780 180214 91792
rect 253566 91780 253572 91792
rect 180208 91752 253572 91780
rect 180208 91740 180214 91752
rect 253566 91740 253572 91752
rect 253624 91740 253630 91792
rect 84378 91196 84384 91248
rect 84436 91236 84442 91248
rect 111058 91236 111064 91248
rect 84436 91208 111064 91236
rect 84436 91196 84442 91208
rect 111058 91196 111064 91208
rect 111116 91196 111122 91248
rect 89070 91128 89076 91180
rect 89128 91168 89134 91180
rect 104250 91168 104256 91180
rect 89128 91140 104256 91168
rect 89128 91128 89134 91140
rect 104250 91128 104256 91140
rect 104308 91128 104314 91180
rect 109678 91060 109684 91112
rect 109736 91100 109742 91112
rect 115198 91100 115204 91112
rect 109736 91072 115204 91100
rect 109736 91060 109742 91072
rect 115198 91060 115204 91072
rect 115256 91060 115262 91112
rect 151446 91060 151452 91112
rect 151504 91100 151510 91112
rect 157334 91100 157340 91112
rect 151504 91072 157340 91100
rect 151504 91060 151510 91072
rect 157334 91060 157340 91072
rect 157392 91060 157398 91112
rect 111518 90992 111524 91044
rect 111576 91032 111582 91044
rect 170398 91032 170404 91044
rect 111576 91004 170404 91032
rect 111576 90992 111582 91004
rect 170398 90992 170404 91004
rect 170456 90992 170462 91044
rect 124122 90924 124128 90976
rect 124180 90964 124186 90976
rect 169110 90964 169116 90976
rect 124180 90936 169116 90964
rect 124180 90924 124186 90936
rect 169110 90924 169116 90936
rect 169168 90924 169174 90976
rect 205082 90380 205088 90432
rect 205140 90420 205146 90432
rect 232774 90420 232780 90432
rect 205140 90392 232780 90420
rect 205140 90380 205146 90392
rect 232774 90380 232780 90392
rect 232832 90380 232838 90432
rect 169018 90312 169024 90364
rect 169076 90352 169082 90364
rect 206278 90352 206284 90364
rect 169076 90324 206284 90352
rect 169076 90312 169082 90324
rect 206278 90312 206284 90324
rect 206336 90312 206342 90364
rect 218698 90312 218704 90364
rect 218756 90352 218762 90364
rect 256142 90352 256148 90364
rect 218756 90324 256148 90352
rect 218756 90312 218762 90324
rect 256142 90312 256148 90324
rect 256200 90312 256206 90364
rect 119798 89632 119804 89684
rect 119856 89672 119862 89684
rect 166534 89672 166540 89684
rect 119856 89644 166540 89672
rect 119856 89632 119862 89644
rect 166534 89632 166540 89644
rect 166592 89632 166598 89684
rect 157334 89564 157340 89616
rect 157392 89604 157398 89616
rect 185670 89604 185676 89616
rect 157392 89576 185676 89604
rect 157392 89564 157398 89576
rect 185670 89564 185676 89576
rect 185728 89564 185734 89616
rect 206278 89020 206284 89072
rect 206336 89060 206342 89072
rect 234154 89060 234160 89072
rect 206336 89032 234160 89060
rect 206336 89020 206342 89032
rect 234154 89020 234160 89032
rect 234212 89020 234218 89072
rect 67266 88952 67272 89004
rect 67324 88992 67330 89004
rect 108298 88992 108304 89004
rect 67324 88964 108304 88992
rect 67324 88952 67330 88964
rect 108298 88952 108304 88964
rect 108356 88952 108362 89004
rect 178954 88952 178960 89004
rect 179012 88992 179018 89004
rect 198090 88992 198096 89004
rect 179012 88964 198096 88992
rect 179012 88952 179018 88964
rect 198090 88952 198096 88964
rect 198148 88952 198154 89004
rect 227070 88952 227076 89004
rect 227128 88992 227134 89004
rect 257614 88992 257620 89004
rect 227128 88964 257620 88992
rect 227128 88952 227134 88964
rect 257614 88952 257620 88964
rect 257672 88952 257678 89004
rect 174722 88816 174728 88868
rect 174780 88856 174786 88868
rect 178862 88856 178868 88868
rect 174780 88828 178868 88856
rect 174780 88816 174786 88828
rect 178862 88816 178868 88828
rect 178920 88816 178926 88868
rect 105538 88272 105544 88324
rect 105596 88312 105602 88324
rect 183094 88312 183100 88324
rect 105596 88284 183100 88312
rect 105596 88272 105602 88284
rect 183094 88272 183100 88284
rect 183152 88272 183158 88324
rect 120718 88204 120724 88256
rect 120776 88244 120782 88256
rect 166258 88244 166264 88256
rect 120776 88216 166264 88244
rect 120776 88204 120782 88216
rect 166258 88204 166264 88216
rect 166316 88204 166322 88256
rect 213178 87660 213184 87712
rect 213236 87700 213242 87712
rect 260374 87700 260380 87712
rect 213236 87672 260380 87700
rect 213236 87660 213242 87672
rect 260374 87660 260380 87672
rect 260432 87660 260438 87712
rect 66162 87592 66168 87644
rect 66220 87632 66226 87644
rect 107010 87632 107016 87644
rect 66220 87604 107016 87632
rect 66220 87592 66226 87604
rect 107010 87592 107016 87604
rect 107068 87592 107074 87644
rect 173250 87592 173256 87644
rect 173308 87632 173314 87644
rect 192662 87632 192668 87644
rect 173308 87604 192668 87632
rect 173308 87592 173314 87604
rect 192662 87592 192668 87604
rect 192720 87592 192726 87644
rect 198090 87592 198096 87644
rect 198148 87632 198154 87644
rect 250714 87632 250720 87644
rect 198148 87604 250720 87632
rect 198148 87592 198154 87604
rect 250714 87592 250720 87604
rect 250772 87592 250778 87644
rect 112714 86912 112720 86964
rect 112772 86952 112778 86964
rect 189902 86952 189908 86964
rect 112772 86924 189908 86952
rect 112772 86912 112778 86924
rect 189902 86912 189908 86924
rect 189960 86912 189966 86964
rect 152458 86844 152464 86896
rect 152516 86884 152522 86896
rect 171870 86884 171876 86896
rect 152516 86856 171876 86884
rect 152516 86844 152522 86856
rect 171870 86844 171876 86856
rect 171928 86844 171934 86896
rect 188430 86300 188436 86352
rect 188488 86340 188494 86352
rect 223022 86340 223028 86352
rect 188488 86312 223028 86340
rect 188488 86300 188494 86312
rect 223022 86300 223028 86312
rect 223080 86300 223086 86352
rect 67726 86232 67732 86284
rect 67784 86272 67790 86284
rect 150434 86272 150440 86284
rect 67784 86244 150440 86272
rect 67784 86232 67790 86244
rect 150434 86232 150440 86244
rect 150492 86232 150498 86284
rect 196710 86232 196716 86284
rect 196768 86272 196774 86284
rect 236914 86272 236920 86284
rect 196768 86244 236920 86272
rect 196768 86232 196774 86244
rect 236914 86232 236920 86244
rect 236972 86232 236978 86284
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 14458 85524 14464 85536
rect 3200 85496 14464 85524
rect 3200 85484 3206 85496
rect 14458 85484 14464 85496
rect 14516 85484 14522 85536
rect 104434 85484 104440 85536
rect 104492 85524 104498 85536
rect 184474 85524 184480 85536
rect 104492 85496 184480 85524
rect 104492 85484 104498 85496
rect 184474 85484 184480 85496
rect 184532 85484 184538 85536
rect 115750 85416 115756 85468
rect 115808 85456 115814 85468
rect 193950 85456 193956 85468
rect 115808 85428 193956 85456
rect 115808 85416 115814 85428
rect 193950 85416 193956 85428
rect 194008 85416 194014 85468
rect 225598 84872 225604 84924
rect 225656 84912 225662 84924
rect 232682 84912 232688 84924
rect 225656 84884 232688 84912
rect 225656 84872 225662 84884
rect 232682 84872 232688 84884
rect 232740 84872 232746 84924
rect 49602 84804 49608 84856
rect 49660 84844 49666 84856
rect 83458 84844 83464 84856
rect 49660 84816 83464 84844
rect 49660 84804 49666 84816
rect 83458 84804 83464 84816
rect 83516 84804 83522 84856
rect 195238 84804 195244 84856
rect 195296 84844 195302 84856
rect 281534 84844 281540 84856
rect 195296 84816 281540 84844
rect 195296 84804 195302 84816
rect 281534 84804 281540 84816
rect 281592 84804 281598 84856
rect 97810 84124 97816 84176
rect 97868 84164 97874 84176
rect 171962 84164 171968 84176
rect 97868 84136 171968 84164
rect 97868 84124 97874 84136
rect 171962 84124 171968 84136
rect 172020 84124 172026 84176
rect 126790 84056 126796 84108
rect 126848 84096 126854 84108
rect 185762 84096 185768 84108
rect 126848 84068 185768 84096
rect 126848 84056 126854 84068
rect 185762 84056 185768 84068
rect 185820 84056 185826 84108
rect 222838 83512 222844 83564
rect 222896 83552 222902 83564
rect 249242 83552 249248 83564
rect 222896 83524 249248 83552
rect 222896 83512 222902 83524
rect 249242 83512 249248 83524
rect 249300 83512 249306 83564
rect 86862 83444 86868 83496
rect 86920 83484 86926 83496
rect 126238 83484 126244 83496
rect 86920 83456 126244 83484
rect 86920 83444 86926 83456
rect 126238 83444 126244 83456
rect 126296 83444 126302 83496
rect 211798 83444 211804 83496
rect 211856 83484 211862 83496
rect 239582 83484 239588 83496
rect 211856 83456 239588 83484
rect 211856 83444 211862 83456
rect 239582 83444 239588 83456
rect 239640 83444 239646 83496
rect 88242 82764 88248 82816
rect 88300 82804 88306 82816
rect 170674 82804 170680 82816
rect 88300 82776 170680 82804
rect 88300 82764 88306 82776
rect 170674 82764 170680 82776
rect 170732 82764 170738 82816
rect 111058 82696 111064 82748
rect 111116 82736 111122 82748
rect 169294 82736 169300 82748
rect 111116 82708 169300 82736
rect 111116 82696 111122 82708
rect 169294 82696 169300 82708
rect 169352 82696 169358 82748
rect 195238 82084 195244 82136
rect 195296 82124 195302 82136
rect 247862 82124 247868 82136
rect 195296 82096 247868 82124
rect 195296 82084 195302 82096
rect 247862 82084 247868 82096
rect 247920 82084 247926 82136
rect 67634 81336 67640 81388
rect 67692 81376 67698 81388
rect 181530 81376 181536 81388
rect 67692 81348 181536 81376
rect 67692 81336 67698 81348
rect 181530 81336 181536 81348
rect 181588 81336 181594 81388
rect 95142 81268 95148 81320
rect 95200 81308 95206 81320
rect 202322 81308 202328 81320
rect 95200 81280 202328 81308
rect 95200 81268 95206 81280
rect 202322 81268 202328 81280
rect 202380 81268 202386 81320
rect 204898 80656 204904 80708
rect 204956 80696 204962 80708
rect 235442 80696 235448 80708
rect 204956 80668 235448 80696
rect 204956 80656 204962 80668
rect 235442 80656 235448 80668
rect 235500 80656 235506 80708
rect 97902 79976 97908 80028
rect 97960 80016 97966 80028
rect 195330 80016 195336 80028
rect 97960 79988 195336 80016
rect 97960 79976 97966 79988
rect 195330 79976 195336 79988
rect 195388 79976 195394 80028
rect 126882 79908 126888 79960
rect 126940 79948 126946 79960
rect 159358 79948 159364 79960
rect 126940 79920 159364 79948
rect 126940 79908 126946 79920
rect 159358 79908 159364 79920
rect 159416 79908 159422 79960
rect 224310 79296 224316 79348
rect 224368 79336 224374 79348
rect 238386 79336 238392 79348
rect 224368 79308 238392 79336
rect 224368 79296 224374 79308
rect 238386 79296 238392 79308
rect 238444 79296 238450 79348
rect 122742 78616 122748 78668
rect 122800 78656 122806 78668
rect 174630 78656 174636 78668
rect 122800 78628 174636 78656
rect 122800 78616 122806 78628
rect 174630 78616 174636 78628
rect 174688 78616 174694 78668
rect 151630 78548 151636 78600
rect 151688 78588 151694 78600
rect 169202 78588 169208 78600
rect 151688 78560 169208 78588
rect 151688 78548 151694 78560
rect 169202 78548 169208 78560
rect 169260 78548 169266 78600
rect 175918 77936 175924 77988
rect 175976 77976 175982 77988
rect 273254 77976 273260 77988
rect 175976 77948 273260 77976
rect 175976 77936 175982 77948
rect 273254 77936 273260 77948
rect 273312 77936 273318 77988
rect 128262 77188 128268 77240
rect 128320 77228 128326 77240
rect 173434 77228 173440 77240
rect 128320 77200 173440 77228
rect 128320 77188 128326 77200
rect 173434 77188 173440 77200
rect 173492 77188 173498 77240
rect 106182 76508 106188 76560
rect 106240 76548 106246 76560
rect 240870 76548 240876 76560
rect 106240 76520 240876 76548
rect 106240 76508 106246 76520
rect 240870 76508 240876 76520
rect 240928 76508 240934 76560
rect 107010 75828 107016 75880
rect 107068 75868 107074 75880
rect 178954 75868 178960 75880
rect 107068 75840 178960 75868
rect 107068 75828 107074 75840
rect 178954 75828 178960 75840
rect 179012 75828 179018 75880
rect 111702 75148 111708 75200
rect 111760 75188 111766 75200
rect 229922 75188 229928 75200
rect 111760 75160 229928 75188
rect 111760 75148 111766 75160
rect 229922 75148 229928 75160
rect 229980 75148 229986 75200
rect 91002 74468 91008 74520
rect 91060 74508 91066 74520
rect 176010 74508 176016 74520
rect 91060 74480 176016 74508
rect 91060 74468 91066 74480
rect 176010 74468 176016 74480
rect 176068 74468 176074 74520
rect 117222 73788 117228 73840
rect 117280 73828 117286 73840
rect 252002 73828 252008 73840
rect 117280 73800 252008 73828
rect 117280 73788 117286 73800
rect 252002 73788 252008 73800
rect 252060 73788 252066 73840
rect 151538 73108 151544 73160
rect 151596 73148 151602 73160
rect 192570 73148 192576 73160
rect 151596 73120 192576 73148
rect 151596 73108 151602 73120
rect 192570 73108 192576 73120
rect 192628 73108 192634 73160
rect 126238 73040 126244 73092
rect 126296 73080 126302 73092
rect 164970 73080 164976 73092
rect 126296 73052 164976 73080
rect 126296 73040 126302 73052
rect 164970 73040 164976 73052
rect 165028 73040 165034 73092
rect 583846 72768 583852 72820
rect 583904 72768 583910 72820
rect 583864 72616 583892 72768
rect 583846 72564 583852 72616
rect 583904 72564 583910 72616
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 22738 71720 22744 71732
rect 3476 71692 22744 71720
rect 3476 71680 3482 71692
rect 22738 71680 22744 71692
rect 22796 71680 22802 71732
rect 99190 71680 99196 71732
rect 99248 71720 99254 71732
rect 177482 71720 177488 71732
rect 99248 71692 177488 71720
rect 99248 71680 99254 71692
rect 177482 71680 177488 71692
rect 177540 71680 177546 71732
rect 119982 71000 119988 71052
rect 120040 71040 120046 71052
rect 250622 71040 250628 71052
rect 120040 71012 250628 71040
rect 120040 71000 120046 71012
rect 250622 71000 250628 71012
rect 250680 71000 250686 71052
rect 102042 70320 102048 70372
rect 102100 70360 102106 70372
rect 210510 70360 210516 70372
rect 102100 70332 210516 70360
rect 102100 70320 102106 70332
rect 210510 70320 210516 70332
rect 210568 70320 210574 70372
rect 125410 70252 125416 70304
rect 125468 70292 125474 70304
rect 180242 70292 180248 70304
rect 125468 70264 180248 70292
rect 125468 70252 125474 70264
rect 180242 70252 180248 70264
rect 180300 70252 180306 70304
rect 103422 68960 103428 69012
rect 103480 69000 103486 69012
rect 164878 69000 164884 69012
rect 103480 68972 164884 69000
rect 103480 68960 103486 68972
rect 164878 68960 164884 68972
rect 164936 68960 164942 69012
rect 101398 68280 101404 68332
rect 101456 68320 101462 68332
rect 254670 68320 254676 68332
rect 101456 68292 254676 68320
rect 101456 68280 101462 68292
rect 254670 68280 254676 68292
rect 254728 68280 254734 68332
rect 107562 67532 107568 67584
rect 107620 67572 107626 67584
rect 203518 67572 203524 67584
rect 107620 67544 203524 67572
rect 107620 67532 107626 67544
rect 203518 67532 203524 67544
rect 203576 67532 203582 67584
rect 116578 67464 116584 67516
rect 116636 67504 116642 67516
rect 173250 67504 173256 67516
rect 116636 67476 173256 67504
rect 116636 67464 116642 67476
rect 173250 67464 173256 67476
rect 173308 67464 173314 67516
rect 108298 66172 108304 66224
rect 108356 66212 108362 66224
rect 214742 66212 214748 66224
rect 108356 66184 214748 66212
rect 108356 66172 108362 66184
rect 214742 66172 214748 66184
rect 214800 66172 214806 66224
rect 106090 66104 106096 66156
rect 106148 66144 106154 66156
rect 182910 66144 182916 66156
rect 106148 66116 182916 66144
rect 106148 66104 106154 66116
rect 182910 66104 182916 66116
rect 182968 66104 182974 66156
rect 104250 64812 104256 64864
rect 104308 64852 104314 64864
rect 211890 64852 211896 64864
rect 104308 64824 211896 64852
rect 104308 64812 104314 64824
rect 211890 64812 211896 64824
rect 211948 64812 211954 64864
rect 124030 64744 124036 64796
rect 124088 64784 124094 64796
rect 191098 64784 191104 64796
rect 124088 64756 191104 64784
rect 124088 64744 124094 64756
rect 191098 64744 191104 64756
rect 191156 64744 191162 64796
rect 125502 63452 125508 63504
rect 125560 63492 125566 63504
rect 206370 63492 206376 63504
rect 125560 63464 206376 63492
rect 125560 63452 125566 63464
rect 206370 63452 206376 63464
rect 206428 63452 206434 63504
rect 124858 63384 124864 63436
rect 124916 63424 124922 63436
rect 169018 63424 169024 63436
rect 124916 63396 169024 63424
rect 124916 63384 124922 63396
rect 169018 63384 169024 63396
rect 169076 63384 169082 63436
rect 132402 62024 132408 62076
rect 132460 62064 132466 62076
rect 198182 62064 198188 62076
rect 132460 62036 198188 62064
rect 132460 62024 132466 62036
rect 198182 62024 198188 62036
rect 198240 62024 198246 62076
rect 115842 61956 115848 62008
rect 115900 61996 115906 62008
rect 171778 61996 171784 62008
rect 115900 61968 171784 61996
rect 115900 61956 115906 61968
rect 171778 61956 171784 61968
rect 171836 61956 171842 62008
rect 114370 60664 114376 60716
rect 114428 60704 114434 60716
rect 189718 60704 189724 60716
rect 114428 60676 189724 60704
rect 114428 60664 114434 60676
rect 189718 60664 189724 60676
rect 189776 60664 189782 60716
rect 77202 59984 77208 60036
rect 77260 60024 77266 60036
rect 258902 60024 258908 60036
rect 77260 59996 258908 60024
rect 77260 59984 77266 59996
rect 258902 59984 258908 59996
rect 258960 59984 258966 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 33778 59344 33784 59356
rect 3108 59316 33784 59344
rect 3108 59304 3114 59316
rect 33778 59304 33784 59316
rect 33836 59304 33842 59356
rect 129642 59304 129648 59356
rect 129700 59344 129706 59356
rect 202230 59344 202236 59356
rect 129700 59316 202236 59344
rect 129700 59304 129706 59316
rect 202230 59304 202236 59316
rect 202288 59304 202294 59356
rect 79962 58624 79968 58676
rect 80020 58664 80026 58676
rect 252094 58664 252100 58676
rect 80020 58636 252100 58664
rect 80020 58624 80026 58636
rect 252094 58624 252100 58636
rect 252152 58624 252158 58676
rect 112438 57876 112444 57928
rect 112496 57916 112502 57928
rect 210418 57916 210424 57928
rect 112496 57888 210424 57916
rect 112496 57876 112502 57888
rect 210418 57876 210424 57888
rect 210476 57876 210482 57928
rect 93762 57196 93768 57248
rect 93820 57236 93826 57248
rect 231210 57236 231216 57248
rect 93820 57208 231216 57236
rect 93820 57196 93826 57208
rect 231210 57196 231216 57208
rect 231268 57196 231274 57248
rect 110138 56516 110144 56568
rect 110196 56556 110202 56568
rect 206462 56556 206468 56568
rect 110196 56528 206468 56556
rect 110196 56516 110202 56528
rect 206462 56516 206468 56528
rect 206520 56516 206526 56568
rect 91002 55836 91008 55888
rect 91060 55876 91066 55888
rect 250530 55876 250536 55888
rect 91060 55848 250536 55876
rect 91060 55836 91066 55848
rect 250530 55836 250536 55848
rect 250588 55836 250594 55888
rect 115198 55156 115204 55208
rect 115256 55196 115262 55208
rect 177298 55196 177304 55208
rect 115256 55168 177304 55196
rect 115256 55156 115262 55168
rect 177298 55156 177304 55168
rect 177356 55156 177362 55208
rect 97902 54476 97908 54528
rect 97960 54516 97966 54528
rect 242250 54516 242256 54528
rect 97960 54488 242256 54516
rect 97960 54476 97966 54488
rect 242250 54476 242256 54488
rect 242308 54476 242314 54528
rect 118510 53728 118516 53780
rect 118568 53768 118574 53780
rect 191282 53768 191288 53780
rect 118568 53740 191288 53768
rect 118568 53728 118574 53740
rect 191282 53728 191288 53740
rect 191340 53728 191346 53780
rect 47578 53048 47584 53100
rect 47636 53088 47642 53100
rect 101398 53088 101404 53100
rect 47636 53060 101404 53088
rect 47636 53048 47642 53060
rect 101398 53048 101404 53060
rect 101456 53048 101462 53100
rect 102042 53048 102048 53100
rect 102100 53088 102106 53100
rect 267734 53088 267740 53100
rect 102100 53060 267740 53088
rect 102100 53048 102106 53060
rect 267734 53048 267740 53060
rect 267792 53048 267798 53100
rect 114278 52368 114284 52420
rect 114336 52408 114342 52420
rect 174722 52408 174728 52420
rect 114336 52380 174728 52408
rect 114336 52368 114342 52380
rect 174722 52368 174728 52380
rect 174780 52368 174786 52420
rect 199378 51756 199384 51808
rect 199436 51796 199442 51808
rect 240134 51796 240140 51808
rect 199436 51768 240140 51796
rect 199436 51756 199442 51768
rect 240134 51756 240140 51768
rect 240192 51756 240198 51808
rect 108942 51688 108948 51740
rect 109000 51728 109006 51740
rect 264330 51728 264336 51740
rect 109000 51700 264336 51728
rect 109000 51688 109006 51700
rect 264330 51688 264336 51700
rect 264388 51688 264394 51740
rect 119890 51008 119896 51060
rect 119948 51048 119954 51060
rect 192478 51048 192484 51060
rect 119948 51020 192484 51048
rect 119948 51008 119954 51020
rect 192478 51008 192484 51020
rect 192536 51008 192542 51060
rect 103422 50328 103428 50380
rect 103480 50368 103486 50380
rect 239398 50368 239404 50380
rect 103480 50340 239404 50368
rect 103480 50328 103486 50340
rect 239398 50328 239404 50340
rect 239456 50328 239462 50380
rect 115842 49036 115848 49088
rect 115900 49076 115906 49088
rect 247770 49076 247776 49088
rect 115900 49048 247776 49076
rect 115900 49036 115906 49048
rect 247770 49036 247776 49048
rect 247828 49036 247834 49088
rect 38562 48968 38568 49020
rect 38620 49008 38626 49020
rect 236638 49008 236644 49020
rect 38620 48980 236644 49008
rect 38620 48968 38626 48980
rect 236638 48968 236644 48980
rect 236696 48968 236702 49020
rect 118602 48220 118608 48272
rect 118660 48260 118666 48272
rect 177390 48260 177396 48272
rect 118660 48232 177396 48260
rect 118660 48220 118666 48232
rect 177390 48220 177396 48232
rect 177448 48220 177454 48272
rect 180058 47608 180064 47660
rect 180116 47648 180122 47660
rect 222930 47648 222936 47660
rect 180116 47620 222936 47648
rect 180116 47608 180122 47620
rect 222930 47608 222936 47620
rect 222988 47608 222994 47660
rect 146938 47540 146944 47592
rect 146996 47580 147002 47592
rect 218698 47580 218704 47592
rect 146996 47552 218704 47580
rect 146996 47540 147002 47552
rect 218698 47540 218704 47552
rect 218756 47540 218762 47592
rect 223022 47540 223028 47592
rect 223080 47580 223086 47592
rect 267734 47580 267740 47592
rect 223080 47552 267740 47580
rect 223080 47540 223086 47552
rect 267734 47540 267740 47552
rect 267792 47540 267798 47592
rect 97258 46248 97264 46300
rect 97316 46288 97322 46300
rect 227070 46288 227076 46300
rect 97316 46260 227076 46288
rect 97316 46248 97322 46260
rect 227070 46248 227076 46260
rect 227128 46248 227134 46300
rect 45370 46180 45376 46232
rect 45428 46220 45434 46232
rect 262858 46220 262864 46232
rect 45428 46192 262864 46220
rect 45428 46180 45434 46192
rect 262858 46180 262864 46192
rect 262916 46180 262922 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 21358 45540 21364 45552
rect 3476 45512 21364 45540
rect 3476 45500 3482 45512
rect 21358 45500 21364 45512
rect 21416 45500 21422 45552
rect 125502 44888 125508 44940
rect 125560 44928 125566 44940
rect 236730 44928 236736 44940
rect 125560 44900 236736 44928
rect 125560 44888 125566 44900
rect 236730 44888 236736 44900
rect 236788 44888 236794 44940
rect 86770 44820 86776 44872
rect 86828 44860 86834 44872
rect 251910 44860 251916 44872
rect 86828 44832 251916 44860
rect 86828 44820 86834 44832
rect 251910 44820 251916 44832
rect 251968 44820 251974 44872
rect 174538 43460 174544 43512
rect 174596 43500 174602 43512
rect 241514 43500 241520 43512
rect 174596 43472 241520 43500
rect 174596 43460 174602 43472
rect 241514 43460 241520 43472
rect 241572 43460 241578 43512
rect 88242 43392 88248 43444
rect 88300 43432 88306 43444
rect 205082 43432 205088 43444
rect 88300 43404 205088 43432
rect 88300 43392 88306 43404
rect 205082 43392 205088 43404
rect 205140 43392 205146 43444
rect 231210 43392 231216 43444
rect 231268 43432 231274 43444
rect 269114 43432 269120 43444
rect 231268 43404 269120 43432
rect 231268 43392 231274 43404
rect 269114 43392 269120 43404
rect 269172 43392 269178 43444
rect 56502 42100 56508 42152
rect 56560 42140 56566 42152
rect 249058 42140 249064 42152
rect 56560 42112 249064 42140
rect 56560 42100 56566 42112
rect 249058 42100 249064 42112
rect 249116 42100 249122 42152
rect 19242 42032 19248 42084
rect 19300 42072 19306 42084
rect 235350 42072 235356 42084
rect 19300 42044 235356 42072
rect 19300 42032 19306 42044
rect 235350 42032 235356 42044
rect 235408 42032 235414 42084
rect 62022 40672 62028 40724
rect 62080 40712 62086 40724
rect 324406 40712 324412 40724
rect 62080 40684 324412 40712
rect 62080 40672 62086 40684
rect 324406 40672 324412 40684
rect 324464 40672 324470 40724
rect 112438 39380 112444 39432
rect 112496 39420 112502 39432
rect 230474 39420 230480 39432
rect 112496 39392 230480 39420
rect 112496 39380 112502 39392
rect 230474 39380 230480 39392
rect 230532 39380 230538 39432
rect 53650 39312 53656 39364
rect 53708 39352 53714 39364
rect 254578 39352 254584 39364
rect 53708 39324 254584 39352
rect 53708 39312 53714 39324
rect 254578 39312 254584 39324
rect 254636 39312 254642 39364
rect 62022 37952 62028 38004
rect 62080 37992 62086 38004
rect 260190 37992 260196 38004
rect 62080 37964 260196 37992
rect 62080 37952 62086 37964
rect 260190 37952 260196 37964
rect 260248 37952 260254 38004
rect 30282 37884 30288 37936
rect 30340 37924 30346 37936
rect 242158 37924 242164 37936
rect 30340 37896 242164 37924
rect 30340 37884 30346 37896
rect 242158 37884 242164 37896
rect 242216 37884 242222 37936
rect 60642 36592 60648 36644
rect 60700 36632 60706 36644
rect 248414 36632 248420 36644
rect 60700 36604 248420 36632
rect 60700 36592 60706 36604
rect 248414 36592 248420 36604
rect 248472 36592 248478 36644
rect 49602 36524 49608 36576
rect 49660 36564 49666 36576
rect 266998 36564 267004 36576
rect 49660 36536 267004 36564
rect 49660 36524 49666 36536
rect 266998 36524 267004 36536
rect 267056 36524 267062 36576
rect 111610 35232 111616 35284
rect 111668 35272 111674 35284
rect 261478 35272 261484 35284
rect 111668 35244 261484 35272
rect 111668 35232 111674 35244
rect 261478 35232 261484 35244
rect 261536 35232 261542 35284
rect 43990 35164 43996 35216
rect 44048 35204 44054 35216
rect 253198 35204 253204 35216
rect 44048 35176 253204 35204
rect 44048 35164 44054 35176
rect 253198 35164 253204 35176
rect 253256 35164 253262 35216
rect 71038 33804 71044 33856
rect 71096 33844 71102 33856
rect 215938 33844 215944 33856
rect 71096 33816 215944 33844
rect 71096 33804 71102 33816
rect 215938 33804 215944 33816
rect 215996 33804 216002 33856
rect 59170 33736 59176 33788
rect 59228 33776 59234 33788
rect 267090 33776 267096 33788
rect 59228 33748 267096 33776
rect 59228 33736 59234 33748
rect 267090 33736 267096 33748
rect 267148 33736 267154 33788
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 36538 33096 36544 33108
rect 2924 33068 36544 33096
rect 2924 33056 2930 33068
rect 36538 33056 36544 33068
rect 36596 33056 36602 33108
rect 110322 32444 110328 32496
rect 110380 32484 110386 32496
rect 243538 32484 243544 32496
rect 110380 32456 243544 32484
rect 110380 32444 110386 32456
rect 243538 32444 243544 32456
rect 243596 32444 243602 32496
rect 50982 32376 50988 32428
rect 51040 32416 51046 32428
rect 249794 32416 249800 32428
rect 51040 32388 249800 32416
rect 51040 32376 51046 32388
rect 249794 32376 249800 32388
rect 249852 32376 249858 32428
rect 83458 31084 83464 31136
rect 83516 31124 83522 31136
rect 266998 31124 267004 31136
rect 83516 31096 267004 31124
rect 83516 31084 83522 31096
rect 266998 31084 267004 31096
rect 267056 31084 267062 31136
rect 37090 31016 37096 31068
rect 37148 31056 37154 31068
rect 245102 31056 245108 31068
rect 37148 31028 245108 31056
rect 37148 31016 37154 31028
rect 245102 31016 245108 31028
rect 245160 31016 245166 31068
rect 55030 29588 55036 29640
rect 55088 29628 55094 29640
rect 233970 29628 233976 29640
rect 55088 29600 233976 29628
rect 55088 29588 55094 29600
rect 233970 29588 233976 29600
rect 234028 29588 234034 29640
rect 184290 28296 184296 28348
rect 184348 28336 184354 28348
rect 258074 28336 258080 28348
rect 184348 28308 258080 28336
rect 184348 28296 184354 28308
rect 258074 28296 258080 28308
rect 258132 28296 258138 28348
rect 122742 28228 122748 28280
rect 122800 28268 122806 28280
rect 213178 28268 213184 28280
rect 122800 28240 213184 28268
rect 122800 28228 122806 28240
rect 213178 28228 213184 28240
rect 213236 28228 213242 28280
rect 83458 26936 83464 26988
rect 83516 26976 83522 26988
rect 238110 26976 238116 26988
rect 83516 26948 238116 26976
rect 83516 26936 83522 26948
rect 238110 26936 238116 26948
rect 238168 26936 238174 26988
rect 95050 26868 95056 26920
rect 95108 26908 95114 26920
rect 258718 26908 258724 26920
rect 95108 26880 258724 26908
rect 95108 26868 95114 26880
rect 258718 26868 258724 26880
rect 258776 26868 258782 26920
rect 20622 25576 20628 25628
rect 20680 25616 20686 25628
rect 221458 25616 221464 25628
rect 20680 25588 221464 25616
rect 20680 25576 20686 25588
rect 221458 25576 221464 25588
rect 221516 25576 221522 25628
rect 63402 25508 63408 25560
rect 63460 25548 63466 25560
rect 310514 25548 310520 25560
rect 63460 25520 310520 25548
rect 63460 25508 63466 25520
rect 310514 25508 310520 25520
rect 310572 25508 310578 25560
rect 188522 24148 188528 24200
rect 188580 24188 188586 24200
rect 263594 24188 263600 24200
rect 188580 24160 263600 24188
rect 188580 24148 188586 24160
rect 263594 24148 263600 24160
rect 263652 24148 263658 24200
rect 82722 24080 82728 24132
rect 82780 24120 82786 24132
rect 222838 24120 222844 24132
rect 82780 24092 222844 24120
rect 82780 24080 82786 24092
rect 222838 24080 222844 24092
rect 222896 24080 222902 24132
rect 84102 22720 84108 22772
rect 84160 22760 84166 22772
rect 231118 22760 231124 22772
rect 84160 22732 231124 22760
rect 84160 22720 84166 22732
rect 231118 22720 231124 22732
rect 231176 22720 231182 22772
rect 126238 21428 126244 21480
rect 126296 21468 126302 21480
rect 217318 21468 217324 21480
rect 126296 21440 217324 21468
rect 126296 21428 126302 21440
rect 217318 21428 217324 21440
rect 217376 21428 217382 21480
rect 31662 21360 31668 21412
rect 31720 21400 31726 21412
rect 235258 21400 235264 21412
rect 31720 21372 235264 21400
rect 31720 21360 31726 21372
rect 235258 21360 235264 21372
rect 235316 21360 235322 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 51718 20652 51724 20664
rect 3476 20624 51724 20652
rect 3476 20612 3482 20624
rect 51718 20612 51724 20624
rect 51776 20612 51782 20664
rect 100662 20000 100668 20052
rect 100720 20040 100726 20052
rect 196710 20040 196716 20052
rect 100720 20012 196716 20040
rect 100720 20000 100726 20012
rect 196710 20000 196716 20012
rect 196768 20000 196774 20052
rect 55122 19932 55128 19984
rect 55180 19972 55186 19984
rect 317414 19972 317420 19984
rect 55180 19944 317420 19972
rect 55180 19932 55186 19944
rect 317414 19932 317420 19944
rect 317472 19932 317478 19984
rect 96522 18640 96528 18692
rect 96580 18680 96586 18692
rect 224218 18680 224224 18692
rect 96580 18652 224224 18680
rect 96580 18640 96586 18652
rect 224218 18640 224224 18652
rect 224276 18640 224282 18692
rect 48222 18572 48228 18624
rect 48280 18612 48286 18624
rect 289814 18612 289820 18624
rect 48280 18584 289820 18612
rect 48280 18572 48286 18584
rect 289814 18572 289820 18584
rect 289872 18572 289878 18624
rect 13722 17280 13728 17332
rect 13780 17320 13786 17332
rect 250438 17320 250444 17332
rect 13780 17292 250444 17320
rect 13780 17280 13786 17292
rect 250438 17280 250444 17292
rect 250496 17280 250502 17332
rect 44082 17212 44088 17264
rect 44140 17252 44146 17264
rect 296714 17252 296720 17264
rect 44140 17224 296720 17252
rect 44140 17212 44146 17224
rect 296714 17212 296720 17224
rect 296772 17212 296778 17264
rect 61930 15920 61936 15972
rect 61988 15960 61994 15972
rect 195238 15960 195244 15972
rect 61988 15932 195244 15960
rect 61988 15920 61994 15932
rect 195238 15920 195244 15932
rect 195296 15920 195302 15972
rect 200758 15920 200764 15972
rect 200816 15960 200822 15972
rect 253474 15960 253480 15972
rect 200816 15932 253480 15960
rect 200816 15920 200822 15932
rect 253474 15920 253480 15932
rect 253532 15920 253538 15972
rect 27522 15852 27528 15904
rect 27580 15892 27586 15904
rect 220170 15892 220176 15904
rect 27580 15864 220176 15892
rect 27580 15852 27586 15864
rect 220170 15852 220176 15864
rect 220228 15852 220234 15904
rect 318058 15852 318064 15904
rect 318116 15892 318122 15904
rect 328730 15892 328736 15904
rect 318116 15864 328736 15892
rect 318116 15852 318122 15864
rect 328730 15852 328736 15864
rect 328788 15852 328794 15904
rect 85482 14492 85488 14544
rect 85540 14532 85546 14544
rect 181438 14532 181444 14544
rect 85540 14504 181444 14532
rect 85540 14492 85546 14504
rect 181438 14492 181444 14504
rect 181496 14492 181502 14544
rect 209038 14492 209044 14544
rect 209096 14532 209102 14544
rect 299658 14532 299664 14544
rect 209096 14504 299664 14532
rect 209096 14492 209102 14504
rect 299658 14492 299664 14504
rect 299716 14492 299722 14544
rect 12158 14424 12164 14476
rect 12216 14464 12222 14476
rect 226978 14464 226984 14476
rect 12216 14436 226984 14464
rect 12216 14424 12222 14436
rect 226978 14424 226984 14436
rect 227036 14424 227042 14476
rect 1670 13132 1676 13184
rect 1728 13172 1734 13184
rect 112438 13172 112444 13184
rect 1728 13144 112444 13172
rect 1728 13132 1734 13144
rect 112438 13132 112444 13144
rect 112496 13132 112502 13184
rect 118602 13132 118608 13184
rect 118660 13172 118666 13184
rect 229738 13172 229744 13184
rect 118660 13144 229744 13172
rect 118660 13132 118666 13144
rect 229738 13132 229744 13144
rect 229796 13132 229802 13184
rect 60642 13064 60648 13116
rect 60700 13104 60706 13116
rect 206278 13104 206284 13116
rect 60700 13076 206284 13104
rect 60700 13064 60706 13076
rect 206278 13064 206284 13076
rect 206336 13064 206342 13116
rect 214558 13064 214564 13116
rect 214616 13104 214622 13116
rect 307938 13104 307944 13116
rect 214616 13076 307944 13104
rect 214616 13064 214622 13076
rect 307938 13064 307944 13076
rect 307996 13064 308002 13116
rect 71498 11772 71504 11824
rect 71556 11812 71562 11824
rect 209130 11812 209136 11824
rect 71556 11784 209136 11812
rect 71556 11772 71562 11784
rect 209130 11772 209136 11784
rect 209188 11772 209194 11824
rect 39942 11704 39948 11756
rect 40000 11744 40006 11756
rect 251174 11744 251180 11756
rect 40000 11716 251180 11744
rect 40000 11704 40006 11716
rect 251174 11704 251180 11716
rect 251232 11704 251238 11756
rect 332686 11704 332692 11756
rect 332744 11744 332750 11756
rect 333882 11744 333888 11756
rect 332744 11716 333888 11744
rect 332744 11704 332750 11716
rect 333882 11704 333888 11716
rect 333940 11704 333946 11756
rect 112806 10344 112812 10396
rect 112864 10384 112870 10396
rect 204898 10384 204904 10396
rect 112864 10356 204904 10384
rect 112864 10344 112870 10356
rect 204898 10344 204904 10356
rect 204956 10344 204962 10396
rect 104526 10276 104532 10328
rect 104584 10316 104590 10328
rect 251818 10316 251824 10328
rect 104584 10288 251824 10316
rect 104584 10276 104590 10288
rect 251818 10276 251824 10288
rect 251876 10276 251882 10328
rect 77386 8984 77392 9036
rect 77444 9024 77450 9036
rect 228358 9024 228364 9036
rect 77444 8996 228364 9024
rect 77444 8984 77450 8996
rect 228358 8984 228364 8996
rect 228416 8984 228422 9036
rect 19426 8916 19432 8968
rect 19484 8956 19490 8968
rect 104158 8956 104164 8968
rect 19484 8928 104164 8956
rect 19484 8916 19490 8928
rect 104158 8916 104164 8928
rect 104216 8916 104222 8968
rect 107010 8916 107016 8968
rect 107068 8956 107074 8968
rect 142798 8956 142804 8968
rect 107068 8928 142804 8956
rect 107068 8916 107074 8928
rect 142798 8916 142804 8928
rect 142856 8916 142862 8968
rect 186958 8916 186964 8968
rect 187016 8956 187022 8968
rect 346946 8956 346952 8968
rect 187016 8928 346952 8956
rect 187016 8916 187022 8928
rect 346946 8916 346952 8928
rect 347004 8916 347010 8968
rect 66714 7624 66720 7676
rect 66772 7664 66778 7676
rect 238018 7664 238024 7676
rect 66772 7636 238024 7664
rect 66772 7624 66778 7636
rect 238018 7624 238024 7636
rect 238076 7624 238082 7676
rect 41874 7556 41880 7608
rect 41932 7596 41938 7608
rect 233878 7596 233884 7608
rect 41932 7568 233884 7596
rect 41932 7556 41938 7568
rect 233878 7556 233884 7568
rect 233936 7556 233942 7608
rect 119890 6196 119896 6248
rect 119948 6236 119954 6248
rect 224310 6236 224316 6248
rect 119948 6208 224316 6236
rect 119948 6196 119954 6208
rect 224310 6196 224316 6208
rect 224368 6196 224374 6248
rect 47854 6128 47860 6180
rect 47912 6168 47918 6180
rect 146938 6168 146944 6180
rect 47912 6140 146944 6168
rect 47912 6128 47918 6140
rect 146938 6128 146944 6140
rect 146996 6128 147002 6180
rect 178770 6128 178776 6180
rect 178828 6168 178834 6180
rect 303154 6168 303160 6180
rect 178828 6140 303160 6168
rect 178828 6128 178834 6140
rect 303154 6128 303160 6140
rect 303212 6128 303218 6180
rect 340966 6128 340972 6180
rect 341024 6168 341030 6180
rect 349154 6168 349160 6180
rect 341024 6140 349160 6168
rect 341024 6128 341030 6140
rect 349154 6128 349160 6140
rect 349212 6128 349218 6180
rect 232590 5516 232596 5568
rect 232648 5556 232654 5568
rect 235810 5556 235816 5568
rect 232648 5528 235816 5556
rect 232648 5516 232654 5528
rect 235810 5516 235816 5528
rect 235868 5516 235874 5568
rect 69106 4836 69112 4888
rect 69164 4876 69170 4888
rect 180150 4876 180156 4888
rect 69164 4848 180156 4876
rect 69164 4836 69170 4848
rect 180150 4836 180156 4848
rect 180208 4836 180214 4888
rect 45462 4768 45468 4820
rect 45520 4808 45526 4820
rect 240778 4808 240784 4820
rect 45520 4780 240784 4808
rect 45520 4768 45526 4780
rect 240778 4768 240784 4780
rect 240836 4768 240842 4820
rect 313826 4428 313832 4480
rect 313884 4468 313890 4480
rect 316034 4468 316040 4480
rect 313884 4440 316040 4468
rect 313884 4428 313890 4440
rect 316034 4428 316040 4440
rect 316092 4428 316098 4480
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 12250 3584 12256 3596
rect 11204 3556 12256 3584
rect 11204 3544 11210 3556
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 27706 3544 27712 3596
rect 27764 3584 27770 3596
rect 27764 3556 35894 3584
rect 27764 3544 27770 3556
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3970 3516 3976 3528
rect 2924 3488 3976 3516
rect 2924 3476 2930 3488
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 9582 3516 9588 3528
rect 8812 3488 9588 3516
rect 8812 3476 8818 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 16482 3516 16488 3528
rect 15988 3488 16488 3516
rect 15988 3476 15994 3488
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 17862 3516 17868 3528
rect 17092 3488 17868 3516
rect 17092 3476 17098 3488
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 19242 3516 19248 3528
rect 18288 3488 19248 3516
rect 18288 3476 18294 3488
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 24762 3516 24768 3528
rect 24268 3488 24768 3516
rect 24268 3476 24274 3488
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 25314 3476 25320 3528
rect 25372 3516 25378 3528
rect 26142 3516 26148 3528
rect 25372 3488 26148 3516
rect 25372 3476 25378 3488
rect 26142 3476 26148 3488
rect 26200 3476 26206 3528
rect 26510 3476 26516 3528
rect 26568 3516 26574 3528
rect 27522 3516 27528 3528
rect 26568 3488 27528 3516
rect 26568 3476 26574 3488
rect 27522 3476 27528 3488
rect 27580 3476 27586 3528
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 33042 3516 33048 3528
rect 32456 3488 33048 3516
rect 32456 3476 32462 3488
rect 33042 3476 33048 3488
rect 33100 3476 33106 3528
rect 33594 3476 33600 3528
rect 33652 3516 33658 3528
rect 34422 3516 34428 3528
rect 33652 3488 34428 3516
rect 33652 3476 33658 3488
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
rect 35866 3516 35894 3556
rect 35986 3544 35992 3596
rect 36044 3584 36050 3596
rect 37090 3584 37096 3596
rect 36044 3556 37096 3584
rect 36044 3544 36050 3556
rect 37090 3544 37096 3556
rect 37148 3544 37154 3596
rect 71038 3584 71044 3596
rect 64846 3556 71044 3584
rect 47578 3516 47584 3528
rect 35866 3488 47584 3516
rect 47578 3476 47584 3488
rect 47636 3476 47642 3528
rect 48958 3476 48964 3528
rect 49016 3516 49022 3528
rect 49602 3516 49608 3528
rect 49016 3488 49608 3516
rect 49016 3476 49022 3488
rect 49602 3476 49608 3488
rect 49660 3476 49666 3528
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50890 3516 50896 3528
rect 50212 3488 50896 3516
rect 50212 3476 50218 3488
rect 50890 3476 50896 3488
rect 50948 3476 50954 3528
rect 56042 3476 56048 3528
rect 56100 3516 56106 3528
rect 56502 3516 56508 3528
rect 56100 3488 56508 3516
rect 56100 3476 56106 3488
rect 56502 3476 56508 3488
rect 56560 3476 56566 3528
rect 57238 3476 57244 3528
rect 57296 3516 57302 3528
rect 57882 3516 57888 3528
rect 57296 3488 57888 3516
rect 57296 3476 57302 3488
rect 57882 3476 57888 3488
rect 57940 3476 57946 3528
rect 58434 3476 58440 3528
rect 58492 3516 58498 3528
rect 59170 3516 59176 3528
rect 58492 3488 59176 3516
rect 58492 3476 58498 3488
rect 59170 3476 59176 3488
rect 59228 3476 59234 3528
rect 59630 3476 59636 3528
rect 59688 3516 59694 3528
rect 60642 3516 60648 3528
rect 59688 3488 60648 3516
rect 59688 3476 59694 3488
rect 60642 3476 60648 3488
rect 60700 3476 60706 3528
rect 63218 3476 63224 3528
rect 63276 3516 63282 3528
rect 64846 3516 64874 3556
rect 71038 3544 71044 3556
rect 71096 3544 71102 3596
rect 85666 3544 85672 3596
rect 85724 3584 85730 3596
rect 86770 3584 86776 3596
rect 85724 3556 86776 3584
rect 85724 3544 85730 3556
rect 86770 3544 86776 3556
rect 86828 3544 86834 3596
rect 126238 3584 126244 3596
rect 122806 3556 126244 3584
rect 63276 3488 64874 3516
rect 63276 3476 63282 3488
rect 65518 3476 65524 3528
rect 65576 3516 65582 3528
rect 66162 3516 66168 3528
rect 65576 3488 66168 3516
rect 65576 3476 65582 3488
rect 66162 3476 66168 3488
rect 66220 3476 66226 3528
rect 67910 3476 67916 3528
rect 67968 3516 67974 3528
rect 68922 3516 68928 3528
rect 67968 3488 68928 3516
rect 67968 3476 67974 3488
rect 68922 3476 68928 3488
rect 68980 3476 68986 3528
rect 72602 3476 72608 3528
rect 72660 3516 72666 3528
rect 73062 3516 73068 3528
rect 72660 3488 73068 3516
rect 72660 3476 72666 3488
rect 73062 3476 73068 3488
rect 73120 3476 73126 3528
rect 73798 3476 73804 3528
rect 73856 3516 73862 3528
rect 74442 3516 74448 3528
rect 73856 3488 74448 3516
rect 73856 3476 73862 3488
rect 74442 3476 74448 3488
rect 74500 3476 74506 3528
rect 74994 3476 75000 3528
rect 75052 3516 75058 3528
rect 75822 3516 75828 3528
rect 75052 3488 75828 3516
rect 75052 3476 75058 3488
rect 75822 3476 75828 3488
rect 75880 3476 75886 3528
rect 76190 3476 76196 3528
rect 76248 3516 76254 3528
rect 77202 3516 77208 3528
rect 76248 3488 77208 3516
rect 76248 3476 76254 3488
rect 77202 3476 77208 3488
rect 77260 3476 77266 3528
rect 80882 3476 80888 3528
rect 80940 3516 80946 3528
rect 81342 3516 81348 3528
rect 80940 3488 81348 3516
rect 80940 3476 80946 3488
rect 81342 3476 81348 3488
rect 81400 3476 81406 3528
rect 82078 3476 82084 3528
rect 82136 3516 82142 3528
rect 82722 3516 82728 3528
rect 82136 3488 82728 3516
rect 82136 3476 82142 3488
rect 82722 3476 82728 3488
rect 82780 3476 82786 3528
rect 83274 3476 83280 3528
rect 83332 3516 83338 3528
rect 84102 3516 84108 3528
rect 83332 3488 84108 3516
rect 83332 3476 83338 3488
rect 84102 3476 84108 3488
rect 84160 3476 84166 3528
rect 84470 3476 84476 3528
rect 84528 3516 84534 3528
rect 85482 3516 85488 3528
rect 84528 3488 85488 3516
rect 84528 3476 84534 3488
rect 85482 3476 85488 3488
rect 85540 3476 85546 3528
rect 90358 3476 90364 3528
rect 90416 3516 90422 3528
rect 91002 3516 91008 3528
rect 90416 3488 91008 3516
rect 90416 3476 90422 3488
rect 91002 3476 91008 3488
rect 91060 3476 91066 3528
rect 91554 3476 91560 3528
rect 91612 3516 91618 3528
rect 122806 3516 122834 3556
rect 126238 3544 126244 3556
rect 126296 3544 126302 3596
rect 276014 3544 276020 3596
rect 276072 3584 276078 3596
rect 277118 3584 277124 3596
rect 276072 3556 277124 3584
rect 276072 3544 276078 3556
rect 277118 3544 277124 3556
rect 277176 3544 277182 3596
rect 91612 3488 122834 3516
rect 91612 3476 91618 3488
rect 123478 3476 123484 3528
rect 123536 3516 123542 3528
rect 124122 3516 124128 3528
rect 123536 3488 124128 3516
rect 123536 3476 123542 3488
rect 124122 3476 124128 3488
rect 124180 3476 124186 3528
rect 124674 3476 124680 3528
rect 124732 3516 124738 3528
rect 125502 3516 125508 3528
rect 124732 3488 125508 3516
rect 124732 3476 124738 3488
rect 125502 3476 125508 3488
rect 125560 3476 125566 3528
rect 129366 3476 129372 3528
rect 129424 3516 129430 3528
rect 130378 3516 130384 3528
rect 129424 3488 130384 3516
rect 129424 3476 129430 3488
rect 130378 3476 130384 3488
rect 130436 3476 130442 3528
rect 202138 3476 202144 3528
rect 202196 3516 202202 3528
rect 257062 3516 257068 3528
rect 202196 3488 257068 3516
rect 202196 3476 202202 3488
rect 257062 3476 257068 3488
rect 257120 3476 257126 3528
rect 281442 3476 281448 3528
rect 281500 3516 281506 3528
rect 283098 3516 283104 3528
rect 281500 3488 283104 3516
rect 281500 3476 281506 3488
rect 283098 3476 283104 3488
rect 283156 3476 283162 3528
rect 296070 3476 296076 3528
rect 296128 3516 296134 3528
rect 299474 3516 299480 3528
rect 296128 3488 299480 3516
rect 296128 3476 296134 3488
rect 299474 3476 299480 3488
rect 299532 3476 299538 3528
rect 307754 3476 307760 3528
rect 307812 3516 307818 3528
rect 309042 3516 309048 3528
rect 307812 3488 309048 3516
rect 307812 3476 307818 3488
rect 309042 3476 309048 3488
rect 309100 3476 309106 3528
rect 313918 3476 313924 3528
rect 313976 3516 313982 3528
rect 315022 3516 315028 3528
rect 313976 3488 315028 3516
rect 313976 3476 313982 3488
rect 315022 3476 315028 3488
rect 315080 3476 315086 3528
rect 324314 3476 324320 3528
rect 324372 3516 324378 3528
rect 325602 3516 325608 3528
rect 324372 3488 325608 3516
rect 324372 3476 324378 3488
rect 325602 3476 325608 3488
rect 325660 3476 325666 3528
rect 335998 3476 336004 3528
rect 336056 3516 336062 3528
rect 337470 3516 337476 3528
rect 336056 3488 337476 3516
rect 336056 3476 336062 3488
rect 337470 3476 337476 3488
rect 337528 3476 337534 3528
rect 340874 3476 340880 3528
rect 340932 3516 340938 3528
rect 342162 3516 342168 3528
rect 340932 3488 342168 3516
rect 340932 3476 340938 3488
rect 342162 3476 342168 3488
rect 342220 3476 342226 3528
rect 582190 3476 582196 3528
rect 582248 3516 582254 3528
rect 583386 3516 583392 3528
rect 582248 3488 583392 3516
rect 582248 3476 582254 3488
rect 583386 3476 583392 3488
rect 583444 3476 583450 3528
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 29638 3448 29644 3460
rect 6512 3420 29644 3448
rect 6512 3408 6518 3420
rect 29638 3408 29644 3420
rect 29696 3408 29702 3460
rect 34790 3408 34796 3460
rect 34848 3448 34854 3460
rect 35802 3448 35808 3460
rect 34848 3420 35808 3448
rect 34848 3408 34854 3420
rect 35802 3408 35808 3420
rect 35860 3408 35866 3460
rect 40678 3408 40684 3460
rect 40736 3448 40742 3460
rect 41322 3448 41328 3460
rect 40736 3420 41328 3448
rect 40736 3408 40742 3420
rect 41322 3408 41328 3420
rect 41380 3408 41386 3460
rect 43070 3408 43076 3460
rect 43128 3448 43134 3460
rect 43990 3448 43996 3460
rect 43128 3420 43996 3448
rect 43128 3408 43134 3420
rect 43990 3408 43996 3420
rect 44048 3408 44054 3460
rect 44266 3408 44272 3460
rect 44324 3448 44330 3460
rect 45370 3448 45376 3460
rect 44324 3420 45376 3448
rect 44324 3408 44330 3420
rect 45370 3408 45376 3420
rect 45428 3408 45434 3460
rect 51350 3408 51356 3460
rect 51408 3448 51414 3460
rect 51408 3420 64874 3448
rect 51408 3408 51414 3420
rect 64846 3380 64874 3420
rect 78582 3408 78588 3460
rect 78640 3448 78646 3460
rect 87598 3448 87604 3460
rect 78640 3420 87604 3448
rect 78640 3408 78646 3420
rect 87598 3408 87604 3420
rect 87656 3408 87662 3460
rect 92750 3408 92756 3460
rect 92808 3448 92814 3460
rect 93762 3448 93768 3460
rect 92808 3420 93768 3448
rect 92808 3408 92814 3420
rect 93762 3408 93768 3420
rect 93820 3408 93826 3460
rect 93946 3408 93952 3460
rect 94004 3448 94010 3460
rect 95050 3448 95056 3460
rect 94004 3420 95056 3448
rect 94004 3408 94010 3420
rect 95050 3408 95056 3420
rect 95108 3408 95114 3460
rect 97442 3408 97448 3460
rect 97500 3448 97506 3460
rect 97902 3448 97908 3460
rect 97500 3420 97908 3448
rect 97500 3408 97506 3420
rect 97902 3408 97908 3420
rect 97960 3408 97966 3460
rect 98638 3408 98644 3460
rect 98696 3448 98702 3460
rect 99282 3448 99288 3460
rect 98696 3420 99288 3448
rect 98696 3408 98702 3420
rect 99282 3408 99288 3420
rect 99340 3408 99346 3460
rect 99834 3408 99840 3460
rect 99892 3448 99898 3460
rect 100662 3448 100668 3460
rect 99892 3420 100668 3448
rect 99892 3408 99898 3420
rect 100662 3408 100668 3420
rect 100720 3408 100726 3460
rect 101030 3408 101036 3460
rect 101088 3448 101094 3460
rect 102042 3448 102048 3460
rect 101088 3420 102048 3448
rect 101088 3408 101094 3420
rect 102042 3408 102048 3420
rect 102100 3408 102106 3460
rect 105722 3408 105728 3460
rect 105780 3448 105786 3460
rect 106182 3448 106188 3460
rect 105780 3420 106188 3448
rect 105780 3408 105786 3420
rect 106182 3408 106188 3420
rect 106240 3408 106246 3460
rect 108114 3408 108120 3460
rect 108172 3448 108178 3460
rect 108942 3448 108948 3460
rect 108172 3420 108948 3448
rect 108172 3408 108178 3420
rect 108942 3408 108948 3420
rect 109000 3408 109006 3460
rect 109310 3408 109316 3460
rect 109368 3448 109374 3460
rect 110322 3448 110328 3460
rect 109368 3420 110328 3448
rect 109368 3408 109374 3420
rect 110322 3408 110328 3420
rect 110380 3408 110386 3460
rect 110506 3408 110512 3460
rect 110564 3448 110570 3460
rect 111702 3448 111708 3460
rect 110564 3420 111708 3448
rect 110564 3408 110570 3420
rect 111702 3408 111708 3420
rect 111760 3408 111766 3460
rect 115198 3408 115204 3460
rect 115256 3448 115262 3460
rect 115842 3448 115848 3460
rect 115256 3420 115848 3448
rect 115256 3408 115262 3420
rect 115842 3408 115848 3420
rect 115900 3408 115906 3460
rect 116394 3408 116400 3460
rect 116452 3448 116458 3460
rect 117222 3448 117228 3460
rect 116452 3420 117228 3448
rect 116452 3408 116458 3420
rect 117222 3408 117228 3420
rect 117280 3408 117286 3460
rect 117590 3408 117596 3460
rect 117648 3448 117654 3460
rect 118602 3448 118608 3460
rect 117648 3420 118608 3448
rect 117648 3408 117654 3420
rect 118602 3408 118608 3420
rect 118660 3408 118666 3460
rect 118786 3408 118792 3460
rect 118844 3448 118850 3460
rect 119982 3448 119988 3460
rect 118844 3420 119988 3448
rect 118844 3408 118850 3420
rect 119982 3408 119988 3420
rect 120040 3408 120046 3460
rect 214650 3448 214656 3460
rect 122806 3420 214656 3448
rect 83458 3380 83464 3392
rect 64846 3352 83464 3380
rect 83458 3340 83464 3352
rect 83516 3340 83522 3392
rect 114002 3340 114008 3392
rect 114060 3380 114066 3392
rect 122806 3380 122834 3420
rect 214650 3408 214656 3420
rect 214708 3408 214714 3460
rect 257338 3408 257344 3460
rect 257396 3448 257402 3460
rect 266538 3448 266544 3460
rect 257396 3420 266544 3448
rect 257396 3408 257402 3420
rect 266538 3408 266544 3420
rect 266596 3408 266602 3460
rect 266998 3408 267004 3460
rect 267056 3448 267062 3460
rect 274818 3448 274824 3460
rect 267056 3420 274824 3448
rect 267056 3408 267062 3420
rect 274818 3408 274824 3420
rect 274876 3408 274882 3460
rect 285398 3408 285404 3460
rect 285456 3448 285462 3460
rect 306466 3448 306472 3460
rect 285456 3420 306472 3448
rect 285456 3408 285462 3420
rect 306466 3408 306472 3420
rect 306524 3408 306530 3460
rect 315298 3408 315304 3460
rect 315356 3448 315362 3460
rect 323302 3448 323308 3460
rect 315356 3420 323308 3448
rect 315356 3408 315362 3420
rect 323302 3408 323308 3420
rect 323360 3408 323366 3460
rect 351638 3408 351644 3460
rect 351696 3448 351702 3460
rect 358814 3448 358820 3460
rect 351696 3420 358820 3448
rect 351696 3408 351702 3420
rect 358814 3408 358820 3420
rect 358872 3408 358878 3460
rect 114060 3352 122834 3380
rect 114060 3340 114066 3352
rect 52546 3272 52552 3324
rect 52604 3312 52610 3324
rect 53650 3312 53656 3324
rect 52604 3284 53656 3312
rect 52604 3272 52610 3284
rect 53650 3272 53656 3284
rect 53708 3272 53714 3324
rect 89162 3272 89168 3324
rect 89220 3312 89226 3324
rect 89622 3312 89628 3324
rect 89220 3284 89628 3312
rect 89220 3272 89226 3284
rect 89622 3272 89628 3284
rect 89680 3272 89686 3324
rect 122282 3272 122288 3324
rect 122340 3312 122346 3324
rect 122742 3312 122748 3324
rect 122340 3284 122748 3312
rect 122340 3272 122346 3284
rect 122742 3272 122748 3284
rect 122800 3272 122806 3324
rect 350442 3136 350448 3188
rect 350500 3176 350506 3188
rect 353294 3176 353300 3188
rect 350500 3148 353300 3176
rect 350500 3136 350506 3148
rect 353294 3136 353300 3148
rect 353352 3136 353358 3188
rect 269758 3068 269764 3120
rect 269816 3108 269822 3120
rect 272426 3108 272432 3120
rect 269816 3080 272432 3108
rect 269816 3068 269822 3080
rect 272426 3068 272432 3080
rect 272484 3068 272490 3120
rect 314010 3068 314016 3120
rect 314068 3108 314074 3120
rect 317322 3108 317328 3120
rect 314068 3080 317328 3108
rect 314068 3068 314074 3080
rect 317322 3068 317328 3080
rect 317380 3068 317386 3120
rect 580994 3068 581000 3120
rect 581052 3108 581058 3120
rect 583570 3108 583576 3120
rect 581052 3080 583576 3108
rect 581052 3068 581058 3080
rect 583570 3068 583576 3080
rect 583628 3068 583634 3120
rect 60826 3000 60832 3052
rect 60884 3040 60890 3052
rect 61930 3040 61936 3052
rect 60884 3012 61936 3040
rect 60884 3000 60890 3012
rect 61930 3000 61936 3012
rect 61988 3000 61994 3052
rect 347038 3000 347044 3052
rect 347096 3040 347102 3052
rect 349246 3040 349252 3052
rect 347096 3012 349252 3040
rect 347096 3000 347102 3012
rect 349246 3000 349252 3012
rect 349304 3000 349310 3052
rect 292574 2836 292580 2848
rect 291120 2808 292580 2836
rect 222930 2728 222936 2780
rect 222988 2768 222994 2780
rect 291120 2768 291148 2808
rect 292574 2796 292580 2808
rect 292632 2796 292638 2848
rect 222988 2740 291148 2768
rect 222988 2728 222994 2740
rect 28902 2116 28908 2168
rect 28960 2156 28966 2168
rect 106826 2156 106832 2168
rect 28960 2128 106832 2156
rect 28960 2116 28966 2128
rect 106826 2116 106832 2128
rect 106884 2116 106890 2168
rect 121086 2116 121092 2168
rect 121144 2156 121150 2168
rect 198090 2156 198096 2168
rect 121144 2128 198096 2156
rect 121144 2116 121150 2128
rect 198090 2116 198096 2128
rect 198148 2116 198154 2168
rect 7650 2048 7656 2100
rect 7708 2088 7714 2100
rect 40586 2088 40592 2100
rect 7708 2060 40592 2088
rect 7708 2048 7714 2060
rect 40586 2048 40592 2060
rect 40644 2048 40650 2100
rect 102226 2048 102232 2100
rect 102284 2088 102290 2100
rect 231210 2088 231216 2100
rect 102284 2060 231216 2088
rect 102284 2048 102290 2060
rect 231210 2048 231216 2060
rect 231268 2048 231274 2100
<< via1 >>
rect 75828 703604 75880 703656
rect 202604 703604 202656 703656
rect 86776 703536 86828 703588
rect 234988 703536 235040 703588
rect 67640 703468 67692 703520
rect 267464 703468 267516 703520
rect 93768 703400 93820 703452
rect 300124 703400 300176 703452
rect 59268 703332 59320 703384
rect 283840 703332 283892 703384
rect 73068 703264 73120 703316
rect 332508 703264 332560 703316
rect 130384 703196 130436 703248
rect 413652 703196 413704 703248
rect 61844 703128 61896 703180
rect 348792 703128 348844 703180
rect 101404 703060 101456 703112
rect 397460 703060 397512 703112
rect 124864 702992 124916 703044
rect 429844 702992 429896 703044
rect 57704 702924 57756 702976
rect 364984 702924 365036 702976
rect 126244 702856 126296 702908
rect 462320 702856 462372 702908
rect 71044 702788 71096 702840
rect 494796 702788 494848 702840
rect 97908 702720 97960 702772
rect 478512 702720 478564 702772
rect 129004 702652 129056 702704
rect 543464 702652 543516 702704
rect 8116 702584 8168 702636
rect 89812 702584 89864 702636
rect 94504 702584 94556 702636
rect 527180 702584 527232 702636
rect 53748 702516 53800 702568
rect 580264 702516 580316 702568
rect 66168 702448 66220 702500
rect 559656 702448 559708 702500
rect 84108 700272 84160 700324
rect 89168 700272 89220 700324
rect 88984 700204 89036 700256
rect 105452 700272 105504 700324
rect 133144 700272 133196 700324
rect 218980 700272 219032 700324
rect 24308 698912 24360 698964
rect 79324 698912 79376 698964
rect 3424 683136 3476 683188
rect 18604 683136 18656 683188
rect 3516 656888 3568 656940
rect 22744 656888 22796 656940
rect 3424 639548 3476 639600
rect 39304 639548 39356 639600
rect 3424 632068 3476 632120
rect 11704 632068 11756 632120
rect 3148 618264 3200 618316
rect 15844 618264 15896 618316
rect 3240 600924 3292 600976
rect 88800 600924 88852 600976
rect 67456 599564 67508 599616
rect 88984 599564 89036 599616
rect 79324 598884 79376 598936
rect 80060 598884 80112 598936
rect 40040 598204 40092 598256
rect 91100 598204 91152 598256
rect 80060 597524 80112 597576
rect 106924 597524 106976 597576
rect 67548 596776 67600 596828
rect 169760 596776 169812 596828
rect 72424 595416 72476 595468
rect 84108 595416 84160 595468
rect 92480 595416 92532 595468
rect 74172 594804 74224 594856
rect 95884 594804 95936 594856
rect 83464 593444 83516 593496
rect 110420 593444 110472 593496
rect 90364 593376 90416 593428
rect 582748 593376 582800 593428
rect 22744 592628 22796 592680
rect 69020 592628 69072 592680
rect 75828 592084 75880 592136
rect 96620 592084 96672 592136
rect 84108 592016 84160 592068
rect 112444 592016 112496 592068
rect 78404 590792 78456 590844
rect 89076 590792 89128 590844
rect 71688 590724 71740 590776
rect 86224 590724 86276 590776
rect 90364 590724 90416 590776
rect 70308 590656 70360 590708
rect 74448 590656 74500 590708
rect 75000 590656 75052 590708
rect 75828 590656 75880 590708
rect 88800 590656 88852 590708
rect 132500 590656 132552 590708
rect 3424 589976 3476 590028
rect 71688 589976 71740 590028
rect 74448 589976 74500 590028
rect 89720 589976 89772 590028
rect 67732 589908 67784 589960
rect 580172 589908 580224 589960
rect 81440 589228 81492 589280
rect 88248 589228 88300 589280
rect 69480 588616 69532 588668
rect 88984 588616 89036 588668
rect 85304 588548 85356 588600
rect 86960 588548 87012 588600
rect 113180 588548 113232 588600
rect 79784 588412 79836 588464
rect 63316 587868 63368 587920
rect 66812 587868 66864 587920
rect 105544 587120 105596 587172
rect 59176 586508 59228 586560
rect 66260 586508 66312 586560
rect 91192 586508 91244 586560
rect 141424 586508 141476 586560
rect 89076 585760 89128 585812
rect 103520 585760 103572 585812
rect 50988 585148 51040 585200
rect 67732 585148 67784 585200
rect 92112 584400 92164 584452
rect 93768 584400 93820 584452
rect 115204 584400 115256 584452
rect 91928 583652 91980 583704
rect 93768 583652 93820 583704
rect 94504 583652 94556 583704
rect 48136 582360 48188 582412
rect 66812 582360 66864 582412
rect 64696 581000 64748 581052
rect 66996 581000 67048 581052
rect 91192 581000 91244 581052
rect 102784 581000 102836 581052
rect 91192 578212 91244 578264
rect 121552 578212 121604 578264
rect 104808 577464 104860 577516
rect 582472 577464 582524 577516
rect 91192 576852 91244 576904
rect 104808 576852 104860 576904
rect 11704 576104 11756 576156
rect 51080 576104 51132 576156
rect 51080 575492 51132 575544
rect 52276 575492 52328 575544
rect 66904 575492 66956 575544
rect 88892 575492 88944 575544
rect 105636 575492 105688 575544
rect 55036 574744 55088 574796
rect 67456 574744 67508 574796
rect 91928 574744 91980 574796
rect 93768 574744 93820 574796
rect 101404 574744 101456 574796
rect 41328 572704 41380 572756
rect 66444 572704 66496 572756
rect 91100 572704 91152 572756
rect 120816 572704 120868 572756
rect 91100 571412 91152 571464
rect 97264 571412 97316 571464
rect 49608 571344 49660 571396
rect 66444 571344 66496 571396
rect 91192 571344 91244 571396
rect 126980 571344 127032 571396
rect 91100 569916 91152 569968
rect 125600 569916 125652 569968
rect 93768 569168 93820 569220
rect 123392 569168 123444 569220
rect 64788 568556 64840 568608
rect 66812 568556 66864 568608
rect 91100 567808 91152 567860
rect 91284 567808 91336 567860
rect 128360 567808 128412 567860
rect 57796 567196 57848 567248
rect 66904 567196 66956 567248
rect 53656 566448 53708 566500
rect 67548 566448 67600 566500
rect 91100 565836 91152 565888
rect 101404 565836 101456 565888
rect 60004 564408 60056 564460
rect 66628 564408 66680 564460
rect 91100 564408 91152 564460
rect 120632 564408 120684 564460
rect 50896 564340 50948 564392
rect 53748 564340 53800 564392
rect 66444 564340 66496 564392
rect 91100 563048 91152 563100
rect 133880 563048 133932 563100
rect 45468 561688 45520 561740
rect 66444 561688 66496 561740
rect 43996 560260 44048 560312
rect 66628 560260 66680 560312
rect 56508 558900 56560 558952
rect 66628 558900 66680 558952
rect 48228 557540 48280 557592
rect 67640 557540 67692 557592
rect 91192 557540 91244 557592
rect 124220 557540 124272 557592
rect 91192 556180 91244 556232
rect 122104 556180 122156 556232
rect 58900 554752 58952 554804
rect 66352 554752 66404 554804
rect 91192 554752 91244 554804
rect 108948 554752 109000 554804
rect 582472 554752 582524 554804
rect 59268 554684 59320 554736
rect 65524 554684 65576 554736
rect 66260 554684 66312 554736
rect 2780 553800 2832 553852
rect 4804 553800 4856 553852
rect 107108 553052 107160 553104
rect 109040 553052 109092 553104
rect 91192 552100 91244 552152
rect 107016 552100 107068 552152
rect 91284 552032 91336 552084
rect 130476 552032 130528 552084
rect 100024 551284 100076 551336
rect 117320 551284 117372 551336
rect 63408 549244 63460 549296
rect 66536 549244 66588 549296
rect 91192 549244 91244 549296
rect 111064 549244 111116 549296
rect 91836 548496 91888 548548
rect 121460 548496 121512 548548
rect 62028 547884 62080 547936
rect 66536 547884 66588 547936
rect 61844 547748 61896 547800
rect 66812 547748 66864 547800
rect 53748 547136 53800 547188
rect 61844 547136 61896 547188
rect 91284 546456 91336 546508
rect 104164 546456 104216 546508
rect 57888 545708 57940 545760
rect 66168 545708 66220 545760
rect 108120 545708 108172 545760
rect 126244 545708 126296 545760
rect 52368 545028 52420 545080
rect 57704 545028 57756 545080
rect 66812 545028 66864 545080
rect 91284 544348 91336 544400
rect 96528 544348 96580 544400
rect 129004 544348 129056 544400
rect 18604 542988 18656 543040
rect 39948 542988 40000 543040
rect 39948 542376 40000 542428
rect 66812 542376 66864 542428
rect 91284 542376 91336 542428
rect 94504 542376 94556 542428
rect 39304 541628 39356 541680
rect 67088 541628 67140 541680
rect 91284 541628 91336 541680
rect 136640 541628 136692 541680
rect 67548 540880 67600 540932
rect 68652 540880 68704 540932
rect 582656 540880 582708 540932
rect 3424 540200 3476 540252
rect 91284 539656 91336 539708
rect 93124 539656 93176 539708
rect 55128 539588 55180 539640
rect 67548 539588 67600 539640
rect 69848 539588 69900 539640
rect 115388 539520 115440 539572
rect 582564 539520 582616 539572
rect 67088 539452 67140 539504
rect 67548 539452 67600 539504
rect 67824 538976 67876 539028
rect 74632 538976 74684 539028
rect 3424 538840 3476 538892
rect 89904 538840 89956 538892
rect 81072 538228 81124 538280
rect 115388 538228 115440 538280
rect 4804 538160 4856 538212
rect 70676 538160 70728 538212
rect 86868 538160 86920 538212
rect 133144 538160 133196 538212
rect 72424 537480 72476 537532
rect 579804 537480 579856 537532
rect 82728 536732 82780 536784
rect 130384 536732 130436 536784
rect 85488 536188 85540 536240
rect 86224 536188 86276 536240
rect 66168 536120 66220 536172
rect 76196 536120 76248 536172
rect 15844 536052 15896 536104
rect 44088 536052 44140 536104
rect 73160 536052 73212 536104
rect 73160 535440 73212 535492
rect 73988 535440 74040 535492
rect 78772 535440 78824 535492
rect 79508 535440 79560 535492
rect 7564 534692 7616 534744
rect 91376 534692 91428 534744
rect 56508 534012 56560 534064
rect 580264 534012 580316 534064
rect 5448 533332 5500 533384
rect 91192 533332 91244 533384
rect 66076 531972 66128 532024
rect 77944 531972 77996 532024
rect 15844 530544 15896 530596
rect 91100 530544 91152 530596
rect 3516 514768 3568 514820
rect 14464 514768 14516 514820
rect 43996 511232 44048 511284
rect 580172 511232 580224 511284
rect 3332 502052 3384 502104
rect 7564 502052 7616 502104
rect 4068 475328 4120 475380
rect 5448 475328 5500 475380
rect 11704 475328 11756 475380
rect 67732 467780 67784 467832
rect 76564 467780 76616 467832
rect 63316 465060 63368 465112
rect 87052 465060 87104 465112
rect 56416 464312 56468 464364
rect 78772 464312 78824 464364
rect 2780 462544 2832 462596
rect 4804 462544 4856 462596
rect 59176 461592 59228 461644
rect 85580 461592 85632 461644
rect 64696 460164 64748 460216
rect 78680 460164 78732 460216
rect 64696 458872 64748 458924
rect 70492 458872 70544 458924
rect 53472 458804 53524 458856
rect 77300 458804 77352 458856
rect 102784 458804 102836 458856
rect 123116 458804 123168 458856
rect 50988 457444 51040 457496
rect 83464 457444 83516 457496
rect 105636 457444 105688 457496
rect 122932 457444 122984 457496
rect 60556 456084 60608 456136
rect 76104 456084 76156 456136
rect 101404 456084 101456 456136
rect 123576 456084 123628 456136
rect 61936 456016 61988 456068
rect 91100 456016 91152 456068
rect 97264 456016 97316 456068
rect 124404 456016 124456 456068
rect 59084 454724 59136 454776
rect 73160 454724 73212 454776
rect 55036 454656 55088 454708
rect 72056 454656 72108 454708
rect 91100 454044 91152 454096
rect 161480 454044 161532 454096
rect 49608 453296 49660 453348
rect 67640 453296 67692 453348
rect 72056 452684 72108 452736
rect 126336 452684 126388 452736
rect 112444 452616 112496 452668
rect 179420 452616 179472 452668
rect 61936 451936 61988 451988
rect 78864 451936 78916 451988
rect 3424 451868 3476 451920
rect 120724 451868 120776 451920
rect 14464 451188 14516 451240
rect 112444 451188 112496 451240
rect 116584 449964 116636 450016
rect 160100 449964 160152 450016
rect 49516 449896 49568 449948
rect 74632 449896 74684 449948
rect 95884 449896 95936 449948
rect 178040 449896 178092 449948
rect 41328 449828 41380 449880
rect 69664 449828 69716 449880
rect 48136 449148 48188 449200
rect 80060 449148 80112 449200
rect 173808 449148 173860 449200
rect 582472 449148 582524 449200
rect 77944 448604 77996 448656
rect 124312 448604 124364 448656
rect 3148 448536 3200 448588
rect 14464 448536 14516 448588
rect 80060 448536 80112 448588
rect 80888 448536 80940 448588
rect 173808 448536 173860 448588
rect 52276 447856 52328 447908
rect 73344 447856 73396 447908
rect 4804 447788 4856 447840
rect 68284 447788 68336 447840
rect 115204 447788 115256 447840
rect 125692 447788 125744 447840
rect 68284 447176 68336 447228
rect 68560 447176 68612 447228
rect 103520 447176 103572 447228
rect 98644 447108 98696 447160
rect 170404 447108 170456 447160
rect 78680 446904 78732 446956
rect 79140 446904 79192 446956
rect 64512 446360 64564 446412
rect 74540 446360 74592 446412
rect 106924 445816 106976 445868
rect 124864 445816 124916 445868
rect 50988 445748 51040 445800
rect 79140 445748 79192 445800
rect 98000 445748 98052 445800
rect 102140 445748 102192 445800
rect 105544 445748 105596 445800
rect 201500 445748 201552 445800
rect 66076 445000 66128 445052
rect 72424 445000 72476 445052
rect 67640 444592 67692 444644
rect 67824 444592 67876 444644
rect 68790 444592 68842 444644
rect 73344 444456 73396 444508
rect 144184 444456 144236 444508
rect 4804 444388 4856 444440
rect 119160 444388 119212 444440
rect 120908 444388 120960 444440
rect 124128 444320 124180 444372
rect 132500 444320 132552 444372
rect 133788 444320 133840 444372
rect 133788 443640 133840 443692
rect 166264 443640 166316 443692
rect 67272 442892 67324 442944
rect 67732 442892 67784 442944
rect 124128 441600 124180 441652
rect 133144 441600 133196 441652
rect 64788 439084 64840 439136
rect 66996 439084 67048 439136
rect 67272 439084 67324 439136
rect 121184 438880 121236 438932
rect 169760 438880 169812 438932
rect 123852 438132 123904 438184
rect 125692 438132 125744 438184
rect 157984 438132 158036 438184
rect 57796 437452 57848 437504
rect 60648 437452 60700 437504
rect 66812 437452 66864 437504
rect 53656 436024 53708 436076
rect 57704 436024 57756 436076
rect 57704 434732 57756 434784
rect 66812 434732 66864 434784
rect 58992 433848 59044 433900
rect 60004 433848 60056 433900
rect 124128 432556 124180 432608
rect 135168 432556 135220 432608
rect 582380 432556 582432 432608
rect 58992 432012 59044 432064
rect 66904 432012 66956 432064
rect 50896 431876 50948 431928
rect 66904 431876 66956 431928
rect 48136 430584 48188 430636
rect 50896 430584 50948 430636
rect 40684 429088 40736 429140
rect 45468 429088 45520 429140
rect 66812 429088 66864 429140
rect 61844 426368 61896 426420
rect 66260 426368 66312 426420
rect 56508 425008 56560 425060
rect 66260 425008 66312 425060
rect 3148 422900 3200 422952
rect 15844 422900 15896 422952
rect 48228 421540 48280 421592
rect 61844 421540 61896 421592
rect 66260 421540 66312 421592
rect 123392 421540 123444 421592
rect 148324 421540 148376 421592
rect 121552 418072 121604 418124
rect 126980 418072 127032 418124
rect 58900 416780 58952 416832
rect 63316 416780 63368 416832
rect 66904 416780 66956 416832
rect 65524 415148 65576 415200
rect 66444 415148 66496 415200
rect 123116 415080 123168 415132
rect 124404 415080 124456 415132
rect 126980 415080 127032 415132
rect 57796 414672 57848 414724
rect 65524 414672 65576 414724
rect 123116 413924 123168 413976
rect 125600 413924 125652 413976
rect 121644 409844 121696 409896
rect 162860 409844 162912 409896
rect 63408 408416 63460 408468
rect 65984 408416 66036 408468
rect 66536 408416 66588 408468
rect 124128 408348 124180 408400
rect 128360 408348 128412 408400
rect 128360 407736 128412 407788
rect 135904 407736 135956 407788
rect 122104 407056 122156 407108
rect 123024 407056 123076 407108
rect 123576 405832 123628 405884
rect 124864 405832 124916 405884
rect 62028 405764 62080 405816
rect 64604 405764 64656 405816
rect 66628 405764 66680 405816
rect 57612 404812 57664 404864
rect 57888 404812 57940 404864
rect 57980 403588 58032 403640
rect 66352 403588 66404 403640
rect 162768 403588 162820 403640
rect 582380 403588 582432 403640
rect 120632 402976 120684 403028
rect 161572 402976 161624 403028
rect 162768 402976 162820 403028
rect 53564 402228 53616 402280
rect 57980 402228 58032 402280
rect 50896 401548 50948 401600
rect 57612 401548 57664 401600
rect 66812 401548 66864 401600
rect 124128 401548 124180 401600
rect 133880 401548 133932 401600
rect 135076 401548 135128 401600
rect 135076 400868 135128 400920
rect 158076 400868 158128 400920
rect 52368 398828 52420 398880
rect 53656 398828 53708 398880
rect 66904 398828 66956 398880
rect 123668 398828 123720 398880
rect 124956 398828 125008 398880
rect 2780 398692 2832 398744
rect 4804 398692 4856 398744
rect 39948 396720 40000 396772
rect 66260 396720 66312 396772
rect 121460 396040 121512 396092
rect 177396 396040 177448 396092
rect 55128 392572 55180 392624
rect 65524 392572 65576 392624
rect 124956 391960 125008 392012
rect 166356 391960 166408 392012
rect 15844 391348 15896 391400
rect 124956 391348 125008 391400
rect 111708 389784 111760 389836
rect 121552 389784 121604 389836
rect 59084 389240 59136 389292
rect 77392 389240 77444 389292
rect 11704 389172 11756 389224
rect 111616 389172 111668 389224
rect 64696 389104 64748 389156
rect 73160 389104 73212 389156
rect 73344 389104 73396 389156
rect 91928 389104 91980 389156
rect 93216 389104 93268 389156
rect 102600 389104 102652 389156
rect 105544 389104 105596 389156
rect 117872 389104 117924 389156
rect 130476 389172 130528 389224
rect 168380 389172 168432 389224
rect 66076 389036 66128 389088
rect 74540 389036 74592 389088
rect 111616 388628 111668 388680
rect 112444 388628 112496 388680
rect 93400 388424 93452 388476
rect 100116 388424 100168 388476
rect 101404 388424 101456 388476
rect 120172 388424 120224 388476
rect 94688 387812 94740 387864
rect 64512 387744 64564 387796
rect 79140 387744 79192 387796
rect 93124 387744 93176 387796
rect 128452 387744 128504 387796
rect 78680 387268 78732 387320
rect 79140 387268 79192 387320
rect 60556 386316 60608 386368
rect 82084 386316 82136 386368
rect 110144 385636 110196 385688
rect 155224 385636 155276 385688
rect 56416 384956 56468 385008
rect 87052 384956 87104 385008
rect 104072 384956 104124 385008
rect 136640 384956 136692 385008
rect 137100 384956 137152 385008
rect 87052 384344 87104 384396
rect 88248 384344 88300 384396
rect 5448 384276 5500 384328
rect 123116 384276 123168 384328
rect 137100 384276 137152 384328
rect 169116 384276 169168 384328
rect 36544 382236 36596 382288
rect 118700 382236 118752 382288
rect 119436 382236 119488 382288
rect 88340 382168 88392 382220
rect 115112 382168 115164 382220
rect 115756 382168 115808 382220
rect 115756 380876 115808 380928
rect 130476 380876 130528 380928
rect 67640 380196 67692 380248
rect 123208 380196 123260 380248
rect 61752 380128 61804 380180
rect 158720 380128 158772 380180
rect 44088 379448 44140 379500
rect 75920 379448 75972 379500
rect 76564 379448 76616 379500
rect 63224 378768 63276 378820
rect 87604 378768 87656 378820
rect 67824 375980 67876 376032
rect 145564 375980 145616 376032
rect 67732 374620 67784 374672
rect 124956 374620 125008 374672
rect 150256 374076 150308 374128
rect 242164 374076 242216 374128
rect 57704 374008 57756 374060
rect 193864 374008 193916 374060
rect 107476 373260 107528 373312
rect 164240 373260 164292 373312
rect 150348 372580 150400 372632
rect 248512 372580 248564 372632
rect 137284 372172 137336 372224
rect 137928 372172 137980 372224
rect 70308 371832 70360 371884
rect 155960 371832 156012 371884
rect 137928 371220 137980 371272
rect 180800 371220 180852 371272
rect 133144 370540 133196 370592
rect 164884 370540 164936 370592
rect 64604 370472 64656 370524
rect 108304 370472 108356 370524
rect 108856 370472 108908 370524
rect 160744 370472 160796 370524
rect 121460 368908 121512 368960
rect 122104 368908 122156 368960
rect 85580 368568 85632 368620
rect 215392 368568 215444 368620
rect 62028 368500 62080 368552
rect 121460 368500 121512 368552
rect 144828 368500 144880 368552
rect 306748 368500 306800 368552
rect 119436 367752 119488 367804
rect 167000 367752 167052 367804
rect 126336 367072 126388 367124
rect 209044 367072 209096 367124
rect 86960 366324 87012 366376
rect 95240 366324 95292 366376
rect 99288 366324 99340 366376
rect 173256 366324 173308 366376
rect 102784 365712 102836 365764
rect 305000 365712 305052 365764
rect 81440 365644 81492 365696
rect 82084 365644 82136 365696
rect 71688 365236 71740 365288
rect 73160 365236 73212 365288
rect 136640 364420 136692 364472
rect 204904 364420 204956 364472
rect 81440 364352 81492 364404
rect 240508 364352 240560 364404
rect 122104 363604 122156 363656
rect 208124 363604 208176 363656
rect 100024 362924 100076 362976
rect 196624 362924 196676 362976
rect 147680 361632 147732 361684
rect 155592 361632 155644 361684
rect 107568 361564 107620 361616
rect 186964 361564 187016 361616
rect 124864 360272 124916 360324
rect 125600 360272 125652 360324
rect 128360 360272 128412 360324
rect 166448 360272 166500 360324
rect 120080 360204 120132 360256
rect 214564 360204 214616 360256
rect 132500 358844 132552 358896
rect 174728 358844 174780 358896
rect 88984 358776 89036 358828
rect 91192 358776 91244 358828
rect 213184 358776 213236 358828
rect 3332 358708 3384 358760
rect 36544 358708 36596 358760
rect 107844 358708 107896 358760
rect 108304 358708 108356 358760
rect 135904 357484 135956 357536
rect 192576 357484 192628 357536
rect 107844 357416 107896 357468
rect 241520 357416 241572 357468
rect 92388 356668 92440 356720
rect 121460 356668 121512 356720
rect 132408 356124 132460 356176
rect 176108 356124 176160 356176
rect 122840 356056 122892 356108
rect 225604 356056 225656 356108
rect 155592 355988 155644 356040
rect 159364 355988 159416 356040
rect 52276 355308 52328 355360
rect 93860 355308 93912 355360
rect 95148 355308 95200 355360
rect 97816 355308 97868 355360
rect 154672 355308 154724 355360
rect 51724 355036 51776 355088
rect 52276 355036 52328 355088
rect 123484 354696 123536 354748
rect 184296 354696 184348 354748
rect 93216 353948 93268 354000
rect 118792 353948 118844 354000
rect 122748 353948 122800 354000
rect 126336 353948 126388 354000
rect 132592 353336 132644 353388
rect 222936 353336 222988 353388
rect 61936 353268 61988 353320
rect 218704 353268 218756 353320
rect 104808 352588 104860 352640
rect 120724 352588 120776 352640
rect 83464 352520 83516 352572
rect 101404 352520 101456 352572
rect 105636 352520 105688 352572
rect 155316 352520 155368 352572
rect 144184 352248 144236 352300
rect 144736 352248 144788 352300
rect 144736 351908 144788 351960
rect 184388 351908 184440 351960
rect 79968 351228 80020 351280
rect 111064 351228 111116 351280
rect 67824 351160 67876 351212
rect 122840 351160 122892 351212
rect 118792 350548 118844 350600
rect 178776 350548 178828 350600
rect 112444 349800 112496 349852
rect 156052 349800 156104 349852
rect 129004 349120 129056 349172
rect 180064 349120 180116 349172
rect 117228 347828 117280 347880
rect 235264 347828 235316 347880
rect 89720 347760 89772 347812
rect 91008 347760 91060 347812
rect 255412 347760 255464 347812
rect 3424 347012 3476 347064
rect 78680 347012 78732 347064
rect 124128 347012 124180 347064
rect 140780 347012 140832 347064
rect 122932 346944 122984 346996
rect 142804 346468 142856 346520
rect 162124 346468 162176 346520
rect 101956 346400 102008 346452
rect 221464 346400 221516 346452
rect 3148 346332 3200 346384
rect 7564 346332 7616 346384
rect 74448 345652 74500 345704
rect 89720 345652 89772 345704
rect 129832 345108 129884 345160
rect 231124 345108 231176 345160
rect 84200 345040 84252 345092
rect 85488 345040 85540 345092
rect 195244 345040 195296 345092
rect 90916 343680 90968 343732
rect 211804 343680 211856 343732
rect 77208 343612 77260 343664
rect 204352 343612 204404 343664
rect 79876 342864 79928 342916
rect 88984 342864 89036 342916
rect 105544 342320 105596 342372
rect 220084 342320 220136 342372
rect 93676 342252 93728 342304
rect 251180 342252 251232 342304
rect 75828 341504 75880 341556
rect 101496 341504 101548 341556
rect 142896 340960 142948 341012
rect 160928 340960 160980 341012
rect 102692 340892 102744 340944
rect 258172 340892 258224 340944
rect 77300 340212 77352 340264
rect 93124 340212 93176 340264
rect 64604 340144 64656 340196
rect 72424 340144 72476 340196
rect 134524 340144 134576 340196
rect 114468 339532 114520 339584
rect 177488 339532 177540 339584
rect 134248 339464 134300 339516
rect 236644 339464 236696 339516
rect 77116 338716 77168 338768
rect 87604 338716 87656 338768
rect 106464 338172 106516 338224
rect 191196 338172 191248 338224
rect 85672 338104 85724 338156
rect 249984 338104 250036 338156
rect 63408 336812 63460 336864
rect 163596 336812 163648 336864
rect 115940 336744 115992 336796
rect 247316 336744 247368 336796
rect 66076 335996 66128 336048
rect 74540 335996 74592 336048
rect 104900 335384 104952 335436
rect 228456 335384 228508 335436
rect 67180 335316 67232 335368
rect 206376 335316 206428 335368
rect 65984 334568 66036 334620
rect 142896 334568 142948 334620
rect 144460 334024 144512 334076
rect 160836 334024 160888 334076
rect 146208 333956 146260 334008
rect 171784 333956 171836 334008
rect 67364 332596 67416 332648
rect 67548 332596 67600 332648
rect 115020 332664 115072 332716
rect 141424 332664 141476 332716
rect 158812 332664 158864 332716
rect 115664 332596 115716 332648
rect 169208 332596 169260 332648
rect 86316 331848 86368 331900
rect 97264 331848 97316 331900
rect 102508 331304 102560 331356
rect 164976 331304 165028 331356
rect 49608 331236 49660 331288
rect 83740 331236 83792 331288
rect 97908 331236 97960 331288
rect 215944 331236 215996 331288
rect 159364 331168 159416 331220
rect 161756 331168 161808 331220
rect 76472 331100 76524 331152
rect 77116 331100 77168 331152
rect 95332 331100 95384 331152
rect 95884 331100 95936 331152
rect 101496 331100 101548 331152
rect 101956 331100 102008 331152
rect 107568 331100 107620 331152
rect 108028 331100 108080 331152
rect 114376 331100 114428 331152
rect 116584 331100 116636 331152
rect 117780 331100 117832 331152
rect 118608 331100 118660 331152
rect 118700 331100 118752 331152
rect 119436 331100 119488 331152
rect 122840 331100 122892 331152
rect 123668 331100 123720 331152
rect 125600 331100 125652 331152
rect 126428 331100 126480 331152
rect 137928 331100 137980 331152
rect 139400 331100 139452 331152
rect 144184 331100 144236 331152
rect 144828 331100 144880 331152
rect 95792 331032 95844 331084
rect 96528 331032 96580 331084
rect 140688 331032 140740 331084
rect 142804 331032 142856 331084
rect 144736 331032 144788 331084
rect 146484 331032 146536 331084
rect 108304 330828 108356 330880
rect 115204 330828 115256 330880
rect 196716 330556 196768 330608
rect 251364 330556 251416 330608
rect 72240 330488 72292 330540
rect 97908 330488 97960 330540
rect 115020 330488 115072 330540
rect 140780 330488 140832 330540
rect 162124 330488 162176 330540
rect 239496 330488 239548 330540
rect 110604 330352 110656 330404
rect 111708 330352 111760 330404
rect 104256 330080 104308 330132
rect 105544 330080 105596 330132
rect 127716 330080 127768 330132
rect 129004 330080 129056 330132
rect 100024 330012 100076 330064
rect 102784 330012 102836 330064
rect 79416 329944 79468 329996
rect 79968 329944 80020 329996
rect 113640 329944 113692 329996
rect 114468 329944 114520 329996
rect 153660 329876 153712 329928
rect 159456 329876 159508 329928
rect 44088 329808 44140 329860
rect 69112 329808 69164 329860
rect 91100 329808 91152 329860
rect 111892 329808 111944 329860
rect 134156 329808 134208 329860
rect 135076 329808 135128 329860
rect 135260 329808 135312 329860
rect 135812 329808 135864 329860
rect 151636 329808 151688 329860
rect 195428 329808 195480 329860
rect 134524 329128 134576 329180
rect 196716 329128 196768 329180
rect 43444 329060 43496 329112
rect 49516 329060 49568 329112
rect 135260 329060 135312 329112
rect 160928 329060 160980 329112
rect 224224 329060 224276 329112
rect 36544 328448 36596 328500
rect 124864 328448 124916 328500
rect 152096 328448 152148 328500
rect 161020 328448 161072 328500
rect 213184 327768 213236 327820
rect 248604 327768 248656 327820
rect 60556 327700 60608 327752
rect 91100 327700 91152 327752
rect 158812 327700 158864 327752
rect 185676 327700 185728 327752
rect 187056 327700 187108 327752
rect 331220 327700 331272 327752
rect 33784 327156 33836 327208
rect 114744 327156 114796 327208
rect 149888 327156 149940 327208
rect 153660 327156 153712 327208
rect 154304 327156 154356 327208
rect 158168 327156 158220 327208
rect 91560 327088 91612 327140
rect 92388 327088 92440 327140
rect 180156 327088 180208 327140
rect 70032 327020 70084 327072
rect 71044 327020 71096 327072
rect 139768 327020 139820 327072
rect 151636 327020 151688 327072
rect 152832 326952 152884 327004
rect 154212 326952 154264 327004
rect 68652 326884 68704 326936
rect 71412 326884 71464 326936
rect 143448 326884 143500 326936
rect 149152 326884 149204 326936
rect 162216 326884 162268 326936
rect 66812 326816 66864 326868
rect 68008 326816 68060 326868
rect 20 326340 72 326392
rect 51724 326340 51776 326392
rect 161756 326340 161808 326392
rect 177304 326340 177356 326392
rect 240784 325728 240836 325780
rect 59176 325660 59228 325712
rect 68100 325660 68152 325712
rect 161020 324980 161072 325032
rect 258356 324980 258408 325032
rect 156052 324912 156104 324964
rect 255504 324912 255556 324964
rect 56508 324300 56560 324352
rect 66904 324300 66956 324352
rect 156144 324232 156196 324284
rect 164240 324232 164292 324284
rect 172060 324232 172112 324284
rect 162308 323552 162360 323604
rect 349160 323552 349212 323604
rect 156052 323416 156104 323468
rect 162584 323416 162636 323468
rect 59268 322940 59320 322992
rect 66720 322940 66772 322992
rect 154764 322532 154816 322584
rect 155316 322532 155368 322584
rect 156052 321920 156104 321972
rect 163504 321920 163556 321972
rect 54944 321580 54996 321632
rect 64144 321580 64196 321632
rect 154764 321580 154816 321632
rect 243820 321580 243872 321632
rect 66628 321512 66680 321564
rect 222936 320968 222988 321020
rect 252652 320968 252704 321020
rect 204904 320900 204956 320952
rect 238116 320900 238168 320952
rect 163596 320832 163648 320884
rect 223028 320832 223080 320884
rect 156604 320152 156656 320204
rect 195152 320152 195204 320204
rect 157248 319472 157300 319524
rect 160100 319472 160152 319524
rect 199384 319472 199436 319524
rect 4068 319404 4120 319456
rect 5448 319404 5500 319456
rect 29644 319404 29696 319456
rect 162584 319404 162636 319456
rect 210424 319404 210476 319456
rect 64420 318792 64472 318844
rect 66904 318792 66956 318844
rect 157248 318792 157300 318844
rect 162124 318792 162176 318844
rect 210424 318792 210476 318844
rect 258080 318792 258132 318844
rect 186964 318112 187016 318164
rect 227628 318112 227680 318164
rect 3516 318044 3568 318096
rect 46848 318044 46900 318096
rect 158168 318044 158220 318096
rect 189908 318044 189960 318096
rect 195428 318044 195480 318096
rect 242256 318044 242308 318096
rect 60648 317500 60700 317552
rect 66904 317500 66956 317552
rect 46848 317432 46900 317484
rect 66720 317432 66772 317484
rect 157248 316752 157300 316804
rect 188436 316752 188488 316804
rect 166540 316684 166592 316736
rect 305644 316684 305696 316736
rect 64788 315664 64840 315716
rect 66996 315664 67048 315716
rect 155960 315324 156012 315376
rect 171968 315324 172020 315376
rect 172060 315324 172112 315376
rect 192484 315324 192536 315376
rect 163688 315256 163740 315308
rect 244280 315256 244332 315308
rect 35164 314644 35216 314696
rect 67548 314644 67600 314696
rect 217324 314644 217376 314696
rect 217968 314644 218020 314696
rect 302240 314644 302292 314696
rect 178776 313964 178828 314016
rect 235540 313964 235592 314016
rect 198096 313896 198148 313948
rect 320180 313896 320232 313948
rect 61844 313284 61896 313336
rect 65524 313284 65576 313336
rect 61936 313216 61988 313268
rect 66904 313216 66956 313268
rect 166448 312604 166500 312656
rect 230480 312604 230532 312656
rect 157340 312536 157392 312588
rect 245660 312536 245712 312588
rect 157248 311856 157300 311908
rect 166540 311856 166592 311908
rect 63408 311788 63460 311840
rect 66904 311788 66956 311840
rect 214564 311176 214616 311228
rect 227812 311176 227864 311228
rect 174728 311108 174780 311160
rect 233976 311108 234028 311160
rect 157248 310496 157300 310548
rect 166448 310496 166500 310548
rect 165068 309748 165120 309800
rect 198096 309748 198148 309800
rect 198004 309204 198056 309256
rect 198648 309204 198700 309256
rect 265624 309204 265676 309256
rect 63224 309136 63276 309188
rect 66628 309136 66680 309188
rect 167736 309136 167788 309188
rect 260840 309136 260892 309188
rect 50804 308388 50856 308440
rect 67088 308388 67140 308440
rect 207664 307844 207716 307896
rect 286324 307844 286376 307896
rect 11704 307776 11756 307828
rect 50804 307776 50856 307828
rect 195336 307776 195388 307828
rect 201684 307776 201736 307828
rect 583484 307776 583536 307828
rect 64604 307708 64656 307760
rect 66536 307708 66588 307760
rect 22744 307028 22796 307080
rect 67088 307028 67140 307080
rect 211804 306416 211856 306468
rect 280896 306416 280948 306468
rect 156512 306348 156564 306400
rect 318064 306348 318116 306400
rect 3516 306280 3568 306332
rect 43444 306280 43496 306332
rect 64696 306280 64748 306332
rect 66904 306280 66956 306332
rect 157248 306280 157300 306332
rect 158720 306280 158772 306332
rect 162124 305600 162176 305652
rect 245752 305600 245804 305652
rect 157248 305192 157300 305244
rect 162308 305192 162360 305244
rect 198096 304988 198148 305040
rect 198556 304988 198608 305040
rect 295340 304988 295392 305040
rect 221188 303696 221240 303748
rect 271236 303696 271288 303748
rect 57888 303628 57940 303680
rect 66904 303628 66956 303680
rect 156052 303628 156104 303680
rect 213184 303628 213236 303680
rect 214748 303628 214800 303680
rect 565084 303628 565136 303680
rect 60464 303560 60516 303612
rect 66996 303560 67048 303612
rect 158720 302880 158772 302932
rect 191196 302880 191248 302932
rect 220084 302268 220136 302320
rect 220728 302268 220780 302320
rect 298192 302268 298244 302320
rect 157248 302200 157300 302252
rect 244004 302200 244056 302252
rect 199476 302132 199528 302184
rect 201408 302132 201460 302184
rect 166356 300908 166408 300960
rect 208400 300908 208452 300960
rect 156788 300840 156840 300892
rect 188344 300840 188396 300892
rect 201408 300840 201460 300892
rect 276664 300840 276716 300892
rect 193956 299548 194008 299600
rect 258264 299548 258316 299600
rect 56416 299480 56468 299532
rect 66904 299480 66956 299532
rect 157156 299480 157208 299532
rect 244924 299480 244976 299532
rect 157248 299412 157300 299464
rect 167000 299412 167052 299464
rect 169208 298800 169260 298852
rect 186964 298800 187016 298852
rect 167000 298732 167052 298784
rect 225328 298732 225380 298784
rect 228364 298732 228416 298784
rect 236184 298732 236236 298784
rect 195336 298188 195388 298240
rect 252744 298188 252796 298240
rect 236184 298120 236236 298172
rect 574744 298120 574796 298172
rect 236092 297304 236144 297356
rect 236644 297304 236696 297356
rect 236644 296760 236696 296812
rect 282920 296760 282972 296812
rect 163504 296692 163556 296744
rect 238484 296692 238536 296744
rect 57704 296624 57756 296676
rect 66904 296624 66956 296676
rect 156420 295944 156472 295996
rect 244372 295944 244424 295996
rect 160008 295332 160060 295384
rect 161572 295332 161624 295384
rect 196808 295332 196860 295384
rect 259552 295332 259604 295384
rect 156328 295264 156380 295316
rect 166356 295264 166408 295316
rect 166540 294584 166592 294636
rect 245936 294584 245988 294636
rect 154856 293972 154908 294024
rect 248696 293972 248748 294024
rect 59084 293904 59136 293956
rect 66996 293904 67048 293956
rect 213184 293224 213236 293276
rect 236000 293224 236052 293276
rect 2780 292816 2832 292868
rect 4804 292816 4856 292868
rect 48044 292544 48096 292596
rect 66720 292544 66772 292596
rect 157248 292544 157300 292596
rect 220636 292544 220688 292596
rect 255320 292544 255372 292596
rect 14464 292476 14516 292528
rect 62028 292476 62080 292528
rect 66904 292476 66956 292528
rect 162216 291796 162268 291848
rect 173440 291796 173492 291848
rect 201408 291796 201460 291848
rect 218060 291796 218112 291848
rect 217876 291252 217928 291304
rect 218152 291252 218204 291304
rect 233976 291252 234028 291304
rect 289912 291252 289964 291304
rect 156788 291184 156840 291236
rect 159640 291184 159692 291236
rect 167828 291184 167880 291236
rect 256792 291184 256844 291236
rect 200396 291116 200448 291168
rect 204260 291116 204312 291168
rect 582564 291116 582616 291168
rect 239404 291048 239456 291100
rect 242348 291048 242400 291100
rect 182916 290436 182968 290488
rect 193956 290436 194008 290488
rect 197360 290436 197412 290488
rect 239956 290436 240008 290488
rect 63316 289892 63368 289944
rect 66904 289892 66956 289944
rect 242348 289824 242400 289876
rect 264244 289824 264296 289876
rect 232504 289756 232556 289808
rect 234620 289756 234672 289808
rect 242164 289756 242216 289808
rect 242900 289756 242952 289808
rect 60556 289348 60608 289400
rect 66904 289348 66956 289400
rect 52184 289076 52236 289128
rect 67180 289076 67232 289128
rect 187148 288464 187200 288516
rect 230572 288464 230624 288516
rect 156788 288396 156840 288448
rect 224500 288396 224552 288448
rect 237932 288396 237984 288448
rect 238116 288396 238168 288448
rect 264336 288396 264388 288448
rect 156236 287104 156288 287156
rect 231308 287104 231360 287156
rect 238116 287104 238168 287156
rect 267096 287104 267148 287156
rect 64696 287036 64748 287088
rect 66720 287036 66772 287088
rect 156328 287036 156380 287088
rect 244464 287036 244516 287088
rect 240784 286492 240836 286544
rect 241980 286492 242032 286544
rect 217968 286424 218020 286476
rect 221556 286424 221608 286476
rect 224224 286220 224276 286272
rect 225052 286220 225104 286272
rect 63408 285744 63460 285796
rect 66904 285744 66956 285796
rect 199384 285744 199436 285796
rect 205548 285744 205600 285796
rect 213828 285744 213880 285796
rect 215392 285744 215444 285796
rect 55128 285676 55180 285728
rect 66812 285676 66864 285728
rect 157248 285676 157300 285728
rect 166356 285676 166408 285728
rect 169300 285676 169352 285728
rect 173256 285676 173308 285728
rect 194048 285676 194100 285728
rect 204628 285676 204680 285728
rect 206376 285676 206428 285728
rect 207020 285676 207072 285728
rect 214564 285676 214616 285728
rect 223580 285744 223632 285796
rect 227628 285744 227680 285796
rect 228916 285744 228968 285796
rect 231124 285744 231176 285796
rect 232228 285744 232280 285796
rect 251824 285744 251876 285796
rect 219716 285676 219768 285728
rect 220728 285676 220780 285728
rect 222844 285676 222896 285728
rect 226524 285676 226576 285728
rect 228456 285676 228508 285728
rect 229284 285676 229336 285728
rect 233148 285676 233200 285728
rect 233884 285676 233936 285728
rect 200120 285268 200172 285320
rect 200488 285268 200540 285320
rect 208400 285268 208452 285320
rect 208676 285268 208728 285320
rect 218152 285268 218204 285320
rect 218336 285268 218388 285320
rect 192576 284928 192628 284980
rect 214564 284928 214616 284980
rect 216772 284384 216824 284436
rect 248420 284384 248472 284436
rect 157248 284316 157300 284368
rect 247040 284316 247092 284368
rect 180156 284248 180208 284300
rect 197360 284248 197412 284300
rect 242256 283908 242308 283960
rect 313280 283840 313332 283892
rect 177304 283568 177356 283620
rect 185768 283568 185820 283620
rect 246396 283568 246448 283620
rect 247316 283568 247368 283620
rect 252836 283568 252888 283620
rect 39948 282888 40000 282940
rect 66720 282888 66772 282940
rect 157248 282888 157300 282940
rect 179512 282888 179564 282940
rect 157156 282820 157208 282872
rect 182916 282820 182968 282872
rect 246120 282820 246172 282872
rect 252560 282820 252612 282872
rect 582748 282820 582800 282872
rect 179512 282140 179564 282192
rect 180708 282140 180760 282192
rect 197360 282140 197412 282192
rect 245936 281664 245988 281716
rect 250076 281664 250128 281716
rect 52276 281528 52328 281580
rect 66352 281528 66404 281580
rect 157248 281460 157300 281512
rect 196808 281460 196860 281512
rect 246120 281460 246172 281512
rect 258356 281460 258408 281512
rect 259368 281460 259420 281512
rect 171876 281392 171928 281444
rect 177304 281392 177356 281444
rect 191196 281392 191248 281444
rect 197360 281392 197412 281444
rect 259368 280848 259420 280900
rect 271144 280848 271196 280900
rect 157064 280780 157116 280832
rect 167828 280780 167880 280832
rect 245936 280780 245988 280832
rect 248512 280780 248564 280832
rect 273904 280780 273956 280832
rect 59084 280168 59136 280220
rect 66812 280168 66864 280220
rect 245936 279828 245988 279880
rect 249892 279828 249944 279880
rect 251088 279828 251140 279880
rect 162308 279420 162360 279472
rect 191748 279420 191800 279472
rect 197452 279420 197504 279472
rect 251088 279420 251140 279472
rect 583576 279420 583628 279472
rect 157248 279012 157300 279064
rect 161388 279012 161440 279064
rect 156972 278808 157024 278860
rect 160100 278808 160152 278860
rect 14464 278740 14516 278792
rect 60464 278740 60516 278792
rect 67272 278740 67324 278792
rect 245936 278672 245988 278724
rect 254124 278672 254176 278724
rect 181444 277992 181496 278044
rect 197360 277992 197412 278044
rect 254124 277992 254176 278044
rect 583300 277992 583352 278044
rect 191840 277788 191892 277840
rect 197452 277788 197504 277840
rect 54852 277380 54904 277432
rect 66720 277380 66772 277432
rect 157248 277380 157300 277432
rect 166540 277380 166592 277432
rect 186964 277380 187016 277432
rect 191840 277380 191892 277432
rect 185768 276700 185820 276752
rect 197544 276700 197596 276752
rect 160100 276632 160152 276684
rect 194508 276632 194560 276684
rect 197360 276632 197412 276684
rect 245752 276632 245804 276684
rect 278044 276632 278096 276684
rect 177488 276496 177540 276548
rect 181536 276496 181588 276548
rect 156880 276020 156932 276072
rect 167828 276020 167880 276072
rect 245936 275952 245988 276004
rect 253940 275952 253992 276004
rect 582656 275952 582708 276004
rect 186964 275340 187016 275392
rect 199660 275340 199712 275392
rect 166448 275272 166500 275324
rect 188620 275272 188672 275324
rect 61752 274660 61804 274712
rect 66812 274660 66864 274712
rect 162216 274660 162268 274712
rect 169300 274660 169352 274712
rect 156512 274592 156564 274644
rect 167736 274592 167788 274644
rect 264336 273980 264388 274032
rect 280804 273980 280856 274032
rect 57704 273912 57756 273964
rect 66904 273912 66956 273964
rect 159456 273912 159508 273964
rect 187148 273912 187200 273964
rect 245844 273912 245896 273964
rect 311900 273912 311952 273964
rect 62028 273232 62080 273284
rect 66812 273232 66864 273284
rect 187056 273232 187108 273284
rect 197360 273232 197412 273284
rect 245844 273232 245896 273284
rect 249892 273232 249944 273284
rect 164976 272552 165028 272604
rect 177488 272552 177540 272604
rect 165068 272484 165120 272536
rect 197452 272484 197504 272536
rect 245752 272484 245804 272536
rect 252652 272484 252704 272536
rect 253848 272484 253900 272536
rect 176108 271804 176160 271856
rect 182916 271804 182968 271856
rect 197360 271872 197412 271924
rect 245844 271464 245896 271516
rect 248604 271464 248656 271516
rect 157156 271124 157208 271176
rect 191196 271124 191248 271176
rect 195520 270580 195572 270632
rect 197820 270580 197872 270632
rect 48228 270512 48280 270564
rect 66904 270512 66956 270564
rect 157248 270512 157300 270564
rect 175924 270512 175976 270564
rect 186228 270512 186280 270564
rect 197360 270512 197412 270564
rect 245936 270444 245988 270496
rect 251180 270444 251232 270496
rect 252652 270444 252704 270496
rect 256884 270444 256936 270496
rect 583392 270444 583444 270496
rect 194876 269832 194928 269884
rect 197452 269832 197504 269884
rect 246580 269764 246632 269816
rect 256884 269764 256936 269816
rect 181628 269152 181680 269204
rect 197360 269152 197412 269204
rect 64512 269084 64564 269136
rect 66720 269084 66772 269136
rect 157248 269084 157300 269136
rect 195428 269084 195480 269136
rect 171968 269016 172020 269068
rect 197360 269016 197412 269068
rect 245752 269016 245804 269068
rect 263600 269016 263652 269068
rect 157248 268336 157300 268388
rect 192576 268336 192628 268388
rect 263600 268336 263652 268388
rect 582656 268336 582708 268388
rect 38660 267724 38712 267776
rect 40684 267724 40736 267776
rect 157248 267656 157300 267708
rect 195336 267656 195388 267708
rect 38660 267588 38712 267640
rect 43444 267588 43496 267640
rect 3516 266976 3568 267028
rect 38660 266976 38712 267028
rect 159640 266976 159692 267028
rect 193956 266976 194008 267028
rect 246488 266976 246540 267028
rect 294052 266976 294104 267028
rect 195888 266364 195940 266416
rect 198004 266364 198056 266416
rect 245844 266364 245896 266416
rect 276020 266364 276072 266416
rect 157248 266296 157300 266348
rect 198096 266296 198148 266348
rect 245936 266296 245988 266348
rect 267740 266296 267792 266348
rect 269028 266296 269080 266348
rect 191104 266228 191156 266280
rect 197360 266228 197412 266280
rect 245936 265752 245988 265804
rect 249984 265752 250036 265804
rect 269028 265616 269080 265668
rect 583024 265616 583076 265668
rect 41328 264936 41380 264988
rect 66812 264936 66864 264988
rect 50988 264188 51040 264240
rect 65984 264188 66036 264240
rect 66536 264188 66588 264240
rect 156880 264188 156932 264240
rect 174728 264188 174780 264240
rect 189908 264188 189960 264240
rect 199568 264188 199620 264240
rect 246028 264188 246080 264240
rect 296720 264188 296772 264240
rect 56324 263576 56376 263628
rect 66812 263576 66864 263628
rect 164148 263576 164200 263628
rect 197360 263576 197412 263628
rect 247132 263304 247184 263356
rect 247040 263100 247092 263152
rect 52368 262828 52420 262880
rect 63500 262828 63552 262880
rect 169300 262828 169352 262880
rect 185676 262828 185728 262880
rect 246672 262828 246724 262880
rect 310612 262828 310664 262880
rect 63500 262216 63552 262268
rect 64604 262216 64656 262268
rect 66444 262216 66496 262268
rect 157248 262216 157300 262268
rect 178776 262216 178828 262268
rect 185768 262216 185820 262268
rect 197360 262216 197412 262268
rect 245936 262216 245988 262268
rect 251456 262216 251508 262268
rect 160928 261536 160980 261588
rect 169760 261536 169812 261588
rect 189908 261536 189960 261588
rect 199384 261536 199436 261588
rect 29644 261468 29696 261520
rect 52460 261468 52512 261520
rect 167736 261468 167788 261520
rect 195520 261468 195572 261520
rect 246396 261468 246448 261520
rect 247316 261468 247368 261520
rect 251180 261468 251232 261520
rect 251824 261468 251876 261520
rect 281908 261468 281960 261520
rect 52460 260856 52512 260908
rect 53472 260856 53524 260908
rect 66812 260856 66864 260908
rect 245936 260176 245988 260228
rect 248696 260176 248748 260228
rect 160836 260108 160888 260160
rect 171968 260108 172020 260160
rect 60556 259428 60608 259480
rect 66812 259428 66864 259480
rect 188528 259428 188580 259480
rect 197452 259428 197504 259480
rect 244372 259428 244424 259480
rect 291200 259428 291252 259480
rect 184296 259360 184348 259412
rect 197360 259360 197412 259412
rect 245936 259360 245988 259412
rect 259552 259360 259604 259412
rect 260748 259360 260800 259412
rect 171876 258680 171928 258732
rect 197912 258680 197964 258732
rect 260748 258680 260800 258732
rect 300952 258680 301004 258732
rect 53748 258068 53800 258120
rect 66720 258068 66772 258120
rect 156420 258068 156472 258120
rect 170496 258068 170548 258120
rect 67456 258000 67508 258052
rect 68192 258000 68244 258052
rect 156880 257932 156932 257984
rect 159548 257932 159600 257984
rect 198648 257456 198700 257508
rect 199384 257456 199436 257508
rect 195428 257388 195480 257440
rect 200028 257388 200080 257440
rect 260196 257320 260248 257372
rect 580356 257320 580408 257372
rect 157248 256776 157300 256828
rect 177948 256776 178000 256828
rect 181444 256776 181496 256828
rect 158720 256708 158772 256760
rect 184848 256708 184900 256760
rect 197360 256776 197412 256828
rect 188436 256640 188488 256692
rect 197360 256640 197412 256692
rect 192576 256368 192628 256420
rect 193864 256368 193916 256420
rect 245660 256028 245712 256080
rect 260840 256028 260892 256080
rect 247132 255960 247184 256012
rect 288440 255960 288492 256012
rect 60372 255688 60424 255740
rect 66996 255688 67048 255740
rect 157248 255280 157300 255332
rect 168380 255280 168432 255332
rect 3148 255212 3200 255264
rect 11704 255212 11756 255264
rect 178040 255212 178092 255264
rect 195980 255212 196032 255264
rect 159548 254532 159600 254584
rect 178040 254532 178092 254584
rect 260840 254532 260892 254584
rect 295432 254532 295484 254584
rect 63132 253920 63184 253972
rect 66904 253920 66956 253972
rect 157248 253920 157300 253972
rect 179328 253920 179380 253972
rect 192668 253920 192720 253972
rect 197360 253920 197412 253972
rect 245936 253852 245988 253904
rect 258264 253852 258316 253904
rect 259368 253852 259420 253904
rect 156420 253580 156472 253632
rect 158720 253580 158772 253632
rect 177488 253240 177540 253292
rect 186320 253240 186372 253292
rect 158168 253172 158220 253224
rect 165160 253172 165212 253224
rect 166540 253172 166592 253224
rect 180340 253172 180392 253224
rect 245660 253172 245712 253224
rect 256792 253172 256844 253224
rect 259368 253172 259420 253224
rect 296812 253172 296864 253224
rect 186320 252628 186372 252680
rect 187608 252628 187660 252680
rect 197452 252628 197504 252680
rect 55036 252560 55088 252612
rect 57612 252560 57664 252612
rect 66904 252560 66956 252612
rect 179880 252560 179932 252612
rect 197360 252560 197412 252612
rect 246028 252492 246080 252544
rect 259460 252492 259512 252544
rect 260748 252492 260800 252544
rect 245936 252424 245988 252476
rect 251364 252424 251416 252476
rect 58992 252084 59044 252136
rect 66812 252084 66864 252136
rect 159364 251880 159416 251932
rect 170404 251880 170456 251932
rect 168380 251812 168432 251864
rect 195796 251812 195848 251864
rect 197452 251812 197504 251864
rect 260748 251812 260800 251864
rect 583668 251812 583720 251864
rect 156880 251336 156932 251388
rect 162216 251336 162268 251388
rect 191104 251200 191156 251252
rect 197360 251200 197412 251252
rect 245660 250452 245712 250504
rect 252744 250452 252796 250504
rect 253020 250452 253072 250504
rect 256792 250452 256844 250504
rect 287060 250452 287112 250504
rect 164148 249840 164200 249892
rect 169024 249840 169076 249892
rect 185676 249840 185728 249892
rect 197360 249840 197412 249892
rect 157248 249772 157300 249824
rect 196348 249772 196400 249824
rect 157156 249704 157208 249756
rect 164148 249704 164200 249756
rect 167828 249704 167880 249756
rect 169208 249704 169260 249756
rect 191196 249704 191248 249756
rect 195704 249704 195756 249756
rect 197360 249704 197412 249756
rect 178868 249296 178920 249348
rect 179880 249296 179932 249348
rect 169760 249024 169812 249076
rect 199476 249024 199528 249076
rect 253020 249024 253072 249076
rect 285680 249024 285732 249076
rect 61936 248412 61988 248464
rect 66812 248412 66864 248464
rect 156420 248412 156472 248464
rect 177856 248412 177908 248464
rect 67456 248276 67508 248328
rect 67916 248276 67968 248328
rect 171784 247732 171836 247784
rect 194416 247732 194468 247784
rect 158628 247664 158680 247716
rect 182732 247664 182784 247716
rect 245936 247664 245988 247716
rect 248696 247664 248748 247716
rect 582840 247664 582892 247716
rect 50988 247052 51040 247104
rect 66628 247052 66680 247104
rect 191196 247052 191248 247104
rect 197452 247052 197504 247104
rect 195244 246984 195296 247036
rect 197360 246984 197412 247036
rect 245936 246372 245988 246424
rect 254032 246372 254084 246424
rect 245016 246304 245068 246356
rect 306564 246304 306616 246356
rect 194508 246032 194560 246084
rect 195336 246032 195388 246084
rect 156788 245692 156840 245744
rect 185768 245692 185820 245744
rect 154856 245624 154908 245676
rect 187056 245624 187108 245676
rect 254032 245624 254084 245676
rect 254584 245624 254636 245676
rect 53564 245556 53616 245608
rect 66628 245556 66680 245608
rect 190368 245420 190420 245472
rect 191840 245420 191892 245472
rect 194416 245148 194468 245200
rect 197360 245148 197412 245200
rect 196348 245012 196400 245064
rect 198740 245012 198792 245064
rect 177856 244876 177908 244928
rect 190000 244876 190052 244928
rect 280896 244876 280948 244928
rect 310520 244876 310572 244928
rect 155316 244332 155368 244384
rect 156972 244264 157024 244316
rect 160836 244264 160888 244316
rect 192576 244264 192628 244316
rect 192760 244264 192812 244316
rect 155408 243380 155460 243432
rect 155868 243380 155920 243432
rect 155868 242972 155920 243024
rect 174636 242972 174688 243024
rect 156052 242904 156104 242956
rect 188436 242904 188488 242956
rect 245936 242904 245988 242956
rect 271328 242904 271380 242956
rect 265624 242224 265676 242276
rect 278872 242224 278924 242276
rect 67456 242020 67508 242072
rect 73896 242020 73948 242072
rect 150072 242020 150124 242072
rect 169760 242156 169812 242208
rect 173808 242156 173860 242208
rect 197360 242156 197412 242208
rect 271236 242156 271288 242208
rect 298284 242156 298336 242208
rect 70308 241884 70360 241936
rect 76380 241884 76432 241936
rect 3516 241408 3568 241460
rect 36544 241408 36596 241460
rect 43444 241408 43496 241460
rect 92894 241408 92946 241460
rect 144230 241408 144282 241460
rect 192760 241476 192812 241528
rect 246396 241476 246448 241528
rect 247224 241476 247276 241528
rect 268384 241476 268436 241528
rect 106096 240796 106148 240848
rect 124864 240796 124916 240848
rect 152464 240796 152516 240848
rect 162308 240796 162360 240848
rect 67548 240728 67600 240780
rect 74724 240728 74776 240780
rect 82544 240728 82596 240780
rect 116584 240728 116636 240780
rect 138848 240728 138900 240780
rect 147680 240728 147732 240780
rect 149520 240728 149572 240780
rect 195704 240456 195756 240508
rect 200120 240456 200172 240508
rect 69020 240116 69072 240168
rect 69756 240116 69808 240168
rect 115940 240116 115992 240168
rect 116860 240116 116912 240168
rect 120724 240116 120776 240168
rect 136088 240116 136140 240168
rect 198648 240116 198700 240168
rect 200304 240116 200356 240168
rect 218152 240116 218204 240168
rect 224960 240116 225012 240168
rect 227812 240116 227864 240168
rect 242808 240116 242860 240168
rect 302332 240116 302384 240168
rect 68928 240048 68980 240100
rect 71412 240048 71464 240100
rect 76564 240048 76616 240100
rect 77300 240048 77352 240100
rect 86040 240048 86092 240100
rect 86868 240048 86920 240100
rect 90456 240048 90508 240100
rect 90916 240048 90968 240100
rect 91928 240048 91980 240100
rect 92388 240048 92440 240100
rect 99380 240048 99432 240100
rect 100668 240048 100720 240100
rect 115296 240048 115348 240100
rect 115848 240048 115900 240100
rect 120448 240048 120500 240100
rect 121368 240048 121420 240100
rect 121736 240048 121788 240100
rect 122748 240048 122800 240100
rect 124680 240048 124732 240100
rect 125416 240048 125468 240100
rect 126980 240048 127032 240100
rect 127532 240048 127584 240100
rect 130384 240048 130436 240100
rect 130936 240048 130988 240100
rect 131856 240048 131908 240100
rect 132408 240048 132460 240100
rect 134616 240048 134668 240100
rect 135168 240048 135220 240100
rect 138020 240048 138072 240100
rect 138940 240048 138992 240100
rect 144000 240048 144052 240100
rect 144828 240048 144880 240100
rect 147680 240048 147732 240100
rect 165068 240048 165120 240100
rect 242256 240048 242308 240100
rect 245660 240048 245712 240100
rect 74816 239980 74868 240032
rect 83464 239980 83516 240032
rect 127440 239980 127492 240032
rect 128268 239980 128320 240032
rect 106832 239912 106884 239964
rect 107568 239912 107620 239964
rect 111064 239912 111116 239964
rect 111616 239912 111668 239964
rect 121000 239912 121052 239964
rect 122932 239912 122984 239964
rect 133144 239912 133196 239964
rect 133788 239912 133840 239964
rect 142252 239912 142304 239964
rect 143448 239912 143500 239964
rect 88984 239776 89036 239828
rect 89628 239776 89680 239828
rect 148232 239776 148284 239828
rect 148968 239776 149020 239828
rect 71688 239640 71740 239692
rect 73804 239640 73856 239692
rect 75368 239640 75420 239692
rect 75828 239640 75880 239692
rect 101128 239640 101180 239692
rect 102048 239640 102100 239692
rect 149060 239572 149112 239624
rect 149612 239572 149664 239624
rect 79048 239504 79100 239556
rect 79968 239504 80020 239556
rect 141056 239504 141108 239556
rect 142068 239504 142120 239556
rect 200120 239504 200172 239556
rect 236736 239504 236788 239556
rect 198740 239436 198792 239488
rect 238760 239436 238812 239488
rect 81808 239368 81860 239420
rect 82728 239368 82780 239420
rect 84752 239368 84804 239420
rect 200120 239368 200172 239420
rect 80520 239232 80572 239284
rect 81256 239232 81308 239284
rect 109592 239232 109644 239284
rect 110328 239232 110380 239284
rect 128912 239232 128964 239284
rect 129648 239232 129700 239284
rect 153936 239232 153988 239284
rect 154488 239232 154540 239284
rect 69480 238824 69532 238876
rect 75276 238824 75328 238876
rect 240140 238756 240192 238808
rect 241244 238756 241296 238808
rect 257436 238756 257488 238808
rect 96620 238688 96672 238740
rect 214196 238688 214248 238740
rect 218152 238688 218204 238740
rect 240324 238688 240376 238740
rect 241796 238688 241848 238740
rect 258172 238688 258224 238740
rect 107660 238620 107712 238672
rect 219900 238620 219952 238672
rect 221096 238620 221148 238672
rect 227628 238620 227680 238672
rect 238760 238620 238812 238672
rect 243912 238620 243964 238672
rect 231124 238552 231176 238604
rect 234712 238552 234764 238604
rect 229100 238076 229152 238128
rect 230480 238076 230532 238128
rect 61752 238008 61804 238060
rect 108304 238008 108356 238060
rect 241796 237804 241848 237856
rect 242440 237804 242492 237856
rect 65892 237532 65944 237584
rect 72516 237532 72568 237584
rect 214196 237464 214248 237516
rect 214656 237464 214708 237516
rect 214564 237396 214616 237448
rect 216036 237396 216088 237448
rect 240324 237396 240376 237448
rect 240784 237396 240836 237448
rect 115940 237328 115992 237380
rect 224316 237328 224368 237380
rect 231768 237328 231820 237380
rect 247224 237328 247276 237380
rect 54852 237260 54904 237312
rect 120724 237260 120776 237312
rect 136088 237260 136140 237312
rect 149704 237260 149756 237312
rect 151912 237260 151964 237312
rect 170588 237260 170640 237312
rect 169760 236648 169812 236700
rect 202788 236648 202840 236700
rect 204168 236648 204220 236700
rect 214748 236648 214800 236700
rect 224316 236648 224368 236700
rect 303804 236648 303856 236700
rect 225696 236036 225748 236088
rect 229652 236036 229704 236088
rect 65984 235900 66036 235952
rect 167644 235900 167696 235952
rect 48136 235832 48188 235884
rect 118884 235832 118936 235884
rect 138020 235832 138072 235884
rect 155408 235832 155460 235884
rect 155684 235764 155736 235816
rect 159548 235764 159600 235816
rect 199936 235288 199988 235340
rect 204996 235288 205048 235340
rect 124128 235220 124180 235272
rect 135352 235220 135404 235272
rect 173440 235220 173492 235272
rect 198832 235220 198884 235272
rect 205088 235220 205140 235272
rect 582748 235220 582800 235272
rect 118884 234608 118936 234660
rect 119344 234608 119396 234660
rect 200304 234608 200356 234660
rect 202144 234608 202196 234660
rect 225604 234608 225656 234660
rect 226156 234608 226208 234660
rect 292580 234608 292632 234660
rect 60372 234540 60424 234592
rect 153844 234540 153896 234592
rect 188436 234540 188488 234592
rect 240140 234540 240192 234592
rect 123024 234472 123076 234524
rect 181628 234472 181680 234524
rect 209136 233248 209188 233300
rect 221004 233248 221056 233300
rect 222108 233248 222160 233300
rect 233976 233248 234028 233300
rect 295524 233248 295576 233300
rect 126980 233180 127032 233232
rect 230480 233180 230532 233232
rect 231768 233180 231820 233232
rect 108304 233112 108356 233164
rect 156788 233112 156840 233164
rect 180064 233112 180116 233164
rect 203616 233112 203668 233164
rect 204076 233112 204128 233164
rect 218980 233112 219032 233164
rect 220360 233112 220412 233164
rect 53472 232500 53524 232552
rect 106740 232500 106792 232552
rect 102140 231820 102192 231872
rect 104164 231820 104216 231872
rect 219532 231820 219584 231872
rect 220360 231820 220412 231872
rect 292672 231820 292724 231872
rect 124864 231752 124916 231804
rect 189908 231752 189960 231804
rect 190000 231752 190052 231804
rect 243636 231752 243688 231804
rect 114376 231684 114428 231736
rect 133512 231684 133564 231736
rect 147588 231684 147640 231736
rect 159456 231684 159508 231736
rect 48044 231616 48096 231668
rect 125324 231616 125376 231668
rect 217140 231480 217192 231532
rect 221464 231480 221516 231532
rect 198740 231072 198792 231124
rect 217324 231072 217376 231124
rect 231768 231072 231820 231124
rect 311992 231072 312044 231124
rect 133604 230460 133656 230512
rect 146116 230460 146168 230512
rect 142068 230392 142120 230444
rect 233976 230392 234028 230444
rect 144828 230324 144880 230376
rect 148324 230324 148376 230376
rect 166908 230324 166960 230376
rect 167736 230324 167788 230376
rect 198832 230324 198884 230376
rect 222844 230324 222896 230376
rect 85580 229712 85632 229764
rect 144184 229712 144236 229764
rect 148876 229712 148928 229764
rect 166908 229712 166960 229764
rect 181536 229712 181588 229764
rect 195612 229712 195664 229764
rect 146116 229032 146168 229084
rect 156880 229032 156932 229084
rect 180340 229032 180392 229084
rect 220452 229032 220504 229084
rect 227260 228420 227312 228472
rect 309232 228420 309284 228472
rect 63316 228352 63368 228404
rect 106924 228352 106976 228404
rect 125416 228352 125468 228404
rect 190828 228352 190880 228404
rect 195796 228352 195848 228404
rect 299756 228352 299808 228404
rect 220268 227808 220320 227860
rect 227260 227808 227312 227860
rect 220084 227740 220136 227792
rect 220452 227740 220504 227792
rect 151084 227672 151136 227724
rect 249984 227672 250036 227724
rect 66076 227604 66128 227656
rect 155316 227604 155368 227656
rect 63224 226992 63276 227044
rect 134524 226992 134576 227044
rect 214748 226992 214800 227044
rect 272524 226992 272576 227044
rect 276664 226992 276716 227044
rect 305092 226992 305144 227044
rect 160744 226312 160796 226364
rect 116584 226244 116636 226296
rect 185676 226244 185728 226296
rect 188620 226244 188672 226296
rect 206836 226244 206888 226296
rect 240692 226244 240744 226296
rect 151084 225564 151136 225616
rect 162400 225564 162452 225616
rect 201408 225292 201460 225344
rect 203616 225292 203668 225344
rect 206284 225156 206336 225208
rect 206836 225156 206888 225208
rect 203524 224952 203576 225004
rect 214748 224952 214800 225004
rect 240968 224952 241020 225004
rect 243268 224952 243320 225004
rect 70400 224884 70452 224936
rect 215944 224884 215996 224936
rect 110236 224816 110288 224868
rect 178868 224816 178920 224868
rect 195612 224816 195664 224868
rect 224316 224816 224368 224868
rect 224868 224816 224920 224868
rect 229008 224204 229060 224256
rect 307852 224204 307904 224256
rect 82728 223524 82780 223576
rect 248512 223524 248564 223576
rect 155224 222844 155276 222896
rect 195244 222844 195296 222896
rect 201592 222844 201644 222896
rect 226984 222844 227036 222896
rect 72516 222096 72568 222148
rect 159364 222096 159416 222148
rect 174728 222096 174780 222148
rect 247040 222096 247092 222148
rect 133880 221416 133932 221468
rect 191840 221416 191892 221468
rect 202144 221416 202196 221468
rect 294144 221416 294196 221468
rect 580908 221144 580960 221196
rect 583576 221144 583628 221196
rect 4804 220804 4856 220856
rect 93768 220804 93820 220856
rect 148324 220736 148376 220788
rect 236920 220736 236972 220788
rect 107476 220668 107528 220720
rect 158076 220668 158128 220720
rect 166356 220668 166408 220720
rect 223764 220668 223816 220720
rect 236920 220056 236972 220108
rect 306656 220056 306708 220108
rect 223764 219920 223816 219972
rect 224224 219920 224276 219972
rect 130936 219376 130988 219428
rect 186964 219376 187016 219428
rect 565084 219376 565136 219428
rect 580172 219376 580224 219428
rect 171968 219308 172020 219360
rect 223396 219308 223448 219360
rect 81256 218764 81308 218816
rect 128360 218764 128412 218816
rect 21364 218696 21416 218748
rect 156604 218696 156656 218748
rect 224408 218696 224460 218748
rect 238852 218696 238904 218748
rect 222936 218084 222988 218136
rect 223396 218084 223448 218136
rect 186964 218016 187016 218068
rect 187148 218016 187200 218068
rect 104808 217268 104860 217320
rect 172796 217268 172848 217320
rect 187516 217268 187568 217320
rect 198004 217268 198056 217320
rect 206284 217268 206336 217320
rect 236644 217268 236696 217320
rect 236736 217268 236788 217320
rect 254032 217268 254084 217320
rect 254584 217268 254636 217320
rect 317420 217268 317472 217320
rect 142804 216656 142856 216708
rect 234620 216656 234672 216708
rect 131028 216588 131080 216640
rect 191196 216588 191248 216640
rect 191840 216588 191892 216640
rect 241520 216588 241572 216640
rect 242256 216588 242308 216640
rect 111800 215908 111852 215960
rect 191656 215908 191708 215960
rect 200028 215908 200080 215960
rect 230480 215908 230532 215960
rect 67732 215228 67784 215280
rect 206468 215228 206520 215280
rect 73896 215160 73948 215212
rect 151084 215160 151136 215212
rect 205088 214616 205140 214668
rect 245660 214616 245712 214668
rect 238116 214548 238168 214600
rect 309324 214548 309376 214600
rect 233240 214344 233292 214396
rect 234436 214344 234488 214396
rect 213000 213936 213052 213988
rect 233240 213936 233292 213988
rect 64696 213868 64748 213920
rect 191932 213868 191984 213920
rect 191656 213800 191708 213852
rect 222292 213800 222344 213852
rect 223028 213800 223080 213852
rect 197360 213256 197412 213308
rect 214840 213256 214892 213308
rect 134524 213188 134576 213240
rect 186964 213188 187016 213240
rect 214656 213188 214708 213240
rect 302516 213188 302568 213240
rect 249064 212780 249116 212832
rect 251272 212780 251324 212832
rect 122840 212440 122892 212492
rect 227812 212440 227864 212492
rect 228364 212440 228416 212492
rect 77392 212372 77444 212424
rect 147680 212372 147732 212424
rect 195244 212372 195296 212424
rect 245752 212372 245804 212424
rect 148968 211760 149020 211812
rect 171784 211760 171836 211812
rect 172428 211148 172480 211200
rect 192484 211148 192536 211200
rect 237380 211148 237432 211200
rect 238300 211148 238352 211200
rect 246304 211148 246356 211200
rect 76656 211080 76708 211132
rect 213000 211080 213052 211132
rect 104900 211012 104952 211064
rect 188528 211012 188580 211064
rect 214840 210468 214892 210520
rect 251272 210468 251324 210520
rect 214748 210400 214800 210452
rect 302424 210400 302476 210452
rect 132408 209720 132460 209772
rect 244464 209720 244516 209772
rect 75276 209652 75328 209704
rect 142804 209652 142856 209704
rect 144184 209040 144236 209092
rect 213736 209040 213788 209092
rect 213736 208360 213788 208412
rect 238116 208360 238168 208412
rect 113088 208292 113140 208344
rect 247132 208292 247184 208344
rect 69020 207612 69072 207664
rect 200028 207612 200080 207664
rect 57704 206932 57756 206984
rect 209044 206932 209096 206984
rect 99472 206864 99524 206916
rect 211804 206864 211856 206916
rect 212448 206864 212500 206916
rect 212448 206320 212500 206372
rect 231124 206320 231176 206372
rect 220176 206252 220228 206304
rect 295616 206252 295668 206304
rect 95240 205572 95292 205624
rect 244280 205572 244332 205624
rect 195336 204960 195388 205012
rect 218888 204960 218940 205012
rect 83464 204892 83516 204944
rect 167000 204892 167052 204944
rect 218796 204892 218848 204944
rect 283012 204892 283064 204944
rect 137928 204212 137980 204264
rect 232136 204212 232188 204264
rect 233148 204212 233200 204264
rect 191196 203668 191248 203720
rect 231952 203668 232004 203720
rect 146208 203532 146260 203584
rect 191288 203532 191340 203584
rect 233148 203532 233200 203584
rect 303712 203532 303764 203584
rect 3056 202784 3108 202836
rect 124128 202784 124180 202836
rect 125508 202784 125560 202836
rect 251456 202784 251508 202836
rect 167000 202716 167052 202768
rect 202880 202716 202932 202768
rect 203524 202716 203576 202768
rect 83096 202104 83148 202156
rect 166816 202104 166868 202156
rect 200028 201424 200080 201476
rect 282184 201492 282236 201544
rect 76564 201356 76616 201408
rect 200856 201356 200908 201408
rect 225696 200812 225748 200864
rect 291292 200812 291344 200864
rect 86868 200744 86920 200796
rect 189724 200744 189776 200796
rect 204996 200744 205048 200796
rect 285772 200744 285824 200796
rect 93124 200064 93176 200116
rect 198740 200064 198792 200116
rect 223028 199452 223080 199504
rect 279056 199452 279108 199504
rect 118608 199384 118660 199436
rect 202144 199384 202196 199436
rect 211896 199384 211948 199436
rect 305184 199384 305236 199436
rect 50804 198636 50856 198688
rect 180248 198636 180300 198688
rect 191288 198636 191340 198688
rect 97816 198568 97868 198620
rect 158720 198568 158772 198620
rect 166816 198568 166868 198620
rect 207664 198568 207716 198620
rect 244280 198500 244332 198552
rect 244924 198500 244976 198552
rect 46848 197276 46900 197328
rect 173256 197276 173308 197328
rect 143448 197208 143500 197260
rect 163504 197208 163556 197260
rect 174636 196596 174688 196648
rect 212080 196596 212132 196648
rect 213828 196596 213880 196648
rect 226984 196596 227036 196648
rect 223028 195984 223080 196036
rect 249892 195984 249944 196036
rect 79876 195916 79928 195968
rect 226340 195916 226392 195968
rect 106924 195848 106976 195900
rect 214564 195848 214616 195900
rect 218888 195236 218940 195288
rect 237472 195236 237524 195288
rect 63132 194488 63184 194540
rect 210424 194488 210476 194540
rect 212080 193876 212132 193928
rect 232504 193876 232556 193928
rect 81348 193808 81400 193860
rect 176016 193808 176068 193860
rect 199384 193808 199436 193860
rect 230572 193808 230624 193860
rect 238024 193808 238076 193860
rect 281724 193808 281776 193860
rect 166908 192516 166960 192568
rect 237380 192516 237432 192568
rect 72424 192448 72476 192500
rect 171968 192448 172020 192500
rect 207664 192448 207716 192500
rect 287336 192448 287388 192500
rect 73160 191768 73212 191820
rect 202604 191768 202656 191820
rect 206376 191156 206428 191208
rect 301044 191156 301096 191208
rect 192576 191088 192628 191140
rect 292764 191088 292816 191140
rect 133788 190476 133840 190528
rect 192668 190476 192720 190528
rect 89536 189728 89588 189780
rect 191196 189728 191248 189780
rect 194508 189728 194560 189780
rect 220728 189728 220780 189780
rect 267004 189728 267056 189780
rect 307944 189728 307996 189780
rect 113088 189048 113140 189100
rect 170588 189116 170640 189168
rect 221464 189116 221516 189168
rect 234712 189116 234764 189168
rect 169760 189048 169812 189100
rect 335360 189048 335412 189100
rect 3516 188980 3568 189032
rect 35164 188980 35216 189032
rect 89628 188980 89680 189032
rect 223028 188980 223080 189032
rect 240784 188368 240836 188420
rect 279148 188368 279200 188420
rect 191748 188300 191800 188352
rect 214564 188300 214616 188352
rect 224316 188300 224368 188352
rect 236092 188300 236144 188352
rect 236736 188300 236788 188352
rect 283196 188300 283248 188352
rect 304264 188300 304316 188352
rect 325700 188300 325752 188352
rect 131028 187688 131080 187740
rect 188620 187688 188672 187740
rect 52276 187620 52328 187672
rect 221464 187620 221516 187672
rect 280804 187620 280856 187672
rect 288624 187620 288676 187672
rect 180708 186940 180760 186992
rect 237564 186940 237616 186992
rect 128268 186328 128320 186380
rect 174636 186328 174688 186380
rect 222108 186328 222160 186380
rect 293960 186328 294012 186380
rect 188528 185648 188580 185700
rect 231216 185648 231268 185700
rect 220268 185580 220320 185632
rect 280160 185580 280212 185632
rect 106188 184968 106240 185020
rect 182916 184968 182968 185020
rect 121368 184900 121420 184952
rect 207664 184900 207716 184952
rect 200764 184220 200816 184272
rect 236000 184220 236052 184272
rect 184848 184152 184900 184204
rect 303896 184152 303948 184204
rect 243820 183744 243872 183796
rect 245752 183744 245804 183796
rect 100668 183608 100720 183660
rect 180248 183608 180300 183660
rect 108948 183540 109000 183592
rect 195336 183540 195388 183592
rect 203616 182860 203668 182912
rect 238760 182860 238812 182912
rect 271328 182860 271380 182912
rect 281816 182860 281868 182912
rect 178868 182792 178920 182844
rect 284484 182792 284536 182844
rect 132408 182248 132460 182300
rect 172060 182248 172112 182300
rect 102048 182180 102100 182232
rect 167736 182180 167788 182232
rect 209136 181500 209188 181552
rect 233332 181500 233384 181552
rect 236000 181500 236052 181552
rect 274548 181500 274600 181552
rect 167644 181432 167696 181484
rect 245752 181432 245804 181484
rect 269856 181432 269908 181484
rect 298376 181432 298428 181484
rect 125968 180888 126020 180940
rect 166448 180888 166500 180940
rect 148232 180820 148284 180872
rect 209044 180820 209096 180872
rect 232504 180208 232556 180260
rect 241704 180208 241756 180260
rect 214564 180140 214616 180192
rect 233148 180140 233200 180192
rect 272524 180140 272576 180192
rect 292856 180140 292908 180192
rect 169024 180072 169076 180124
rect 224224 180072 224276 180124
rect 239404 180072 239456 180124
rect 252652 180072 252704 180124
rect 257436 180072 257488 180124
rect 288532 180072 288584 180124
rect 192484 179868 192536 179920
rect 198004 179868 198056 179920
rect 129464 179460 129516 179512
rect 165436 179460 165488 179512
rect 121920 179392 121972 179444
rect 192576 179392 192628 179444
rect 224316 179392 224368 179444
rect 229468 179392 229520 179444
rect 574744 179324 574796 179376
rect 580172 179324 580224 179376
rect 224224 179256 224276 179308
rect 229928 179256 229980 179308
rect 171968 178712 172020 178764
rect 197360 178712 197412 178764
rect 278044 178712 278096 178764
rect 294236 178712 294288 178764
rect 184296 178644 184348 178696
rect 242900 178644 242952 178696
rect 243544 178644 243596 178696
rect 287152 178644 287204 178696
rect 123300 178100 123352 178152
rect 164976 178100 165028 178152
rect 115848 178032 115900 178084
rect 171876 178032 171928 178084
rect 222844 177352 222896 177404
rect 232136 177352 232188 177404
rect 271144 177352 271196 177404
rect 285864 177352 285916 177404
rect 193864 177284 193916 177336
rect 229376 177284 229428 177336
rect 231216 177284 231268 177336
rect 238852 177284 238904 177336
rect 268384 177284 268436 177336
rect 287244 177284 287296 177336
rect 128176 176808 128228 176860
rect 207020 176808 207072 176860
rect 158996 176740 159048 176792
rect 174728 176740 174780 176792
rect 67548 176672 67600 176724
rect 70492 176672 70544 176724
rect 136088 176672 136140 176724
rect 213920 176604 213972 176656
rect 164884 176196 164936 176248
rect 167000 176196 167052 176248
rect 231124 176128 231176 176180
rect 236000 176128 236052 176180
rect 220084 175992 220136 176044
rect 231860 175992 231912 176044
rect 233148 175992 233200 176044
rect 244372 175992 244424 176044
rect 276664 175992 276716 176044
rect 284576 175992 284628 176044
rect 119436 175924 119488 175976
rect 165068 175924 165120 175976
rect 207020 175924 207072 175976
rect 214104 175924 214156 175976
rect 215208 175924 215260 175976
rect 229192 175924 229244 175976
rect 246304 175924 246356 175976
rect 278780 175924 278832 175976
rect 224960 175788 225012 175840
rect 273352 175788 273404 175840
rect 135260 175176 135312 175228
rect 213920 175176 213972 175228
rect 243636 175244 243688 175296
rect 264980 175244 265032 175296
rect 229284 175176 229336 175228
rect 229928 175176 229980 175228
rect 230848 175176 230900 175228
rect 231124 175176 231176 175228
rect 249892 175176 249944 175228
rect 279424 175176 279476 175228
rect 192668 175108 192720 175160
rect 214012 175108 214064 175160
rect 263140 173952 263192 174004
rect 264980 173952 265032 174004
rect 214564 173884 214616 173936
rect 242992 173884 243044 173936
rect 245016 173884 245068 173936
rect 265072 173884 265124 173936
rect 172060 173816 172112 173868
rect 213920 173816 213972 173868
rect 231584 173816 231636 173868
rect 239404 173816 239456 173868
rect 282460 173816 282512 173868
rect 289912 173816 289964 173868
rect 188620 173748 188672 173800
rect 214012 173748 214064 173800
rect 229100 173612 229152 173664
rect 229468 173612 229520 173664
rect 250536 172592 250588 172644
rect 264980 172592 265032 172644
rect 238208 172524 238260 172576
rect 265072 172524 265124 172576
rect 165436 172456 165488 172508
rect 213920 172456 213972 172508
rect 231584 172456 231636 172508
rect 240232 172456 240284 172508
rect 282092 172456 282144 172508
rect 295616 172456 295668 172508
rect 240232 171776 240284 171828
rect 248420 171776 248472 171828
rect 258816 171232 258868 171284
rect 264980 171232 265032 171284
rect 240784 171096 240836 171148
rect 265072 171096 265124 171148
rect 166448 171028 166500 171080
rect 214012 171028 214064 171080
rect 231124 171028 231176 171080
rect 233516 171028 233568 171080
rect 282828 171028 282880 171080
rect 298192 171028 298244 171080
rect 174636 170960 174688 171012
rect 213920 170960 213972 171012
rect 236828 169804 236880 169856
rect 264980 169804 265032 169856
rect 233976 169736 234028 169788
rect 265072 169736 265124 169788
rect 164976 169668 165028 169720
rect 214012 169668 214064 169720
rect 167828 169600 167880 169652
rect 213920 169600 213972 169652
rect 281540 169464 281592 169516
rect 283196 169464 283248 169516
rect 282828 169396 282880 169448
rect 287336 169396 287388 169448
rect 238392 169056 238444 169108
rect 241612 169056 241664 169108
rect 231676 168988 231728 169040
rect 247040 168988 247092 169040
rect 247776 168444 247828 168496
rect 264980 168444 265032 168496
rect 242256 168376 242308 168428
rect 265072 168376 265124 168428
rect 192576 168308 192628 168360
rect 213920 168308 213972 168360
rect 231768 168308 231820 168360
rect 240232 168308 240284 168360
rect 282828 167696 282880 167748
rect 288716 167696 288768 167748
rect 174728 167628 174780 167680
rect 214564 167628 214616 167680
rect 229744 167628 229796 167680
rect 239036 167628 239088 167680
rect 248052 167084 248104 167136
rect 264980 167084 265032 167136
rect 239496 167016 239548 167068
rect 265072 167016 265124 167068
rect 280068 167016 280120 167068
rect 280436 167016 280488 167068
rect 165068 166948 165120 167000
rect 213920 166948 213972 167000
rect 282828 166948 282880 167000
rect 291384 166948 291436 167000
rect 170496 166880 170548 166932
rect 214012 166880 214064 166932
rect 231768 166676 231820 166728
rect 234896 166676 234948 166728
rect 230480 166268 230532 166320
rect 230848 166268 230900 166320
rect 236092 166268 236144 166320
rect 258080 166268 258132 166320
rect 262864 165656 262916 165708
rect 265348 165656 265400 165708
rect 232780 165588 232832 165640
rect 264980 165588 265032 165640
rect 166540 165520 166592 165572
rect 214012 165520 214064 165572
rect 231492 165520 231544 165572
rect 244372 165520 244424 165572
rect 282000 165520 282052 165572
rect 284576 165520 284628 165572
rect 171876 165452 171928 165504
rect 213920 165452 213972 165504
rect 231124 164840 231176 164892
rect 248512 164840 248564 164892
rect 257620 164296 257672 164348
rect 265072 164296 265124 164348
rect 251824 164228 251876 164280
rect 264980 164228 265032 164280
rect 3240 164160 3292 164212
rect 25504 164160 25556 164212
rect 169208 164160 169260 164212
rect 213920 164160 213972 164212
rect 282828 164160 282880 164212
rect 303804 164160 303856 164212
rect 170588 164092 170640 164144
rect 214012 164092 214064 164144
rect 282460 164092 282512 164144
rect 285956 164092 286008 164144
rect 231768 163956 231820 164008
rect 236092 163956 236144 164008
rect 250628 162936 250680 162988
rect 264980 162936 265032 162988
rect 235540 162868 235592 162920
rect 265072 162868 265124 162920
rect 173256 162800 173308 162852
rect 214012 162800 214064 162852
rect 282828 162800 282880 162852
rect 292764 162800 292816 162852
rect 177396 162732 177448 162784
rect 213920 162732 213972 162784
rect 231308 162528 231360 162580
rect 237564 162528 237616 162580
rect 236736 162120 236788 162172
rect 265164 162120 265216 162172
rect 254584 161440 254636 161492
rect 264980 161440 265032 161492
rect 169024 161372 169076 161424
rect 214012 161372 214064 161424
rect 231768 161372 231820 161424
rect 242992 161372 243044 161424
rect 195336 161304 195388 161356
rect 213920 161304 213972 161356
rect 230940 160964 230992 161016
rect 233240 160964 233292 161016
rect 245292 160692 245344 160744
rect 262864 160692 262916 160744
rect 281540 160216 281592 160268
rect 281816 160216 281868 160268
rect 282828 160148 282880 160200
rect 288624 160148 288676 160200
rect 238024 160080 238076 160132
rect 264980 160080 265032 160132
rect 182916 160012 182968 160064
rect 213920 160012 213972 160064
rect 231768 160012 231820 160064
rect 241704 160012 241756 160064
rect 281908 160012 281960 160064
rect 294236 160012 294288 160064
rect 198096 159944 198148 159996
rect 214012 159944 214064 159996
rect 282368 159944 282420 159996
rect 290096 159944 290148 159996
rect 243912 158788 243964 158840
rect 265072 158788 265124 158840
rect 233884 158720 233936 158772
rect 264980 158720 265032 158772
rect 167736 158652 167788 158704
rect 214012 158652 214064 158704
rect 282092 158652 282144 158704
rect 300952 158652 301004 158704
rect 181536 158584 181588 158636
rect 213920 158584 213972 158636
rect 231216 158584 231268 158636
rect 240140 158584 240192 158636
rect 241152 157428 241204 157480
rect 265072 157428 265124 157480
rect 235264 157360 235316 157412
rect 264980 157360 265032 157412
rect 166356 157292 166408 157344
rect 213920 157292 213972 157344
rect 180248 157224 180300 157276
rect 214012 157224 214064 157276
rect 230940 156952 230992 157004
rect 233424 156952 233476 157004
rect 236644 156612 236696 156664
rect 265256 156612 265308 156664
rect 242440 155932 242492 155984
rect 264980 155932 265032 155984
rect 178960 155864 179012 155916
rect 213920 155864 213972 155916
rect 230848 155864 230900 155916
rect 236000 155864 236052 155916
rect 282276 155864 282328 155916
rect 310612 155864 310664 155916
rect 185768 155796 185820 155848
rect 214012 155796 214064 155848
rect 246580 154640 246632 154692
rect 265072 154640 265124 154692
rect 241060 154572 241112 154624
rect 264980 154572 265032 154624
rect 282276 154504 282328 154556
rect 302516 154504 302568 154556
rect 282828 154436 282880 154488
rect 292856 154436 292908 154488
rect 231308 154368 231360 154420
rect 237380 154368 237432 154420
rect 234160 153824 234212 153876
rect 265716 153824 265768 153876
rect 192576 153280 192628 153332
rect 213920 153280 213972 153332
rect 185676 153212 185728 153264
rect 214012 153212 214064 153264
rect 262956 153212 263008 153264
rect 265348 153212 265400 153264
rect 230480 153144 230532 153196
rect 234620 153144 234672 153196
rect 167644 152464 167696 152516
rect 194508 152464 194560 152516
rect 242164 151852 242216 151904
rect 264980 151852 265032 151904
rect 206284 151784 206336 151836
rect 213920 151784 213972 151836
rect 238116 151784 238168 151836
rect 265072 151784 265124 151836
rect 281908 151716 281960 151768
rect 307852 151716 307904 151768
rect 231584 151104 231636 151156
rect 251272 151104 251324 151156
rect 232872 151036 232924 151088
rect 265624 151036 265676 151088
rect 206376 150492 206428 150544
rect 213920 150492 213972 150544
rect 183008 150424 183060 150476
rect 214104 150424 214156 150476
rect 261484 150424 261536 150476
rect 264980 150424 265032 150476
rect 194508 150356 194560 150408
rect 214012 150356 214064 150408
rect 230572 150356 230624 150408
rect 241520 150356 241572 150408
rect 2780 150288 2832 150340
rect 4804 150288 4856 150340
rect 209044 150288 209096 150340
rect 213920 150288 213972 150340
rect 249248 149676 249300 149728
rect 265164 149676 265216 149728
rect 256056 149064 256108 149116
rect 264980 149064 265032 149116
rect 231768 148996 231820 149048
rect 247224 148996 247276 149048
rect 282828 148996 282880 149048
rect 306564 148996 306616 149048
rect 234068 148316 234120 148368
rect 265256 148316 265308 148368
rect 282644 147840 282696 147892
rect 287244 147840 287296 147892
rect 166356 147636 166408 147688
rect 213920 147636 213972 147688
rect 259092 147636 259144 147688
rect 264980 147636 265032 147688
rect 282828 147568 282880 147620
rect 305184 147568 305236 147620
rect 282276 147500 282328 147552
rect 298284 147500 298336 147552
rect 239680 146888 239732 146940
rect 265072 146888 265124 146940
rect 231124 146820 231176 146872
rect 236828 146820 236880 146872
rect 231308 146548 231360 146600
rect 238208 146548 238260 146600
rect 184388 146276 184440 146328
rect 213920 146276 213972 146328
rect 247960 146276 248012 146328
rect 264980 146276 265032 146328
rect 282828 146208 282880 146260
rect 313280 146208 313332 146260
rect 282736 146140 282788 146192
rect 294144 146140 294196 146192
rect 231216 145528 231268 145580
rect 240784 145528 240836 145580
rect 198188 144984 198240 145036
rect 214012 144984 214064 145036
rect 240968 144984 241020 145036
rect 264980 144984 265032 145036
rect 169024 144916 169076 144968
rect 213920 144916 213972 144968
rect 235356 144916 235408 144968
rect 265072 144916 265124 144968
rect 282828 144848 282880 144900
rect 299756 144848 299808 144900
rect 173164 144168 173216 144220
rect 184296 144168 184348 144220
rect 230572 144168 230624 144220
rect 249064 144168 249116 144220
rect 231768 144032 231820 144084
rect 238392 144032 238444 144084
rect 202236 143624 202288 143676
rect 214012 143624 214064 143676
rect 250812 143624 250864 143676
rect 265072 143624 265124 143676
rect 189816 143556 189868 143608
rect 213920 143556 213972 143608
rect 242348 143556 242400 143608
rect 264980 143556 265032 143608
rect 231768 143488 231820 143540
rect 243820 143488 243872 143540
rect 282828 143488 282880 143540
rect 295340 143488 295392 143540
rect 171784 142808 171836 142860
rect 193864 142808 193916 142860
rect 209228 142196 209280 142248
rect 213920 142196 213972 142248
rect 254768 142196 254820 142248
rect 265072 142196 265124 142248
rect 180340 142128 180392 142180
rect 214012 142128 214064 142180
rect 238208 142128 238260 142180
rect 264980 142128 265032 142180
rect 282552 142060 282604 142112
rect 285864 142060 285916 142112
rect 169116 141380 169168 141432
rect 209044 141380 209096 141432
rect 230940 141380 230992 141432
rect 263140 141380 263192 141432
rect 282828 141312 282880 141364
rect 288440 141312 288492 141364
rect 263048 140836 263100 140888
rect 265256 140836 265308 140888
rect 180248 140768 180300 140820
rect 213920 140768 213972 140820
rect 236828 140768 236880 140820
rect 264980 140768 265032 140820
rect 231768 140700 231820 140752
rect 245752 140700 245804 140752
rect 282828 140700 282880 140752
rect 291476 140700 291528 140752
rect 180156 140020 180208 140072
rect 199384 140020 199436 140072
rect 240784 140020 240836 140072
rect 263232 140020 263284 140072
rect 210608 139476 210660 139528
rect 214104 139476 214156 139528
rect 259000 139476 259052 139528
rect 265164 139476 265216 139528
rect 211804 139408 211856 139460
rect 213920 139408 213972 139460
rect 263140 139408 263192 139460
rect 264980 139408 265032 139460
rect 177304 138660 177356 138712
rect 200856 138660 200908 138712
rect 229928 138660 229980 138712
rect 264980 138660 265032 138712
rect 281540 138320 281592 138372
rect 284484 138320 284536 138372
rect 192484 137980 192536 138032
rect 213920 137980 213972 138032
rect 231492 137912 231544 137964
rect 254032 137912 254084 137964
rect 231768 137844 231820 137896
rect 242900 137844 242952 137896
rect 282828 137436 282880 137488
rect 287060 137436 287112 137488
rect 181536 137232 181588 137284
rect 214012 137232 214064 137284
rect 3516 136892 3568 136944
rect 7564 136892 7616 136944
rect 257528 136688 257580 136740
rect 264980 136688 265032 136740
rect 171784 136620 171836 136672
rect 213920 136620 213972 136672
rect 243728 136620 243780 136672
rect 265072 136620 265124 136672
rect 231768 136552 231820 136604
rect 256700 136552 256752 136604
rect 282828 136552 282880 136604
rect 296904 136552 296956 136604
rect 231676 136484 231728 136536
rect 245016 136484 245068 136536
rect 170404 135872 170456 135924
rect 209136 135872 209188 135924
rect 187056 135260 187108 135312
rect 213920 135260 213972 135312
rect 256240 135260 256292 135312
rect 264980 135260 265032 135312
rect 231768 135192 231820 135244
rect 256148 135192 256200 135244
rect 231676 135124 231728 135176
rect 249156 135124 249208 135176
rect 166264 134580 166316 134632
rect 185584 134580 185636 134632
rect 178868 134512 178920 134564
rect 214012 134512 214064 134564
rect 261760 133968 261812 134020
rect 265072 133968 265124 134020
rect 204996 133900 205048 133952
rect 213920 133900 213972 133952
rect 257436 133900 257488 133952
rect 264980 133900 265032 133952
rect 231492 133832 231544 133884
rect 250536 133832 250588 133884
rect 282828 133832 282880 133884
rect 309324 133832 309376 133884
rect 230756 133152 230808 133204
rect 239496 133152 239548 133204
rect 202420 132540 202472 132592
rect 213920 132540 213972 132592
rect 173164 132472 173216 132524
rect 214012 132472 214064 132524
rect 230940 132404 230992 132456
rect 244924 132404 244976 132456
rect 282828 132404 282880 132456
rect 311900 132404 311952 132456
rect 181444 131724 181496 131776
rect 209228 131724 209280 131776
rect 264244 131588 264296 131640
rect 267188 131588 267240 131640
rect 230480 131316 230532 131368
rect 233976 131316 234028 131368
rect 209320 131180 209372 131232
rect 213920 131180 213972 131232
rect 205088 131112 205140 131164
rect 214012 131112 214064 131164
rect 245200 131112 245252 131164
rect 264980 131112 265032 131164
rect 231768 131044 231820 131096
rect 260288 131044 260340 131096
rect 231492 130976 231544 131028
rect 242256 130976 242308 131028
rect 282276 130976 282328 131028
rect 285680 130976 285732 131028
rect 207664 129820 207716 129872
rect 213920 129820 213972 129872
rect 164884 129752 164936 129804
rect 214012 129752 214064 129804
rect 253388 129752 253440 129804
rect 264980 129752 265032 129804
rect 231768 129684 231820 129736
rect 247776 129684 247828 129736
rect 282092 129684 282144 129736
rect 301044 129684 301096 129736
rect 231492 129548 231544 129600
rect 236736 129548 236788 129600
rect 167828 129004 167880 129056
rect 206376 129004 206428 129056
rect 210424 128392 210476 128444
rect 214012 128392 214064 128444
rect 261576 128392 261628 128444
rect 265164 128392 265216 128444
rect 196808 128324 196860 128376
rect 213920 128324 213972 128376
rect 244924 128324 244976 128376
rect 264980 128324 265032 128376
rect 231768 128256 231820 128308
rect 253296 128256 253348 128308
rect 282000 128256 282052 128308
rect 311992 128256 312044 128308
rect 231676 128188 231728 128240
rect 248052 128188 248104 128240
rect 282828 128188 282880 128240
rect 306656 128188 306708 128240
rect 174636 127576 174688 127628
rect 211804 127576 211856 127628
rect 247868 127576 247920 127628
rect 265072 127576 265124 127628
rect 59176 126964 59228 127016
rect 65524 126964 65576 127016
rect 195336 126964 195388 127016
rect 213920 126964 213972 127016
rect 231768 126896 231820 126948
rect 245292 126896 245344 126948
rect 282276 126896 282328 126948
rect 296720 126896 296772 126948
rect 173256 126216 173308 126268
rect 214564 126216 214616 126268
rect 231124 126216 231176 126268
rect 246580 126216 246632 126268
rect 253296 125672 253348 125724
rect 265072 125672 265124 125724
rect 206376 125604 206428 125656
rect 213920 125604 213972 125656
rect 249156 125604 249208 125656
rect 264980 125604 265032 125656
rect 282828 125536 282880 125588
rect 317420 125536 317472 125588
rect 282736 125468 282788 125520
rect 314660 125468 314712 125520
rect 230848 124924 230900 124976
rect 242440 124924 242492 124976
rect 171876 124856 171928 124908
rect 206284 124856 206336 124908
rect 230940 124856 230992 124908
rect 250628 124856 250680 124908
rect 252008 124244 252060 124296
rect 265072 124244 265124 124296
rect 191104 124176 191156 124228
rect 213920 124176 213972 124228
rect 243544 124176 243596 124228
rect 264980 124176 265032 124228
rect 282276 124108 282328 124160
rect 296812 124108 296864 124160
rect 282828 124040 282880 124092
rect 294052 124040 294104 124092
rect 231768 123836 231820 123888
rect 235540 123836 235592 123888
rect 230664 123428 230716 123480
rect 243912 123428 243964 123480
rect 250720 123428 250772 123480
rect 263140 123428 263192 123480
rect 187148 122884 187200 122936
rect 214012 122884 214064 122936
rect 166264 122816 166316 122868
rect 213920 122816 213972 122868
rect 240876 122816 240928 122868
rect 264980 122816 265032 122868
rect 282828 122748 282880 122800
rect 307944 122748 307996 122800
rect 231584 122680 231636 122732
rect 254584 122680 254636 122732
rect 230756 122476 230808 122528
rect 232596 122476 232648 122528
rect 169116 122068 169168 122120
rect 214564 122068 214616 122120
rect 203616 121456 203668 121508
rect 213920 121456 213972 121508
rect 253480 121456 253532 121508
rect 264980 121456 265032 121508
rect 231768 121388 231820 121440
rect 255964 121388 256016 121440
rect 282828 121388 282880 121440
rect 302424 121388 302476 121440
rect 231676 120912 231728 120964
rect 238024 120912 238076 120964
rect 193956 120164 194008 120216
rect 213920 120164 213972 120216
rect 177580 120096 177632 120148
rect 214012 120096 214064 120148
rect 260288 120096 260340 120148
rect 264980 120096 265032 120148
rect 231768 120028 231820 120080
rect 258724 120028 258776 120080
rect 282828 120028 282880 120080
rect 302240 120028 302292 120080
rect 282736 119960 282788 120012
rect 288532 119960 288584 120012
rect 211804 118736 211856 118788
rect 214012 118736 214064 118788
rect 263140 118736 263192 118788
rect 265440 118736 265492 118788
rect 176108 118668 176160 118720
rect 213920 118668 213972 118720
rect 231216 118668 231268 118720
rect 238116 118668 238168 118720
rect 255964 118668 256016 118720
rect 264980 118668 265032 118720
rect 231400 118600 231452 118652
rect 251916 118600 251968 118652
rect 282828 118600 282880 118652
rect 309232 118600 309284 118652
rect 282276 118532 282328 118584
rect 292672 118532 292724 118584
rect 238392 117920 238444 117972
rect 249156 117920 249208 117972
rect 231492 117648 231544 117700
rect 236644 117648 236696 117700
rect 206468 117376 206520 117428
rect 213920 117376 213972 117428
rect 254584 117376 254636 117428
rect 264980 117376 265032 117428
rect 170404 117308 170456 117360
rect 214012 117308 214064 117360
rect 249064 117308 249116 117360
rect 265072 117308 265124 117360
rect 231768 117240 231820 117292
rect 241152 117240 241204 117292
rect 282828 117240 282880 117292
rect 303712 117240 303764 117292
rect 231676 116832 231728 116884
rect 235264 116832 235316 116884
rect 199476 116016 199528 116068
rect 213920 116016 213972 116068
rect 240784 116016 240836 116068
rect 265072 116016 265124 116068
rect 177304 115948 177356 116000
rect 214012 115948 214064 116000
rect 236644 115948 236696 116000
rect 264980 115948 265032 116000
rect 231492 115880 231544 115932
rect 264336 115880 264388 115932
rect 282368 115880 282420 115932
rect 305092 115880 305144 115932
rect 282828 115812 282880 115864
rect 303896 115812 303948 115864
rect 168288 115200 168340 115252
rect 183008 115200 183060 115252
rect 203524 114588 203576 114640
rect 214012 114588 214064 114640
rect 230572 114588 230624 114640
rect 232688 114588 232740 114640
rect 183100 114520 183152 114572
rect 213920 114520 213972 114572
rect 249156 114520 249208 114572
rect 264980 114520 265032 114572
rect 231768 114452 231820 114504
rect 267096 114452 267148 114504
rect 282092 114452 282144 114504
rect 307760 114452 307812 114504
rect 231492 114384 231544 114436
rect 241060 114384 241112 114436
rect 167736 113772 167788 113824
rect 184388 113772 184440 113824
rect 261668 113568 261720 113620
rect 264980 113568 265032 113620
rect 211988 113296 212040 113348
rect 214288 113296 214340 113348
rect 184480 113160 184532 113212
rect 213920 113160 213972 113212
rect 231768 113092 231820 113144
rect 262956 113092 263008 113144
rect 282828 113092 282880 113144
rect 291200 113092 291252 113144
rect 231400 113024 231452 113076
rect 249248 113024 249300 113076
rect 282460 113024 282512 113076
rect 285772 113024 285824 113076
rect 202512 112412 202564 112464
rect 214748 112412 214800 112464
rect 210516 111800 210568 111852
rect 213920 111800 213972 111852
rect 260380 111800 260432 111852
rect 264980 111800 265032 111852
rect 230756 111732 230808 111784
rect 234068 111732 234120 111784
rect 282828 111732 282880 111784
rect 289820 111732 289872 111784
rect 281724 111596 281776 111648
rect 284300 111596 284352 111648
rect 231584 111052 231636 111104
rect 250812 111052 250864 111104
rect 177488 110508 177540 110560
rect 213920 110508 213972 110560
rect 261484 110508 261536 110560
rect 265072 110508 265124 110560
rect 167644 110440 167696 110492
rect 214012 110440 214064 110492
rect 247776 110440 247828 110492
rect 264980 110440 265032 110492
rect 231768 110372 231820 110424
rect 242164 110372 242216 110424
rect 282276 110372 282328 110424
rect 299572 110372 299624 110424
rect 282828 110304 282880 110356
rect 298100 110304 298152 110356
rect 231400 109692 231452 109744
rect 249340 109692 249392 109744
rect 173348 109080 173400 109132
rect 213920 109080 213972 109132
rect 251824 109080 251876 109132
rect 265072 109080 265124 109132
rect 171968 109012 172020 109064
rect 214012 109012 214064 109064
rect 242256 109012 242308 109064
rect 264980 109012 265032 109064
rect 168012 108944 168064 108996
rect 169208 108944 169260 108996
rect 231584 108944 231636 108996
rect 256056 108944 256108 108996
rect 282368 108944 282420 108996
rect 295524 108944 295576 108996
rect 231768 108536 231820 108588
rect 236920 108536 236972 108588
rect 192668 108264 192720 108316
rect 202420 108264 202472 108316
rect 236736 108264 236788 108316
rect 246396 108264 246448 108316
rect 282828 107924 282880 107976
rect 287152 107924 287204 107976
rect 202328 107720 202380 107772
rect 213920 107720 213972 107772
rect 258724 107720 258776 107772
rect 265072 107720 265124 107772
rect 165068 107652 165120 107704
rect 214012 107652 214064 107704
rect 250536 107652 250588 107704
rect 264980 107652 265032 107704
rect 231308 107584 231360 107636
rect 259092 107584 259144 107636
rect 231768 107516 231820 107568
rect 239680 107516 239732 107568
rect 209228 106360 209280 106412
rect 214012 106360 214064 106412
rect 258908 106360 258960 106412
rect 265072 106360 265124 106412
rect 181628 106292 181680 106344
rect 213920 106292 213972 106344
rect 252100 106292 252152 106344
rect 264980 106292 265032 106344
rect 231400 106224 231452 106276
rect 262864 106224 262916 106276
rect 282828 106224 282880 106276
rect 291292 106224 291344 106276
rect 231768 106156 231820 106208
rect 247960 106156 248012 106208
rect 166540 105544 166592 105596
rect 203616 105544 203668 105596
rect 205180 104932 205232 104984
rect 213920 104932 213972 104984
rect 262956 104932 263008 104984
rect 265072 104932 265124 104984
rect 176016 104864 176068 104916
rect 214012 104864 214064 104916
rect 253572 104864 253624 104916
rect 264980 104864 265032 104916
rect 282828 104796 282880 104848
rect 292580 104796 292632 104848
rect 231768 104728 231820 104780
rect 238300 104728 238352 104780
rect 231124 104320 231176 104372
rect 235356 104320 235408 104372
rect 181536 103572 181588 103624
rect 214012 103572 214064 103624
rect 170496 103504 170548 103556
rect 213920 103504 213972 103556
rect 238116 103504 238168 103556
rect 264980 103504 265032 103556
rect 231768 103436 231820 103488
rect 240968 103436 241020 103488
rect 282828 103436 282880 103488
rect 290004 103436 290056 103488
rect 241060 102824 241112 102876
rect 263140 102824 263192 102876
rect 169208 102756 169260 102808
rect 213184 102756 213236 102808
rect 231032 102756 231084 102808
rect 256332 102756 256384 102808
rect 262772 102212 262824 102264
rect 265164 102212 265216 102264
rect 256148 102144 256200 102196
rect 264980 102144 265032 102196
rect 231676 102076 231728 102128
rect 254768 102076 254820 102128
rect 230572 102008 230624 102060
rect 242348 102008 242400 102060
rect 281724 102008 281776 102060
rect 284392 102008 284444 102060
rect 173440 101396 173492 101448
rect 189816 101396 189868 101448
rect 169300 100716 169352 100768
rect 213920 100716 213972 100768
rect 246396 100716 246448 100768
rect 264980 100716 265032 100768
rect 230572 100648 230624 100700
rect 263048 100648 263100 100700
rect 281724 100648 281776 100700
rect 302332 100648 302384 100700
rect 231124 100580 231176 100632
rect 238208 100580 238260 100632
rect 211896 99424 211948 99476
rect 214012 99424 214064 99476
rect 263140 99424 263192 99476
rect 265072 99424 265124 99476
rect 170680 99356 170732 99408
rect 213920 99356 213972 99408
rect 257620 99356 257672 99408
rect 264980 99356 265032 99408
rect 231124 99288 231176 99340
rect 236828 99288 236880 99340
rect 282828 99288 282880 99340
rect 310520 99288 310572 99340
rect 231676 98608 231728 98660
rect 246304 98608 246356 98660
rect 253388 98064 253440 98116
rect 265072 98064 265124 98116
rect 167828 97996 167880 98048
rect 213920 97996 213972 98048
rect 246580 97996 246632 98048
rect 264980 97996 265032 98048
rect 3424 97928 3476 97980
rect 17224 97928 17276 97980
rect 231768 97928 231820 97980
rect 259000 97928 259052 97980
rect 282184 97928 282236 97980
rect 298376 97928 298428 97980
rect 282828 97860 282880 97912
rect 295432 97860 295484 97912
rect 177396 97248 177448 97300
rect 214840 97248 214892 97300
rect 206284 96636 206336 96688
rect 213920 96636 213972 96688
rect 214472 96636 214524 96688
rect 264980 97248 265032 97300
rect 219164 96024 219216 96076
rect 219256 96024 219308 96076
rect 259092 96636 259144 96688
rect 265072 96636 265124 96688
rect 209136 95956 209188 96008
rect 220084 95956 220136 96008
rect 164976 95888 165028 95940
rect 214104 95888 214156 95940
rect 230572 95820 230624 95872
rect 232596 95820 232648 95872
rect 224408 95208 224460 95260
rect 227720 95208 227772 95260
rect 230572 95208 230624 95260
rect 240140 95208 240192 95260
rect 260104 95140 260156 95192
rect 278780 95140 278832 95192
rect 67364 94460 67416 94512
rect 124864 94460 124916 94512
rect 135812 94460 135864 94512
rect 167736 94460 167788 94512
rect 191288 94460 191340 94512
rect 213368 94460 213420 94512
rect 217324 94460 217376 94512
rect 253480 94460 253532 94512
rect 267648 94460 267700 94512
rect 269120 94460 269172 94512
rect 100668 93848 100720 93900
rect 166448 93848 166500 93900
rect 228364 93848 228416 93900
rect 229836 93848 229888 93900
rect 213276 93780 213328 93832
rect 281632 93780 281684 93832
rect 217232 93712 217284 93764
rect 230480 93712 230532 93764
rect 240140 93712 240192 93764
rect 273996 93712 274048 93764
rect 67548 93168 67600 93220
rect 97264 93168 97316 93220
rect 117136 93168 117188 93220
rect 177580 93168 177632 93220
rect 185768 93168 185820 93220
rect 202512 93168 202564 93220
rect 65984 93100 66036 93152
rect 106924 93100 106976 93152
rect 121736 93100 121788 93152
rect 187148 93100 187200 93152
rect 106832 92556 106884 92608
rect 116584 92556 116636 92608
rect 99104 92488 99156 92540
rect 112444 92488 112496 92540
rect 110696 92420 110748 92472
rect 133880 92420 133932 92472
rect 136088 92420 136140 92472
rect 166356 92420 166408 92472
rect 267188 92420 267240 92472
rect 281540 92420 281592 92472
rect 159364 91808 159416 91860
rect 181444 91808 181496 91860
rect 214656 91808 214708 91860
rect 265808 91808 265860 91860
rect 59176 91740 59228 91792
rect 88984 91740 89036 91792
rect 180156 91740 180208 91792
rect 253572 91740 253624 91792
rect 84384 91196 84436 91248
rect 111064 91196 111116 91248
rect 89076 91128 89128 91180
rect 104256 91128 104308 91180
rect 109684 91060 109736 91112
rect 115204 91060 115256 91112
rect 151452 91060 151504 91112
rect 157340 91060 157392 91112
rect 111524 90992 111576 91044
rect 170404 90992 170456 91044
rect 124128 90924 124180 90976
rect 169116 90924 169168 90976
rect 205088 90380 205140 90432
rect 232780 90380 232832 90432
rect 169024 90312 169076 90364
rect 206284 90312 206336 90364
rect 218704 90312 218756 90364
rect 256148 90312 256200 90364
rect 119804 89632 119856 89684
rect 166540 89632 166592 89684
rect 157340 89564 157392 89616
rect 185676 89564 185728 89616
rect 206284 89020 206336 89072
rect 234160 89020 234212 89072
rect 67272 88952 67324 89004
rect 108304 88952 108356 89004
rect 178960 88952 179012 89004
rect 198096 88952 198148 89004
rect 227076 88952 227128 89004
rect 257620 88952 257672 89004
rect 174728 88816 174780 88868
rect 178868 88816 178920 88868
rect 105544 88272 105596 88324
rect 183100 88272 183152 88324
rect 120724 88204 120776 88256
rect 166264 88204 166316 88256
rect 213184 87660 213236 87712
rect 260380 87660 260432 87712
rect 66168 87592 66220 87644
rect 107016 87592 107068 87644
rect 173256 87592 173308 87644
rect 192668 87592 192720 87644
rect 198096 87592 198148 87644
rect 250720 87592 250772 87644
rect 112720 86912 112772 86964
rect 189908 86912 189960 86964
rect 152464 86844 152516 86896
rect 171876 86844 171928 86896
rect 188436 86300 188488 86352
rect 223028 86300 223080 86352
rect 67732 86232 67784 86284
rect 150440 86232 150492 86284
rect 196716 86232 196768 86284
rect 236920 86232 236972 86284
rect 3148 85484 3200 85536
rect 14464 85484 14516 85536
rect 104440 85484 104492 85536
rect 184480 85484 184532 85536
rect 115756 85416 115808 85468
rect 193956 85416 194008 85468
rect 225604 84872 225656 84924
rect 232688 84872 232740 84924
rect 49608 84804 49660 84856
rect 83464 84804 83516 84856
rect 195244 84804 195296 84856
rect 281540 84804 281592 84856
rect 97816 84124 97868 84176
rect 171968 84124 172020 84176
rect 126796 84056 126848 84108
rect 185768 84056 185820 84108
rect 222844 83512 222896 83564
rect 249248 83512 249300 83564
rect 86868 83444 86920 83496
rect 126244 83444 126296 83496
rect 211804 83444 211856 83496
rect 239588 83444 239640 83496
rect 88248 82764 88300 82816
rect 170680 82764 170732 82816
rect 111064 82696 111116 82748
rect 169300 82696 169352 82748
rect 195244 82084 195296 82136
rect 247868 82084 247920 82136
rect 67640 81336 67692 81388
rect 181536 81336 181588 81388
rect 95148 81268 95200 81320
rect 202328 81268 202380 81320
rect 204904 80656 204956 80708
rect 235448 80656 235500 80708
rect 97908 79976 97960 80028
rect 195336 79976 195388 80028
rect 126888 79908 126940 79960
rect 159364 79908 159416 79960
rect 224316 79296 224368 79348
rect 238392 79296 238444 79348
rect 122748 78616 122800 78668
rect 174636 78616 174688 78668
rect 151636 78548 151688 78600
rect 169208 78548 169260 78600
rect 175924 77936 175976 77988
rect 273260 77936 273312 77988
rect 128268 77188 128320 77240
rect 173440 77188 173492 77240
rect 106188 76508 106240 76560
rect 240876 76508 240928 76560
rect 107016 75828 107068 75880
rect 178960 75828 179012 75880
rect 111708 75148 111760 75200
rect 229928 75148 229980 75200
rect 91008 74468 91060 74520
rect 176016 74468 176068 74520
rect 117228 73788 117280 73840
rect 252008 73788 252060 73840
rect 151544 73108 151596 73160
rect 192576 73108 192628 73160
rect 126244 73040 126296 73092
rect 164976 73040 165028 73092
rect 583852 72768 583904 72820
rect 583852 72564 583904 72616
rect 3424 71680 3476 71732
rect 22744 71680 22796 71732
rect 99196 71680 99248 71732
rect 177488 71680 177540 71732
rect 119988 71000 120040 71052
rect 250628 71000 250680 71052
rect 102048 70320 102100 70372
rect 210516 70320 210568 70372
rect 125416 70252 125468 70304
rect 180248 70252 180300 70304
rect 103428 68960 103480 69012
rect 164884 68960 164936 69012
rect 101404 68280 101456 68332
rect 254676 68280 254728 68332
rect 107568 67532 107620 67584
rect 203524 67532 203576 67584
rect 116584 67464 116636 67516
rect 173256 67464 173308 67516
rect 108304 66172 108356 66224
rect 214748 66172 214800 66224
rect 106096 66104 106148 66156
rect 182916 66104 182968 66156
rect 104256 64812 104308 64864
rect 211896 64812 211948 64864
rect 124036 64744 124088 64796
rect 191104 64744 191156 64796
rect 125508 63452 125560 63504
rect 206376 63452 206428 63504
rect 124864 63384 124916 63436
rect 169024 63384 169076 63436
rect 132408 62024 132460 62076
rect 198188 62024 198240 62076
rect 115848 61956 115900 62008
rect 171784 61956 171836 62008
rect 114376 60664 114428 60716
rect 189724 60664 189776 60716
rect 77208 59984 77260 60036
rect 258908 59984 258960 60036
rect 3056 59304 3108 59356
rect 33784 59304 33836 59356
rect 129648 59304 129700 59356
rect 202236 59304 202288 59356
rect 79968 58624 80020 58676
rect 252100 58624 252152 58676
rect 112444 57876 112496 57928
rect 210424 57876 210476 57928
rect 93768 57196 93820 57248
rect 231216 57196 231268 57248
rect 110144 56516 110196 56568
rect 206468 56516 206520 56568
rect 91008 55836 91060 55888
rect 250536 55836 250588 55888
rect 115204 55156 115256 55208
rect 177304 55156 177356 55208
rect 97908 54476 97960 54528
rect 242256 54476 242308 54528
rect 118516 53728 118568 53780
rect 191288 53728 191340 53780
rect 47584 53048 47636 53100
rect 101404 53048 101456 53100
rect 102048 53048 102100 53100
rect 267740 53048 267792 53100
rect 114284 52368 114336 52420
rect 174728 52368 174780 52420
rect 199384 51756 199436 51808
rect 240140 51756 240192 51808
rect 108948 51688 109000 51740
rect 264336 51688 264388 51740
rect 119896 51008 119948 51060
rect 192484 51008 192536 51060
rect 103428 50328 103480 50380
rect 239404 50328 239456 50380
rect 115848 49036 115900 49088
rect 247776 49036 247828 49088
rect 38568 48968 38620 49020
rect 236644 48968 236696 49020
rect 118608 48220 118660 48272
rect 177396 48220 177448 48272
rect 180064 47608 180116 47660
rect 222936 47608 222988 47660
rect 146944 47540 146996 47592
rect 218704 47540 218756 47592
rect 223028 47540 223080 47592
rect 267740 47540 267792 47592
rect 97264 46248 97316 46300
rect 227076 46248 227128 46300
rect 45376 46180 45428 46232
rect 262864 46180 262916 46232
rect 3424 45500 3476 45552
rect 21364 45500 21416 45552
rect 125508 44888 125560 44940
rect 236736 44888 236788 44940
rect 86776 44820 86828 44872
rect 251916 44820 251968 44872
rect 174544 43460 174596 43512
rect 241520 43460 241572 43512
rect 88248 43392 88300 43444
rect 205088 43392 205140 43444
rect 231216 43392 231268 43444
rect 269120 43392 269172 43444
rect 56508 42100 56560 42152
rect 249064 42100 249116 42152
rect 19248 42032 19300 42084
rect 235356 42032 235408 42084
rect 62028 40672 62080 40724
rect 324412 40672 324464 40724
rect 112444 39380 112496 39432
rect 230480 39380 230532 39432
rect 53656 39312 53708 39364
rect 254584 39312 254636 39364
rect 62028 37952 62080 38004
rect 260196 37952 260248 38004
rect 30288 37884 30340 37936
rect 242164 37884 242216 37936
rect 60648 36592 60700 36644
rect 248420 36592 248472 36644
rect 49608 36524 49660 36576
rect 267004 36524 267056 36576
rect 111616 35232 111668 35284
rect 261484 35232 261536 35284
rect 43996 35164 44048 35216
rect 253204 35164 253256 35216
rect 71044 33804 71096 33856
rect 215944 33804 215996 33856
rect 59176 33736 59228 33788
rect 267096 33736 267148 33788
rect 2872 33056 2924 33108
rect 36544 33056 36596 33108
rect 110328 32444 110380 32496
rect 243544 32444 243596 32496
rect 50988 32376 51040 32428
rect 249800 32376 249852 32428
rect 83464 31084 83516 31136
rect 267004 31084 267056 31136
rect 37096 31016 37148 31068
rect 245108 31016 245160 31068
rect 55036 29588 55088 29640
rect 233976 29588 234028 29640
rect 184296 28296 184348 28348
rect 258080 28296 258132 28348
rect 122748 28228 122800 28280
rect 213184 28228 213236 28280
rect 83464 26936 83516 26988
rect 238116 26936 238168 26988
rect 95056 26868 95108 26920
rect 258724 26868 258776 26920
rect 20628 25576 20680 25628
rect 221464 25576 221516 25628
rect 63408 25508 63460 25560
rect 310520 25508 310572 25560
rect 188528 24148 188580 24200
rect 263600 24148 263652 24200
rect 82728 24080 82780 24132
rect 222844 24080 222896 24132
rect 84108 22720 84160 22772
rect 231124 22720 231176 22772
rect 126244 21428 126296 21480
rect 217324 21428 217376 21480
rect 31668 21360 31720 21412
rect 235264 21360 235316 21412
rect 3424 20612 3476 20664
rect 51724 20612 51776 20664
rect 100668 20000 100720 20052
rect 196716 20000 196768 20052
rect 55128 19932 55180 19984
rect 317420 19932 317472 19984
rect 96528 18640 96580 18692
rect 224224 18640 224276 18692
rect 48228 18572 48280 18624
rect 289820 18572 289872 18624
rect 13728 17280 13780 17332
rect 250444 17280 250496 17332
rect 44088 17212 44140 17264
rect 296720 17212 296772 17264
rect 61936 15920 61988 15972
rect 195244 15920 195296 15972
rect 200764 15920 200816 15972
rect 253480 15920 253532 15972
rect 27528 15852 27580 15904
rect 220176 15852 220228 15904
rect 318064 15852 318116 15904
rect 328736 15852 328788 15904
rect 85488 14492 85540 14544
rect 181444 14492 181496 14544
rect 209044 14492 209096 14544
rect 299664 14492 299716 14544
rect 12164 14424 12216 14476
rect 226984 14424 227036 14476
rect 1676 13132 1728 13184
rect 112444 13132 112496 13184
rect 118608 13132 118660 13184
rect 229744 13132 229796 13184
rect 60648 13064 60700 13116
rect 206284 13064 206336 13116
rect 214564 13064 214616 13116
rect 307944 13064 307996 13116
rect 71504 11772 71556 11824
rect 209136 11772 209188 11824
rect 39948 11704 40000 11756
rect 251180 11704 251232 11756
rect 332692 11704 332744 11756
rect 333888 11704 333940 11756
rect 112812 10344 112864 10396
rect 204904 10344 204956 10396
rect 104532 10276 104584 10328
rect 251824 10276 251876 10328
rect 77392 8984 77444 9036
rect 228364 8984 228416 9036
rect 19432 8916 19484 8968
rect 104164 8916 104216 8968
rect 107016 8916 107068 8968
rect 142804 8916 142856 8968
rect 186964 8916 187016 8968
rect 346952 8916 347004 8968
rect 66720 7624 66772 7676
rect 238024 7624 238076 7676
rect 41880 7556 41932 7608
rect 233884 7556 233936 7608
rect 119896 6196 119948 6248
rect 224316 6196 224368 6248
rect 47860 6128 47912 6180
rect 146944 6128 146996 6180
rect 178776 6128 178828 6180
rect 303160 6128 303212 6180
rect 340972 6128 341024 6180
rect 349160 6128 349212 6180
rect 232596 5516 232648 5568
rect 235816 5516 235868 5568
rect 69112 4836 69164 4888
rect 180156 4836 180208 4888
rect 45468 4768 45520 4820
rect 240784 4768 240836 4820
rect 313832 4428 313884 4480
rect 316040 4428 316092 4480
rect 11152 3544 11204 3596
rect 12256 3544 12308 3596
rect 27712 3544 27764 3596
rect 2872 3476 2924 3528
rect 3976 3476 4028 3528
rect 8760 3476 8812 3528
rect 9588 3476 9640 3528
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 15936 3476 15988 3528
rect 16488 3476 16540 3528
rect 17040 3476 17092 3528
rect 17868 3476 17920 3528
rect 18236 3476 18288 3528
rect 19248 3476 19300 3528
rect 24216 3476 24268 3528
rect 24768 3476 24820 3528
rect 25320 3476 25372 3528
rect 26148 3476 26200 3528
rect 26516 3476 26568 3528
rect 27528 3476 27580 3528
rect 32404 3476 32456 3528
rect 33048 3476 33100 3528
rect 33600 3476 33652 3528
rect 34428 3476 34480 3528
rect 35992 3544 36044 3596
rect 37096 3544 37148 3596
rect 47584 3476 47636 3528
rect 48964 3476 49016 3528
rect 49608 3476 49660 3528
rect 50160 3476 50212 3528
rect 50896 3476 50948 3528
rect 56048 3476 56100 3528
rect 56508 3476 56560 3528
rect 57244 3476 57296 3528
rect 57888 3476 57940 3528
rect 58440 3476 58492 3528
rect 59176 3476 59228 3528
rect 59636 3476 59688 3528
rect 60648 3476 60700 3528
rect 63224 3476 63276 3528
rect 71044 3544 71096 3596
rect 85672 3544 85724 3596
rect 86776 3544 86828 3596
rect 65524 3476 65576 3528
rect 66168 3476 66220 3528
rect 67916 3476 67968 3528
rect 68928 3476 68980 3528
rect 72608 3476 72660 3528
rect 73068 3476 73120 3528
rect 73804 3476 73856 3528
rect 74448 3476 74500 3528
rect 75000 3476 75052 3528
rect 75828 3476 75880 3528
rect 76196 3476 76248 3528
rect 77208 3476 77260 3528
rect 80888 3476 80940 3528
rect 81348 3476 81400 3528
rect 82084 3476 82136 3528
rect 82728 3476 82780 3528
rect 83280 3476 83332 3528
rect 84108 3476 84160 3528
rect 84476 3476 84528 3528
rect 85488 3476 85540 3528
rect 90364 3476 90416 3528
rect 91008 3476 91060 3528
rect 91560 3476 91612 3528
rect 126244 3544 126296 3596
rect 276020 3544 276072 3596
rect 277124 3544 277176 3596
rect 123484 3476 123536 3528
rect 124128 3476 124180 3528
rect 124680 3476 124732 3528
rect 125508 3476 125560 3528
rect 129372 3476 129424 3528
rect 130384 3476 130436 3528
rect 202144 3476 202196 3528
rect 257068 3476 257120 3528
rect 281448 3476 281500 3528
rect 283104 3476 283156 3528
rect 296076 3476 296128 3528
rect 299480 3476 299532 3528
rect 307760 3476 307812 3528
rect 309048 3476 309100 3528
rect 313924 3476 313976 3528
rect 315028 3476 315080 3528
rect 324320 3476 324372 3528
rect 325608 3476 325660 3528
rect 336004 3476 336056 3528
rect 337476 3476 337528 3528
rect 340880 3476 340932 3528
rect 342168 3476 342220 3528
rect 582196 3476 582248 3528
rect 583392 3476 583444 3528
rect 6460 3408 6512 3460
rect 29644 3408 29696 3460
rect 34796 3408 34848 3460
rect 35808 3408 35860 3460
rect 40684 3408 40736 3460
rect 41328 3408 41380 3460
rect 43076 3408 43128 3460
rect 43996 3408 44048 3460
rect 44272 3408 44324 3460
rect 45376 3408 45428 3460
rect 51356 3408 51408 3460
rect 78588 3408 78640 3460
rect 87604 3408 87656 3460
rect 92756 3408 92808 3460
rect 93768 3408 93820 3460
rect 93952 3408 94004 3460
rect 95056 3408 95108 3460
rect 97448 3408 97500 3460
rect 97908 3408 97960 3460
rect 98644 3408 98696 3460
rect 99288 3408 99340 3460
rect 99840 3408 99892 3460
rect 100668 3408 100720 3460
rect 101036 3408 101088 3460
rect 102048 3408 102100 3460
rect 105728 3408 105780 3460
rect 106188 3408 106240 3460
rect 108120 3408 108172 3460
rect 108948 3408 109000 3460
rect 109316 3408 109368 3460
rect 110328 3408 110380 3460
rect 110512 3408 110564 3460
rect 111708 3408 111760 3460
rect 115204 3408 115256 3460
rect 115848 3408 115900 3460
rect 116400 3408 116452 3460
rect 117228 3408 117280 3460
rect 117596 3408 117648 3460
rect 118608 3408 118660 3460
rect 118792 3408 118844 3460
rect 119988 3408 120040 3460
rect 83464 3340 83516 3392
rect 114008 3340 114060 3392
rect 214656 3408 214708 3460
rect 257344 3408 257396 3460
rect 266544 3408 266596 3460
rect 267004 3408 267056 3460
rect 274824 3408 274876 3460
rect 285404 3408 285456 3460
rect 306472 3408 306524 3460
rect 315304 3408 315356 3460
rect 323308 3408 323360 3460
rect 351644 3408 351696 3460
rect 358820 3408 358872 3460
rect 52552 3272 52604 3324
rect 53656 3272 53708 3324
rect 89168 3272 89220 3324
rect 89628 3272 89680 3324
rect 122288 3272 122340 3324
rect 122748 3272 122800 3324
rect 350448 3136 350500 3188
rect 353300 3136 353352 3188
rect 269764 3068 269816 3120
rect 272432 3068 272484 3120
rect 314016 3068 314068 3120
rect 317328 3068 317380 3120
rect 581000 3068 581052 3120
rect 583576 3068 583628 3120
rect 60832 3000 60884 3052
rect 61936 3000 61988 3052
rect 347044 3000 347096 3052
rect 349252 3000 349304 3052
rect 222936 2728 222988 2780
rect 292580 2796 292632 2848
rect 28908 2116 28960 2168
rect 106832 2116 106884 2168
rect 121092 2116 121144 2168
rect 198096 2116 198148 2168
rect 7656 2048 7708 2100
rect 40592 2048 40644 2100
rect 102232 2048 102284 2100
rect 231216 2048 231268 2100
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 702642 8156 703520
rect 8116 702636 8168 702642
rect 8116 702578 8168 702584
rect 24320 698970 24348 703520
rect 24308 698964 24360 698970
rect 24308 698906 24360 698912
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 18604 683188 18656 683194
rect 18604 683130 18656 683136
rect 3422 671256 3478 671265
rect 3422 671191 3478 671200
rect 3436 639606 3464 671191
rect 3514 658200 3570 658209
rect 3514 658135 3570 658144
rect 3528 656946 3556 658135
rect 3516 656940 3568 656946
rect 3516 656882 3568 656888
rect 3424 639600 3476 639606
rect 3424 639542 3476 639548
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 11704 632120 11756 632126
rect 3476 632088 3478 632097
rect 11704 632062 11756 632068
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 600982 3280 606047
rect 3240 600976 3292 600982
rect 3240 600918 3292 600924
rect 3424 590028 3476 590034
rect 3424 589970 3476 589976
rect 3436 580009 3464 589970
rect 3422 580000 3478 580009
rect 3422 579935 3478 579944
rect 11716 576162 11744 632062
rect 15844 618316 15896 618322
rect 15844 618258 15896 618264
rect 11704 576156 11756 576162
rect 11704 576098 11756 576104
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 2778 553888 2834 553897
rect 2778 553823 2780 553832
rect 2832 553823 2834 553832
rect 2780 553794 2832 553800
rect 3436 540258 3464 566879
rect 4804 553852 4856 553858
rect 4804 553794 4856 553800
rect 3424 540252 3476 540258
rect 3424 540194 3476 540200
rect 3424 538892 3476 538898
rect 3424 538834 3476 538840
rect 3436 527921 3464 538834
rect 4816 538218 4844 553794
rect 4804 538212 4856 538218
rect 4804 538154 4856 538160
rect 15856 536110 15884 618258
rect 18616 543046 18644 683130
rect 22744 656940 22796 656946
rect 22744 656882 22796 656888
rect 22756 592686 22784 656882
rect 39304 639600 39356 639606
rect 39304 639542 39356 639548
rect 22744 592680 22796 592686
rect 22744 592622 22796 592628
rect 18604 543040 18656 543046
rect 18604 542982 18656 542988
rect 39316 541686 39344 639542
rect 40052 598262 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 67640 703520 67692 703526
rect 72946 703520 73058 704960
rect 75828 703656 75880 703662
rect 75828 703598 75880 703604
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 67640 703462 67692 703468
rect 59268 703384 59320 703390
rect 59268 703326 59320 703332
rect 57704 702976 57756 702982
rect 57704 702918 57756 702924
rect 53748 702568 53800 702574
rect 53748 702510 53800 702516
rect 40040 598256 40092 598262
rect 40040 598198 40092 598204
rect 50988 585200 51040 585206
rect 50988 585142 51040 585148
rect 48136 582412 48188 582418
rect 48136 582354 48188 582360
rect 41328 572756 41380 572762
rect 41328 572698 41380 572704
rect 39948 543040 40000 543046
rect 39948 542982 40000 542988
rect 39960 542434 39988 542982
rect 39948 542428 40000 542434
rect 39948 542370 40000 542376
rect 39304 541680 39356 541686
rect 39304 541622 39356 541628
rect 15844 536104 15896 536110
rect 15844 536046 15896 536052
rect 7564 534744 7616 534750
rect 7564 534686 7616 534692
rect 5448 533384 5500 533390
rect 5448 533326 5500 533332
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3332 502104 3384 502110
rect 3332 502046 3384 502052
rect 3344 501809 3372 502046
rect 3330 501800 3386 501809
rect 3330 501735 3386 501744
rect 2778 462632 2834 462641
rect 2778 462567 2780 462576
rect 2832 462567 2834 462576
rect 2780 462538 2832 462544
rect 3436 451926 3464 527847
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 3516 514762 3568 514768
rect 4066 475688 4122 475697
rect 4066 475623 4122 475632
rect 4080 475386 4108 475623
rect 5460 475386 5488 533326
rect 7576 502110 7604 534686
rect 15844 530596 15896 530602
rect 15844 530538 15896 530544
rect 14464 514820 14516 514826
rect 14464 514762 14516 514768
rect 7564 502104 7616 502110
rect 7564 502046 7616 502052
rect 4068 475380 4120 475386
rect 4068 475322 4120 475328
rect 5448 475380 5500 475386
rect 5448 475322 5500 475328
rect 11704 475380 11756 475386
rect 11704 475322 11756 475328
rect 4804 462596 4856 462602
rect 4804 462538 4856 462544
rect 3424 451920 3476 451926
rect 3424 451862 3476 451868
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 4816 447846 4844 462538
rect 4804 447840 4856 447846
rect 4804 447782 4856 447788
rect 4804 444440 4856 444446
rect 4804 444382 4856 444388
rect 3146 423600 3202 423609
rect 3146 423535 3202 423544
rect 3160 422958 3188 423535
rect 3148 422952 3200 422958
rect 3148 422894 3200 422900
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 2780 398744 2832 398750
rect 2780 398686 2832 398692
rect 2792 397497 2820 398686
rect 2778 397488 2834 397497
rect 2778 397423 2834 397432
rect 3436 388929 3464 410479
rect 4816 398750 4844 444382
rect 4804 398744 4856 398750
rect 4804 398686 4856 398692
rect 11716 389230 11744 475322
rect 14476 451246 14504 514762
rect 14464 451240 14516 451246
rect 14464 451182 14516 451188
rect 14464 448588 14516 448594
rect 14464 448530 14516 448536
rect 11704 389224 11756 389230
rect 11704 389166 11756 389172
rect 3422 388920 3478 388929
rect 3422 388855 3478 388864
rect 3422 387016 3478 387025
rect 3422 386951 3478 386960
rect 3436 383654 3464 386951
rect 5448 384328 5500 384334
rect 5448 384270 5500 384276
rect 3436 383626 3556 383654
rect 3528 371385 3556 383626
rect 3514 371376 3570 371385
rect 3514 371311 3570 371320
rect 3332 358760 3384 358766
rect 3332 358702 3384 358708
rect 3344 358465 3372 358702
rect 3330 358456 3386 358465
rect 3330 358391 3386 358400
rect 3424 347064 3476 347070
rect 3424 347006 3476 347012
rect 3148 346384 3200 346390
rect 3148 346326 3200 346332
rect 3160 345409 3188 346326
rect 3146 345400 3202 345409
rect 3146 345335 3202 345344
rect 20 326392 72 326398
rect 20 326334 72 326340
rect 32 6769 60 326334
rect 2778 293176 2834 293185
rect 2778 293111 2834 293120
rect 2792 292874 2820 293111
rect 2780 292868 2832 292874
rect 2780 292810 2832 292816
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3436 214985 3464 347006
rect 3528 318102 3556 371311
rect 5460 319462 5488 384270
rect 7562 381576 7618 381585
rect 7562 381511 7618 381520
rect 7576 346390 7604 381511
rect 7564 346384 7616 346390
rect 7564 346326 7616 346332
rect 7562 328536 7618 328545
rect 7562 328471 7618 328480
rect 4068 319456 4120 319462
rect 4068 319398 4120 319404
rect 5448 319456 5500 319462
rect 5448 319398 5500 319404
rect 4080 319297 4108 319398
rect 4066 319288 4122 319297
rect 4066 319223 4122 319232
rect 3516 318096 3568 318102
rect 3516 318038 3568 318044
rect 3516 306332 3568 306338
rect 3516 306274 3568 306280
rect 3528 306241 3556 306274
rect 3514 306232 3570 306241
rect 3514 306167 3570 306176
rect 4804 292868 4856 292874
rect 4804 292810 4856 292816
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3528 267034 3556 267135
rect 3516 267028 3568 267034
rect 3516 266970 3568 266976
rect 3516 241460 3568 241466
rect 3516 241402 3568 241408
rect 3528 241097 3556 241402
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 4816 237289 4844 292810
rect 4802 237280 4858 237289
rect 4802 237215 4858 237224
rect 4804 220856 4856 220862
rect 4804 220798 4856 220804
rect 3422 214976 3478 214985
rect 3422 214911 3478 214920
rect 3422 210352 3478 210361
rect 3422 210287 3478 210296
rect 3056 202836 3108 202842
rect 3056 202778 3108 202784
rect 3068 201929 3096 202778
rect 3054 201920 3110 201929
rect 3054 201855 3110 201864
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 2780 150340 2832 150346
rect 2780 150282 2832 150288
rect 2792 149841 2820 150282
rect 2778 149832 2834 149841
rect 2778 149767 2834 149776
rect 3436 110673 3464 210287
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3528 188873 3556 188974
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 4816 150346 4844 220798
rect 4804 150340 4856 150346
rect 4804 150282 4856 150288
rect 7576 136950 7604 328471
rect 11704 307828 11756 307834
rect 11704 307770 11756 307776
rect 11716 255270 11744 307770
rect 14476 292534 14504 448530
rect 15856 422958 15884 530538
rect 15844 422952 15896 422958
rect 15844 422894 15896 422900
rect 15856 391406 15884 422894
rect 39960 396778 39988 542370
rect 41340 449886 41368 572698
rect 45468 561740 45520 561746
rect 45468 561682 45520 561688
rect 43996 560312 44048 560318
rect 43996 560254 44048 560260
rect 44008 511290 44036 560254
rect 44088 536104 44140 536110
rect 44088 536046 44140 536052
rect 43996 511284 44048 511290
rect 43996 511226 44048 511232
rect 41328 449880 41380 449886
rect 41328 449822 41380 449828
rect 40684 429140 40736 429146
rect 40684 429082 40736 429088
rect 39948 396772 40000 396778
rect 39948 396714 40000 396720
rect 15844 391400 15896 391406
rect 15844 391342 15896 391348
rect 36544 382288 36596 382294
rect 36544 382230 36596 382236
rect 36556 358766 36584 382230
rect 36544 358760 36596 358766
rect 36544 358702 36596 358708
rect 17222 330440 17278 330449
rect 17222 330375 17278 330384
rect 14464 292528 14516 292534
rect 14464 292470 14516 292476
rect 14464 278792 14516 278798
rect 14464 278734 14516 278740
rect 11704 255264 11756 255270
rect 11704 255206 11756 255212
rect 3516 136944 3568 136950
rect 3516 136886 3568 136892
rect 7564 136944 7616 136950
rect 7564 136886 7616 136892
rect 3528 136785 3556 136886
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 14476 85542 14504 278734
rect 17236 97986 17264 330375
rect 36544 328500 36596 328506
rect 36544 328442 36596 328448
rect 33784 327208 33836 327214
rect 33784 327150 33836 327156
rect 29644 319456 29696 319462
rect 29644 319398 29696 319404
rect 22744 307080 22796 307086
rect 22744 307022 22796 307028
rect 21364 218748 21416 218754
rect 21364 218690 21416 218696
rect 17224 97980 17276 97986
rect 17224 97922 17276 97928
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 14464 85536 14516 85542
rect 14464 85478 14516 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 12346 80744 12402 80753
rect 12346 80679 12402 80688
rect 5446 79520 5502 79529
rect 5446 79455 5502 79464
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 4066 68232 4122 68241
rect 4066 68167 4122 68176
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 3974 28248 4030 28257
rect 3974 28183 4030 28192
rect 110 22672 166 22681
rect 110 22607 166 22616
rect 18 6760 74 6769
rect 18 6695 74 6704
rect 124 490 152 22607
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 1676 13184 1728 13190
rect 1676 13126 1728 13132
rect 400 598 612 626
rect 400 490 428 598
rect 124 462 428 490
rect 584 480 612 598
rect 1688 480 1716 13126
rect 3988 3534 4016 28183
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 2884 480 2912 3470
rect 4080 480 4108 68167
rect 5460 6914 5488 79455
rect 10966 35184 11022 35193
rect 10966 35119 11022 35128
rect 9586 10296 9642 10305
rect 9586 10231 9642 10240
rect 5276 6886 5488 6914
rect 5276 480 5304 6886
rect 9600 3534 9628 10231
rect 10980 3534 11008 35119
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6472 480 6500 3402
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 7668 480 7696 2042
rect 8772 480 8800 3470
rect 9968 480 9996 3470
rect 11164 480 11192 3538
rect 12176 3482 12204 14418
rect 12360 6914 12388 80679
rect 17866 72448 17922 72457
rect 17866 72383 17922 72392
rect 15106 59936 15162 59945
rect 15106 59871 15162 59880
rect 13728 17332 13780 17338
rect 13728 17274 13780 17280
rect 13740 6914 13768 17274
rect 15120 6914 15148 59871
rect 16486 43480 16542 43489
rect 16486 43415 16542 43424
rect 12268 6886 12388 6914
rect 13556 6886 13768 6914
rect 14752 6886 15148 6914
rect 12268 3602 12296 6886
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12176 3454 12388 3482
rect 12360 480 12388 3454
rect 13556 480 13584 6886
rect 14752 480 14780 6886
rect 16500 3534 16528 43415
rect 17880 3534 17908 72383
rect 21376 45558 21404 218690
rect 22756 71738 22784 307022
rect 25502 293992 25558 294001
rect 25502 293927 25558 293936
rect 25516 164218 25544 293927
rect 29656 261526 29684 319398
rect 29644 261520 29696 261526
rect 29644 261462 29696 261468
rect 25504 164212 25556 164218
rect 25504 164154 25556 164160
rect 29642 79384 29698 79393
rect 29642 79319 29698 79328
rect 26146 76528 26202 76537
rect 26146 76463 26202 76472
rect 22744 71732 22796 71738
rect 22744 71674 22796 71680
rect 23386 69592 23442 69601
rect 23386 69527 23442 69536
rect 22006 50280 22062 50289
rect 22006 50215 22062 50224
rect 21364 45552 21416 45558
rect 21364 45494 21416 45500
rect 19248 42084 19300 42090
rect 19248 42026 19300 42032
rect 19260 3534 19288 42026
rect 20628 25628 20680 25634
rect 20628 25570 20680 25576
rect 19432 8968 19484 8974
rect 19432 8910 19484 8916
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 16488 3528 16540 3534
rect 16488 3470 16540 3476
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 15948 480 15976 3470
rect 17052 480 17080 3470
rect 18248 480 18276 3470
rect 19444 480 19472 8910
rect 20640 480 20668 25570
rect 22020 6914 22048 50215
rect 23400 6914 23428 69527
rect 24766 29608 24822 29617
rect 24766 29543 24822 29552
rect 21836 6886 22048 6914
rect 23032 6886 23428 6914
rect 21836 480 21864 6886
rect 23032 480 23060 6886
rect 24780 3534 24808 29543
rect 26160 3534 26188 76463
rect 27528 15904 27580 15910
rect 27528 15846 27580 15852
rect 27540 3534 27568 15846
rect 27712 3596 27764 3602
rect 27712 3538 27764 3544
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 26148 3528 26200 3534
rect 26148 3470 26200 3476
rect 26516 3528 26568 3534
rect 26516 3470 26568 3476
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 24228 480 24256 3470
rect 25332 480 25360 3470
rect 26528 480 26556 3470
rect 27724 480 27752 3538
rect 29656 3466 29684 79319
rect 33046 62792 33102 62801
rect 33046 62727 33102 62736
rect 30288 37936 30340 37942
rect 30288 37878 30340 37884
rect 30300 6914 30328 37878
rect 31668 21412 31720 21418
rect 31668 21354 31720 21360
rect 31680 6914 31708 21354
rect 30116 6886 30328 6914
rect 31312 6886 31708 6914
rect 29644 3460 29696 3466
rect 29644 3402 29696 3408
rect 28908 2168 28960 2174
rect 28908 2110 28960 2116
rect 28920 480 28948 2110
rect 30116 480 30144 6886
rect 31312 480 31340 6886
rect 33060 3534 33088 62727
rect 33796 59362 33824 327150
rect 35164 314696 35216 314702
rect 35164 314638 35216 314644
rect 35176 189038 35204 314638
rect 36556 241466 36584 328442
rect 39948 282940 40000 282946
rect 39948 282882 40000 282888
rect 38660 267776 38712 267782
rect 38660 267718 38712 267724
rect 38672 267646 38700 267718
rect 38660 267640 38712 267646
rect 38660 267582 38712 267588
rect 38672 267034 38700 267582
rect 38660 267028 38712 267034
rect 38660 266970 38712 266976
rect 36544 241460 36596 241466
rect 36544 241402 36596 241408
rect 36542 203688 36598 203697
rect 36542 203623 36598 203632
rect 35164 189032 35216 189038
rect 35164 188974 35216 188980
rect 35806 66872 35862 66881
rect 35806 66807 35862 66816
rect 33784 59356 33836 59362
rect 33784 59298 33836 59304
rect 34426 47560 34482 47569
rect 34426 47495 34482 47504
rect 34440 3534 34468 47495
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 32416 480 32444 3470
rect 33612 480 33640 3470
rect 35820 3466 35848 66807
rect 36556 33114 36584 203623
rect 38568 49020 38620 49026
rect 38568 48962 38620 48968
rect 37186 44840 37242 44849
rect 37186 44775 37242 44784
rect 36544 33108 36596 33114
rect 36544 33050 36596 33056
rect 37096 31068 37148 31074
rect 37096 31010 37148 31016
rect 37108 16574 37136 31010
rect 37016 16546 37136 16574
rect 35992 3596 36044 3602
rect 35992 3538 36044 3544
rect 34796 3460 34848 3466
rect 34796 3402 34848 3408
rect 35808 3460 35860 3466
rect 35808 3402 35860 3408
rect 34808 480 34836 3402
rect 36004 480 36032 3538
rect 37016 3482 37044 16546
rect 37200 6914 37228 44775
rect 38580 6914 38608 48962
rect 39960 11762 39988 282882
rect 40696 267782 40724 429082
rect 44008 427145 44036 511226
rect 43994 427136 44050 427145
rect 43994 427071 44050 427080
rect 44100 379506 44128 536046
rect 45480 429146 45508 561682
rect 48148 449206 48176 582354
rect 49608 571396 49660 571402
rect 49608 571338 49660 571344
rect 48228 557592 48280 557598
rect 48228 557534 48280 557540
rect 48136 449200 48188 449206
rect 48136 449142 48188 449148
rect 48136 430636 48188 430642
rect 48136 430578 48188 430584
rect 45468 429140 45520 429146
rect 45468 429082 45520 429088
rect 44088 379500 44140 379506
rect 44088 379442 44140 379448
rect 44088 329860 44140 329866
rect 44088 329802 44140 329808
rect 43444 329112 43496 329118
rect 43444 329054 43496 329060
rect 43456 306338 43484 329054
rect 43444 306332 43496 306338
rect 43444 306274 43496 306280
rect 40684 267776 40736 267782
rect 40684 267718 40736 267724
rect 43444 267640 43496 267646
rect 43444 267582 43496 267588
rect 41328 264988 41380 264994
rect 41328 264930 41380 264936
rect 41340 75177 41368 264930
rect 43456 241466 43484 267582
rect 43444 241460 43496 241466
rect 43444 241402 43496 241408
rect 41326 75168 41382 75177
rect 41326 75103 41382 75112
rect 41326 73808 41382 73817
rect 41326 73743 41382 73752
rect 40682 64152 40738 64161
rect 40682 64087 40738 64096
rect 39948 11756 40000 11762
rect 39948 11698 40000 11704
rect 40696 6914 40724 64087
rect 37108 6886 37228 6914
rect 38396 6886 38608 6914
rect 40604 6886 40724 6914
rect 37108 3602 37136 6886
rect 37096 3596 37148 3602
rect 37096 3538 37148 3544
rect 37016 3454 37228 3482
rect 37200 480 37228 3454
rect 38396 480 38424 6886
rect 39578 6216 39634 6225
rect 39578 6151 39634 6160
rect 39592 480 39620 6151
rect 40604 2106 40632 6886
rect 41340 3466 41368 73743
rect 43996 35216 44048 35222
rect 43996 35158 44048 35164
rect 41880 7608 41932 7614
rect 41880 7550 41932 7556
rect 40684 3460 40736 3466
rect 40684 3402 40736 3408
rect 41328 3460 41380 3466
rect 41328 3402 41380 3408
rect 40592 2100 40644 2106
rect 40592 2042 40644 2048
rect 40696 480 40724 3402
rect 41892 480 41920 7550
rect 44008 3466 44036 35158
rect 44100 17270 44128 329802
rect 46848 318096 46900 318102
rect 46848 318038 46900 318044
rect 46860 317490 46888 318038
rect 46848 317484 46900 317490
rect 46848 317426 46900 317432
rect 46860 197334 46888 317426
rect 48044 292596 48096 292602
rect 48044 292538 48096 292544
rect 48056 231674 48084 292538
rect 48148 235890 48176 430578
rect 48240 421598 48268 557534
rect 49620 453354 49648 571338
rect 50896 564392 50948 564398
rect 50896 564334 50948 564340
rect 49608 453348 49660 453354
rect 49608 453290 49660 453296
rect 49516 449948 49568 449954
rect 49516 449890 49568 449896
rect 48228 421592 48280 421598
rect 48228 421534 48280 421540
rect 49528 329118 49556 449890
rect 50908 431934 50936 564334
rect 51000 457502 51028 585142
rect 51080 576156 51132 576162
rect 51080 576098 51132 576104
rect 51092 575550 51120 576098
rect 51080 575544 51132 575550
rect 51080 575486 51132 575492
rect 52276 575544 52328 575550
rect 52276 575486 52328 575492
rect 50988 457496 51040 457502
rect 50988 457438 51040 457444
rect 52288 447914 52316 575486
rect 53656 566500 53708 566506
rect 53656 566442 53708 566448
rect 52368 545080 52420 545086
rect 52368 545022 52420 545028
rect 52276 447908 52328 447914
rect 52276 447850 52328 447856
rect 50988 445800 51040 445806
rect 50988 445742 51040 445748
rect 50896 431928 50948 431934
rect 50896 431870 50948 431876
rect 50908 430642 50936 431870
rect 50896 430636 50948 430642
rect 50896 430578 50948 430584
rect 50896 401600 50948 401606
rect 50896 401542 50948 401548
rect 49608 331288 49660 331294
rect 49608 331230 49660 331236
rect 49516 329112 49568 329118
rect 49516 329054 49568 329060
rect 48228 270564 48280 270570
rect 48228 270506 48280 270512
rect 48136 235884 48188 235890
rect 48136 235826 48188 235832
rect 48044 231668 48096 231674
rect 48044 231610 48096 231616
rect 46848 197328 46900 197334
rect 46848 197270 46900 197276
rect 47584 53100 47636 53106
rect 47584 53042 47636 53048
rect 45376 46232 45428 46238
rect 45376 46174 45428 46180
rect 44088 17264 44140 17270
rect 44088 17206 44140 17212
rect 45388 3466 45416 46174
rect 46846 26888 46902 26897
rect 46846 26823 46902 26832
rect 46860 6914 46888 26823
rect 46676 6886 46888 6914
rect 45468 4820 45520 4826
rect 45468 4762 45520 4768
rect 43076 3460 43128 3466
rect 43076 3402 43128 3408
rect 43996 3460 44048 3466
rect 43996 3402 44048 3408
rect 44272 3460 44324 3466
rect 44272 3402 44324 3408
rect 45376 3460 45428 3466
rect 45376 3402 45428 3408
rect 43088 480 43116 3402
rect 44284 480 44312 3402
rect 45480 480 45508 4762
rect 46676 480 46704 6886
rect 47596 3534 47624 53042
rect 48240 18630 48268 270506
rect 49620 84862 49648 331230
rect 50804 308440 50856 308446
rect 50804 308382 50856 308388
rect 50816 307834 50844 308382
rect 50804 307828 50856 307834
rect 50804 307770 50856 307776
rect 50816 198694 50844 307770
rect 50908 240145 50936 401542
rect 51000 264246 51028 445742
rect 52274 440872 52330 440881
rect 52274 440807 52330 440816
rect 52288 355366 52316 440807
rect 52380 398886 52408 545022
rect 53472 458856 53524 458862
rect 53472 458798 53524 458804
rect 52368 398880 52420 398886
rect 52368 398822 52420 398828
rect 53484 387705 53512 458798
rect 53668 436082 53696 566442
rect 53760 564398 53788 702510
rect 55036 574796 55088 574802
rect 55036 574738 55088 574744
rect 53748 564392 53800 564398
rect 53748 564334 53800 564340
rect 53748 547188 53800 547194
rect 53748 547130 53800 547136
rect 53656 436076 53708 436082
rect 53656 436018 53708 436024
rect 53760 402974 53788 547130
rect 55048 454714 55076 574738
rect 56508 558952 56560 558958
rect 56508 558894 56560 558900
rect 55128 539640 55180 539646
rect 55128 539582 55180 539588
rect 55036 454708 55088 454714
rect 55036 454650 55088 454656
rect 55034 444680 55090 444689
rect 55034 444615 55090 444624
rect 54942 411360 54998 411369
rect 54942 411295 54998 411304
rect 53576 402946 53788 402974
rect 53576 402286 53604 402946
rect 53564 402280 53616 402286
rect 53564 402222 53616 402228
rect 53470 387696 53526 387705
rect 53470 387631 53526 387640
rect 52366 385656 52422 385665
rect 52366 385591 52422 385600
rect 52276 355360 52328 355366
rect 52276 355302 52328 355308
rect 52288 355094 52316 355302
rect 51724 355088 51776 355094
rect 51724 355030 51776 355036
rect 52276 355088 52328 355094
rect 52276 355030 52328 355036
rect 51736 326398 51764 355030
rect 51724 326392 51776 326398
rect 51724 326334 51776 326340
rect 52184 289128 52236 289134
rect 52184 289070 52236 289076
rect 50988 264240 51040 264246
rect 50988 264182 51040 264188
rect 50988 247104 51040 247110
rect 50988 247046 51040 247052
rect 50894 240136 50950 240145
rect 50894 240071 50950 240080
rect 50804 198688 50856 198694
rect 50804 198630 50856 198636
rect 49608 84856 49660 84862
rect 49608 84798 49660 84804
rect 50894 54496 50950 54505
rect 50894 54431 50950 54440
rect 49608 36576 49660 36582
rect 49608 36518 49660 36524
rect 48228 18624 48280 18630
rect 48228 18566 48280 18572
rect 47860 6180 47912 6186
rect 47860 6122 47912 6128
rect 47584 3528 47636 3534
rect 47584 3470 47636 3476
rect 47872 480 47900 6122
rect 49620 3534 49648 36518
rect 50908 3534 50936 54431
rect 51000 32434 51028 247046
rect 51722 224224 51778 224233
rect 51722 224159 51778 224168
rect 50988 32428 51040 32434
rect 50988 32370 51040 32376
rect 51736 20670 51764 224159
rect 52196 208321 52224 289070
rect 52276 281580 52328 281586
rect 52276 281522 52328 281528
rect 52182 208312 52238 208321
rect 52182 208247 52238 208256
rect 52288 187678 52316 281522
rect 52380 262886 52408 385591
rect 52368 262880 52420 262886
rect 52368 262822 52420 262828
rect 52460 261520 52512 261526
rect 52460 261462 52512 261468
rect 52472 260914 52500 261462
rect 52460 260908 52512 260914
rect 52460 260850 52512 260856
rect 53472 260908 53524 260914
rect 53472 260850 53524 260856
rect 53484 232558 53512 260850
rect 53576 245614 53604 402222
rect 53656 398880 53708 398886
rect 53656 398822 53708 398828
rect 53564 245608 53616 245614
rect 53564 245550 53616 245556
rect 53668 238513 53696 398822
rect 54956 331129 54984 411295
rect 53838 331120 53894 331129
rect 53838 331055 53894 331064
rect 54942 331120 54998 331129
rect 54942 331055 54998 331064
rect 53852 330449 53880 331055
rect 53838 330440 53894 330449
rect 53838 330375 53894 330384
rect 54944 321632 54996 321638
rect 54944 321574 54996 321580
rect 54852 277432 54904 277438
rect 54852 277374 54904 277380
rect 53748 258120 53800 258126
rect 53748 258062 53800 258068
rect 53654 238504 53710 238513
rect 53654 238439 53710 238448
rect 53472 232552 53524 232558
rect 53472 232494 53524 232500
rect 52276 187672 52328 187678
rect 52276 187614 52328 187620
rect 53760 72593 53788 258062
rect 54864 237318 54892 277374
rect 54852 237312 54904 237318
rect 54852 237254 54904 237260
rect 54956 213897 54984 321574
rect 55048 252618 55076 444615
rect 55140 392630 55168 539582
rect 56520 534070 56548 558894
rect 57716 545086 57744 702918
rect 59176 586560 59228 586566
rect 59176 586502 59228 586508
rect 57796 567248 57848 567254
rect 57796 567190 57848 567196
rect 57704 545080 57756 545086
rect 57704 545022 57756 545028
rect 56508 534064 56560 534070
rect 56508 534006 56560 534012
rect 56416 464364 56468 464370
rect 56416 464306 56468 464312
rect 55128 392624 55180 392630
rect 55128 392566 55180 392572
rect 56428 385014 56456 464306
rect 56520 425066 56548 534006
rect 57808 437510 57836 567190
rect 58900 554804 58952 554810
rect 58900 554746 58952 554752
rect 57888 545760 57940 545766
rect 57888 545702 57940 545708
rect 57796 437504 57848 437510
rect 57796 437446 57848 437452
rect 57704 436076 57756 436082
rect 57704 436018 57756 436024
rect 57716 434790 57744 436018
rect 57704 434784 57756 434790
rect 57704 434726 57756 434732
rect 56508 425060 56560 425066
rect 56508 425002 56560 425008
rect 57612 404864 57664 404870
rect 57612 404806 57664 404812
rect 57624 401606 57652 404806
rect 57612 401600 57664 401606
rect 57612 401542 57664 401548
rect 56416 385008 56468 385014
rect 56416 384950 56468 384956
rect 57716 374066 57744 434726
rect 57796 414724 57848 414730
rect 57796 414666 57848 414672
rect 57704 374060 57756 374066
rect 57704 374002 57756 374008
rect 56508 324352 56560 324358
rect 56508 324294 56560 324300
rect 56416 299532 56468 299538
rect 56416 299474 56468 299480
rect 55128 285728 55180 285734
rect 55128 285670 55180 285676
rect 55036 252612 55088 252618
rect 55036 252554 55088 252560
rect 54942 213888 54998 213897
rect 54942 213823 54998 213832
rect 53746 72584 53802 72593
rect 53746 72519 53802 72528
rect 53746 55856 53802 55865
rect 53746 55791 53802 55800
rect 53656 39364 53708 39370
rect 53656 39306 53708 39312
rect 51724 20664 51776 20670
rect 51724 20606 51776 20612
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 49608 3528 49660 3534
rect 49608 3470 49660 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50896 3528 50948 3534
rect 50896 3470 50948 3476
rect 48976 480 49004 3470
rect 50172 480 50200 3470
rect 51356 3460 51408 3466
rect 51356 3402 51408 3408
rect 51368 480 51396 3402
rect 53668 3330 53696 39306
rect 52552 3324 52604 3330
rect 52552 3266 52604 3272
rect 53656 3324 53708 3330
rect 53656 3266 53708 3272
rect 52564 480 52592 3266
rect 53760 480 53788 55791
rect 55036 29640 55088 29646
rect 55036 29582 55088 29588
rect 55048 6914 55076 29582
rect 55140 19990 55168 285670
rect 56324 263628 56376 263634
rect 56324 263570 56376 263576
rect 56336 240009 56364 263570
rect 56322 240000 56378 240009
rect 56322 239935 56378 239944
rect 56428 235929 56456 299474
rect 56414 235920 56470 235929
rect 56414 235855 56470 235864
rect 56520 65521 56548 324294
rect 57716 296682 57744 374002
rect 57704 296676 57756 296682
rect 57704 296618 57756 296624
rect 57704 273964 57756 273970
rect 57704 273906 57756 273912
rect 57612 252612 57664 252618
rect 57612 252554 57664 252560
rect 57624 220833 57652 252554
rect 57610 220824 57666 220833
rect 57610 220759 57666 220768
rect 57716 206990 57744 273906
rect 57808 241369 57836 414666
rect 57900 404870 57928 545702
rect 58912 416838 58940 554746
rect 59188 461650 59216 586502
rect 59280 554742 59308 703326
rect 61844 703180 61896 703186
rect 61844 703122 61896 703128
rect 60004 564460 60056 564466
rect 60004 564402 60056 564408
rect 59268 554736 59320 554742
rect 59268 554678 59320 554684
rect 59176 461644 59228 461650
rect 59176 461586 59228 461592
rect 59084 454776 59136 454782
rect 59084 454718 59136 454724
rect 58992 433900 59044 433906
rect 58992 433842 59044 433848
rect 59004 432070 59032 433842
rect 58992 432064 59044 432070
rect 58992 432006 59044 432012
rect 58900 416832 58952 416838
rect 58900 416774 58952 416780
rect 57888 404864 57940 404870
rect 57888 404806 57940 404812
rect 57980 403640 58032 403646
rect 57980 403582 58032 403588
rect 57992 402286 58020 403582
rect 57980 402280 58032 402286
rect 57980 402222 58032 402228
rect 59004 377369 59032 432006
rect 59096 389298 59124 454718
rect 59174 445904 59230 445913
rect 59174 445839 59230 445848
rect 59084 389292 59136 389298
rect 59084 389234 59136 389240
rect 58990 377360 59046 377369
rect 58990 377295 59046 377304
rect 59188 354674 59216 445839
rect 60016 433906 60044 564402
rect 61856 547806 61884 703122
rect 66168 702500 66220 702506
rect 66168 702442 66220 702448
rect 61934 590744 61990 590753
rect 61934 590679 61990 590688
rect 61844 547800 61896 547806
rect 61844 547742 61896 547748
rect 61856 547194 61884 547742
rect 61844 547188 61896 547194
rect 61844 547130 61896 547136
rect 60556 456136 60608 456142
rect 60556 456078 60608 456084
rect 60004 433900 60056 433906
rect 60004 433842 60056 433848
rect 60568 386374 60596 456078
rect 61948 456074 61976 590679
rect 63316 587920 63368 587926
rect 63316 587862 63368 587868
rect 62028 547936 62080 547942
rect 62028 547878 62080 547884
rect 61936 456068 61988 456074
rect 61936 456010 61988 456016
rect 61936 451988 61988 451994
rect 61936 451930 61988 451936
rect 60648 437504 60700 437510
rect 60648 437446 60700 437452
rect 60556 386368 60608 386374
rect 60556 386310 60608 386316
rect 59096 354646 59216 354674
rect 59096 352073 59124 354646
rect 60660 353977 60688 437446
rect 61842 427136 61898 427145
rect 61842 427071 61898 427080
rect 61856 426426 61884 427071
rect 61844 426420 61896 426426
rect 61844 426362 61896 426368
rect 61856 423858 61884 426362
rect 61764 423830 61884 423858
rect 61764 380186 61792 423830
rect 61844 421592 61896 421598
rect 61844 421534 61896 421540
rect 61752 380180 61804 380186
rect 61752 380122 61804 380128
rect 61856 364334 61884 421534
rect 61948 366353 61976 451930
rect 62040 405822 62068 547878
rect 63328 465118 63356 587862
rect 64696 581052 64748 581058
rect 64696 580994 64748 581000
rect 63408 549296 63460 549302
rect 63408 549238 63460 549244
rect 63316 465112 63368 465118
rect 63316 465054 63368 465060
rect 63328 451274 63356 465054
rect 63236 451246 63356 451274
rect 62028 405816 62080 405822
rect 62028 405758 62080 405764
rect 63236 378826 63264 451246
rect 63316 416832 63368 416838
rect 63316 416774 63368 416780
rect 63224 378820 63276 378826
rect 63224 378762 63276 378768
rect 62028 368552 62080 368558
rect 62028 368494 62080 368500
rect 61934 366344 61990 366353
rect 61934 366279 61990 366288
rect 61856 364306 61976 364334
rect 60646 353968 60702 353977
rect 60646 353903 60702 353912
rect 61948 353326 61976 364306
rect 61936 353320 61988 353326
rect 61936 353262 61988 353268
rect 59082 352064 59138 352073
rect 59082 351999 59138 352008
rect 57888 303680 57940 303686
rect 57888 303622 57940 303628
rect 57794 241360 57850 241369
rect 57794 241295 57850 241304
rect 57704 206984 57756 206990
rect 57704 206926 57756 206932
rect 56506 65512 56562 65521
rect 56506 65447 56562 65456
rect 57900 57225 57928 303622
rect 59096 293962 59124 351999
rect 60462 335472 60518 335481
rect 60462 335407 60518 335416
rect 59176 325712 59228 325718
rect 59176 325654 59228 325660
rect 59084 293956 59136 293962
rect 59084 293898 59136 293904
rect 59084 280220 59136 280226
rect 59084 280162 59136 280168
rect 58992 252136 59044 252142
rect 58992 252078 59044 252084
rect 59004 231849 59032 252078
rect 58990 231840 59046 231849
rect 58990 231775 59046 231784
rect 59096 212537 59124 280162
rect 59188 234569 59216 325654
rect 59268 322992 59320 322998
rect 59268 322934 59320 322940
rect 59174 234560 59230 234569
rect 59174 234495 59230 234504
rect 59082 212528 59138 212537
rect 59082 212463 59138 212472
rect 59176 127016 59228 127022
rect 59176 126958 59228 126964
rect 59188 91798 59216 126958
rect 59176 91792 59228 91798
rect 59176 91734 59228 91740
rect 57886 57216 57942 57225
rect 57886 57151 57942 57160
rect 57886 51776 57942 51785
rect 57886 51711 57942 51720
rect 56508 42152 56560 42158
rect 56508 42094 56560 42100
rect 55128 19984 55180 19990
rect 55128 19926 55180 19932
rect 54956 6886 55076 6914
rect 54956 480 54984 6886
rect 56520 3534 56548 42094
rect 57900 3534 57928 51711
rect 59176 33788 59228 33794
rect 59176 33730 59228 33736
rect 59188 3534 59216 33730
rect 59280 24177 59308 322934
rect 60476 303618 60504 335407
rect 60556 327752 60608 327758
rect 60556 327694 60608 327700
rect 60464 303612 60516 303618
rect 60464 303554 60516 303560
rect 60568 289406 60596 327694
rect 60648 317552 60700 317558
rect 60648 317494 60700 317500
rect 60556 289400 60608 289406
rect 60556 289342 60608 289348
rect 60464 278792 60516 278798
rect 60464 278734 60516 278740
rect 60372 255740 60424 255746
rect 60372 255682 60424 255688
rect 60384 234598 60412 255682
rect 60476 242049 60504 278734
rect 60556 259480 60608 259486
rect 60556 259422 60608 259428
rect 60462 242040 60518 242049
rect 60462 241975 60518 241984
rect 60372 234592 60424 234598
rect 60372 234534 60424 234540
rect 60568 216617 60596 259422
rect 60554 216608 60610 216617
rect 60554 216543 60610 216552
rect 60660 36650 60688 317494
rect 61844 313336 61896 313342
rect 61844 313278 61896 313284
rect 61752 274712 61804 274718
rect 61752 274654 61804 274660
rect 61764 238066 61792 274654
rect 61752 238060 61804 238066
rect 61752 238002 61804 238008
rect 61856 226273 61884 313278
rect 61948 313274 61976 353262
rect 61936 313268 61988 313274
rect 61936 313210 61988 313216
rect 62040 292534 62068 368494
rect 63224 309188 63276 309194
rect 63224 309130 63276 309136
rect 62028 292528 62080 292534
rect 62028 292470 62080 292476
rect 62028 273284 62080 273290
rect 62028 273226 62080 273232
rect 61936 248464 61988 248470
rect 61936 248406 61988 248412
rect 61842 226264 61898 226273
rect 61842 226199 61898 226208
rect 61948 71097 61976 248406
rect 61934 71088 61990 71097
rect 61934 71023 61990 71032
rect 62040 40730 62068 273226
rect 63132 253972 63184 253978
rect 63132 253914 63184 253920
rect 63144 194546 63172 253914
rect 63236 227050 63264 309130
rect 63328 289950 63356 416774
rect 63420 408474 63448 549238
rect 64708 460222 64736 580994
rect 66074 579728 66130 579737
rect 66074 579663 66130 579672
rect 64788 568608 64840 568614
rect 64788 568550 64840 568556
rect 64696 460216 64748 460222
rect 64696 460158 64748 460164
rect 64696 458924 64748 458930
rect 64696 458866 64748 458872
rect 64512 446412 64564 446418
rect 64512 446354 64564 446360
rect 63408 408468 63460 408474
rect 63408 408410 63460 408416
rect 64524 387802 64552 446354
rect 64604 405816 64656 405822
rect 64604 405758 64656 405764
rect 64512 387796 64564 387802
rect 64512 387738 64564 387744
rect 64616 370530 64644 405758
rect 64708 389162 64736 458866
rect 64800 439142 64828 568550
rect 65524 554736 65576 554742
rect 65524 554678 65576 554684
rect 64788 439136 64840 439142
rect 64788 439078 64840 439084
rect 65536 415206 65564 554678
rect 66088 532030 66116 579663
rect 66180 546417 66208 702442
rect 67456 599616 67508 599622
rect 67456 599558 67508 599564
rect 66810 588296 66866 588305
rect 66810 588231 66866 588240
rect 66824 587926 66852 588231
rect 66812 587920 66864 587926
rect 66812 587862 66864 587868
rect 66260 586560 66312 586566
rect 66258 586528 66260 586537
rect 66312 586528 66314 586537
rect 66258 586463 66314 586472
rect 66810 582448 66866 582457
rect 66810 582383 66812 582392
rect 66864 582383 66866 582392
rect 66812 582354 66864 582360
rect 66994 581088 67050 581097
rect 66994 581023 66996 581032
rect 67048 581023 67050 581032
rect 66996 580994 67048 581000
rect 66902 575648 66958 575657
rect 66902 575583 66958 575592
rect 66916 575550 66944 575583
rect 66904 575544 66956 575550
rect 66904 575486 66956 575492
rect 67468 575385 67496 599558
rect 67548 596828 67600 596834
rect 67548 596770 67600 596776
rect 67454 575376 67510 575385
rect 67454 575311 67510 575320
rect 67468 574802 67496 575311
rect 67456 574796 67508 574802
rect 67456 574738 67508 574744
rect 66442 573200 66498 573209
rect 66442 573135 66498 573144
rect 66456 572762 66484 573135
rect 66444 572756 66496 572762
rect 66444 572698 66496 572704
rect 66442 571840 66498 571849
rect 66442 571775 66498 571784
rect 66456 571402 66484 571775
rect 66444 571396 66496 571402
rect 66444 571338 66496 571344
rect 67270 570208 67326 570217
rect 67270 570143 67326 570152
rect 66810 568848 66866 568857
rect 66810 568783 66866 568792
rect 66824 568614 66852 568783
rect 66812 568608 66864 568614
rect 66812 568550 66864 568556
rect 66902 567488 66958 567497
rect 66902 567423 66958 567432
rect 66916 567254 66944 567423
rect 66904 567248 66956 567254
rect 66904 567190 66956 567196
rect 66626 564632 66682 564641
rect 66626 564567 66682 564576
rect 66640 564466 66668 564567
rect 66628 564460 66680 564466
rect 66628 564402 66680 564408
rect 66444 564392 66496 564398
rect 66444 564334 66496 564340
rect 66456 564097 66484 564334
rect 66442 564088 66498 564097
rect 66442 564023 66498 564032
rect 66442 562048 66498 562057
rect 66442 561983 66498 561992
rect 66456 561746 66484 561983
rect 66444 561740 66496 561746
rect 66444 561682 66496 561688
rect 66626 560416 66682 560425
rect 66626 560351 66682 560360
rect 66640 560318 66668 560351
rect 66628 560312 66680 560318
rect 66628 560254 66680 560260
rect 66626 559056 66682 559065
rect 66626 558991 66682 559000
rect 66640 558958 66668 558991
rect 66628 558952 66680 558958
rect 66628 558894 66680 558900
rect 66350 555248 66406 555257
rect 66350 555183 66406 555192
rect 66364 554810 66392 555183
rect 66352 554804 66404 554810
rect 66352 554746 66404 554752
rect 66260 554736 66312 554742
rect 66258 554704 66260 554713
rect 66312 554704 66314 554713
rect 66258 554639 66314 554648
rect 66534 549672 66590 549681
rect 66534 549607 66590 549616
rect 66548 549302 66576 549607
rect 66536 549296 66588 549302
rect 66536 549238 66588 549244
rect 66534 548312 66590 548321
rect 66534 548247 66590 548256
rect 66548 547942 66576 548247
rect 66536 547936 66588 547942
rect 66536 547878 66588 547884
rect 66812 547800 66864 547806
rect 66812 547742 66864 547748
rect 66824 547641 66852 547742
rect 66810 547632 66866 547641
rect 66810 547567 66866 547576
rect 66166 546408 66222 546417
rect 66166 546343 66222 546352
rect 66180 545766 66208 546343
rect 66168 545760 66220 545766
rect 66168 545702 66220 545708
rect 66812 545080 66864 545086
rect 66812 545022 66864 545028
rect 66824 544921 66852 545022
rect 66810 544912 66866 544921
rect 66810 544847 66866 544856
rect 66810 542736 66866 542745
rect 66810 542671 66866 542680
rect 66824 542434 66852 542671
rect 66812 542428 66864 542434
rect 66812 542370 66864 542376
rect 67086 541784 67142 541793
rect 67086 541719 67142 541728
rect 67100 541686 67128 541719
rect 67088 541680 67140 541686
rect 67088 541622 67140 541628
rect 67100 539510 67128 541622
rect 67088 539504 67140 539510
rect 67088 539446 67140 539452
rect 66168 536172 66220 536178
rect 66168 536114 66220 536120
rect 66076 532024 66128 532030
rect 66076 531966 66128 531972
rect 66076 445052 66128 445058
rect 66076 444994 66128 445000
rect 65524 415200 65576 415206
rect 65524 415142 65576 415148
rect 65536 414730 65564 415142
rect 65524 414724 65576 414730
rect 65524 414666 65576 414672
rect 65984 408468 66036 408474
rect 65984 408410 66036 408416
rect 65536 392630 65564 392661
rect 65524 392624 65576 392630
rect 65522 392592 65524 392601
rect 65576 392592 65578 392601
rect 65522 392527 65578 392536
rect 64696 389156 64748 389162
rect 64696 389098 64748 389104
rect 64604 370524 64656 370530
rect 64604 370466 64656 370472
rect 64142 345672 64198 345681
rect 64142 345607 64198 345616
rect 63408 336864 63460 336870
rect 63408 336806 63460 336812
rect 63420 311846 63448 336806
rect 64156 321638 64184 345607
rect 64604 340196 64656 340202
rect 64604 340138 64656 340144
rect 64144 321632 64196 321638
rect 64144 321574 64196 321580
rect 64420 318844 64472 318850
rect 64420 318786 64472 318792
rect 63408 311840 63460 311846
rect 63408 311782 63460 311788
rect 63316 289944 63368 289950
rect 63316 289886 63368 289892
rect 63328 228410 63356 289886
rect 63408 285796 63460 285802
rect 63408 285738 63460 285744
rect 63316 228404 63368 228410
rect 63316 228346 63368 228352
rect 63224 227044 63276 227050
rect 63224 226986 63276 226992
rect 63132 194540 63184 194546
rect 63132 194482 63184 194488
rect 62028 40724 62080 40730
rect 62028 40666 62080 40672
rect 62028 38004 62080 38010
rect 62028 37946 62080 37952
rect 60648 36644 60700 36650
rect 60648 36586 60700 36592
rect 59266 24168 59322 24177
rect 59266 24103 59322 24112
rect 61936 15972 61988 15978
rect 61936 15914 61988 15920
rect 60648 13116 60700 13122
rect 60648 13058 60700 13064
rect 60660 3534 60688 13058
rect 56048 3528 56100 3534
rect 56048 3470 56100 3476
rect 56508 3528 56560 3534
rect 56508 3470 56560 3476
rect 57244 3528 57296 3534
rect 57244 3470 57296 3476
rect 57888 3528 57940 3534
rect 57888 3470 57940 3476
rect 58440 3528 58492 3534
rect 58440 3470 58492 3476
rect 59176 3528 59228 3534
rect 59176 3470 59228 3476
rect 59636 3528 59688 3534
rect 59636 3470 59688 3476
rect 60648 3528 60700 3534
rect 60648 3470 60700 3476
rect 56060 480 56088 3470
rect 57256 480 57284 3470
rect 58452 480 58480 3470
rect 59648 480 59676 3470
rect 61948 3058 61976 15914
rect 60832 3052 60884 3058
rect 60832 2994 60884 3000
rect 61936 3052 61988 3058
rect 61936 2994 61988 3000
rect 60844 480 60872 2994
rect 62040 480 62068 37946
rect 63420 25566 63448 285738
rect 63500 262880 63552 262886
rect 63500 262822 63552 262828
rect 63512 262274 63540 262822
rect 63500 262268 63552 262274
rect 63500 262210 63552 262216
rect 64432 69737 64460 318786
rect 64616 307766 64644 340138
rect 64694 338328 64750 338337
rect 64694 338263 64750 338272
rect 64604 307760 64656 307766
rect 64604 307702 64656 307708
rect 64708 306338 64736 338263
rect 64786 331800 64842 331809
rect 64786 331735 64842 331744
rect 64800 315722 64828 331735
rect 64788 315716 64840 315722
rect 64788 315658 64840 315664
rect 65536 314265 65564 392527
rect 65996 391105 66024 408410
rect 65982 391096 66038 391105
rect 65982 391031 66038 391040
rect 66088 389094 66116 444994
rect 66180 389201 66208 536114
rect 67284 442950 67312 570143
rect 67560 566817 67588 596770
rect 67546 566808 67602 566817
rect 67546 566743 67602 566752
rect 67560 566506 67588 566743
rect 67548 566500 67600 566506
rect 67548 566442 67600 566448
rect 67652 558929 67680 703462
rect 71044 702840 71096 702846
rect 71044 702782 71096 702788
rect 69020 592680 69072 592686
rect 69020 592622 69072 592628
rect 67732 589960 67784 589966
rect 67732 589902 67784 589908
rect 67744 585857 67772 589902
rect 69032 588962 69060 592622
rect 71056 592034 71084 702782
rect 72988 699825 73016 703520
rect 73068 703316 73120 703322
rect 73068 703258 73120 703264
rect 72974 699816 73030 699825
rect 72974 699751 73030 699760
rect 73080 598934 73108 703258
rect 72988 598906 73108 598934
rect 72424 595468 72476 595474
rect 72424 595410 72476 595416
rect 70872 592006 71084 592034
rect 70872 590753 70900 592006
rect 71688 590776 71740 590782
rect 70858 590744 70914 590753
rect 70308 590708 70360 590714
rect 71688 590718 71740 590724
rect 70858 590679 70914 590688
rect 70308 590650 70360 590656
rect 70320 589098 70348 590650
rect 70104 589070 70348 589098
rect 70872 589098 70900 590679
rect 71700 590034 71728 590718
rect 71688 590028 71740 590034
rect 71688 589970 71740 589976
rect 72436 589098 72464 595410
rect 72988 589393 73016 598906
rect 75840 596174 75868 703598
rect 86776 703588 86828 703594
rect 86776 703530 86828 703536
rect 84108 700324 84160 700330
rect 84108 700266 84160 700272
rect 79324 698964 79376 698970
rect 79324 698906 79376 698912
rect 79336 598942 79364 698906
rect 79324 598936 79376 598942
rect 79324 598878 79376 598884
rect 80060 598936 80112 598942
rect 80060 598878 80112 598884
rect 80072 597582 80100 598878
rect 80060 597576 80112 597582
rect 80060 597518 80112 597524
rect 75748 596146 75868 596174
rect 74172 594856 74224 594862
rect 74172 594798 74224 594804
rect 72974 589384 73030 589393
rect 72974 589319 73030 589328
rect 72988 589274 73016 589319
rect 72988 589246 73062 589274
rect 70872 589070 71208 589098
rect 72128 589070 72464 589098
rect 73034 589084 73062 589246
rect 74184 589098 74212 594798
rect 75748 592034 75776 596146
rect 75828 592136 75880 592142
rect 75828 592078 75880 592084
rect 77942 592104 77998 592113
rect 75656 592006 75776 592034
rect 74448 590708 74500 590714
rect 74448 590650 74500 590656
rect 75000 590708 75052 590714
rect 75000 590650 75052 590656
rect 74460 590034 74488 590650
rect 74448 590028 74500 590034
rect 74448 589970 74500 589976
rect 73968 589070 74212 589098
rect 75012 588962 75040 590650
rect 69032 588934 69520 588962
rect 74888 588934 75040 588962
rect 69492 588674 69520 588934
rect 75656 588713 75684 592006
rect 75840 590714 75868 592078
rect 77942 592039 77998 592048
rect 77022 590744 77078 590753
rect 75828 590708 75880 590714
rect 77022 590679 77078 590688
rect 75828 590650 75880 590656
rect 77036 589098 77064 590679
rect 77956 589098 77984 592039
rect 78404 590844 78456 590850
rect 78404 590786 78456 590792
rect 76728 589070 77064 589098
rect 77648 589070 77984 589098
rect 78416 588826 78444 590786
rect 80072 589098 80100 597518
rect 81346 595504 81402 595513
rect 84120 595474 84148 700266
rect 81346 595439 81402 595448
rect 84108 595468 84160 595474
rect 81360 589274 81388 595439
rect 84108 595410 84160 595416
rect 83464 593496 83516 593502
rect 83464 593438 83516 593444
rect 82542 591016 82598 591025
rect 82542 590951 82598 590960
rect 81438 590744 81494 590753
rect 81438 590679 81494 590688
rect 81452 589286 81480 590679
rect 81314 589246 81388 589274
rect 81440 589280 81492 589286
rect 80072 589070 80408 589098
rect 81314 589084 81342 589246
rect 81440 589222 81492 589228
rect 82556 589098 82584 590951
rect 83476 589098 83504 593438
rect 84108 592068 84160 592074
rect 84108 592010 84160 592016
rect 84120 589274 84148 592010
rect 86788 591002 86816 703530
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 136652 703582 137692 703610
rect 89180 700330 89208 703520
rect 93768 703452 93820 703458
rect 93768 703394 93820 703400
rect 89812 702636 89864 702642
rect 89812 702578 89864 702584
rect 89168 700324 89220 700330
rect 89168 700266 89220 700272
rect 88984 700256 89036 700262
rect 88984 700198 89036 700204
rect 88800 600976 88852 600982
rect 88800 600918 88852 600924
rect 88812 596174 88840 600918
rect 88996 599622 89024 700198
rect 88984 599616 89036 599622
rect 88984 599558 89036 599564
rect 88812 596146 88932 596174
rect 86788 590974 87000 591002
rect 86866 590880 86922 590889
rect 86866 590815 86922 590824
rect 86224 590776 86276 590782
rect 86224 590718 86276 590724
rect 82248 589070 82584 589098
rect 83168 589070 83504 589098
rect 84074 589246 84148 589274
rect 84074 589084 84102 589246
rect 86236 589098 86264 590718
rect 86880 589274 86908 590815
rect 85928 589070 86264 589098
rect 86834 589246 86908 589274
rect 86834 589084 86862 589246
rect 78416 588798 78568 588826
rect 75642 588704 75698 588713
rect 69480 588668 69532 588674
rect 75642 588639 75698 588648
rect 69480 588610 69532 588616
rect 75656 588554 75684 588639
rect 86972 588606 87000 590974
rect 88800 590708 88852 590714
rect 88800 590650 88852 590656
rect 88248 589280 88300 589286
rect 88248 589222 88300 589228
rect 88260 588849 88288 589222
rect 88812 589098 88840 590650
rect 88688 589070 88840 589098
rect 88246 588840 88302 588849
rect 88246 588775 88302 588784
rect 85304 588600 85356 588606
rect 75656 588526 75808 588554
rect 79488 588526 79824 588554
rect 85008 588548 85304 588554
rect 85008 588542 85356 588548
rect 86960 588600 87012 588606
rect 88062 588568 88118 588577
rect 86960 588542 87012 588548
rect 85008 588526 85344 588542
rect 87768 588526 88062 588554
rect 79796 588470 79824 588526
rect 88062 588503 88118 588512
rect 79784 588464 79836 588470
rect 79784 588406 79836 588412
rect 67730 585848 67786 585857
rect 67730 585783 67786 585792
rect 67744 585206 67772 585783
rect 67732 585200 67784 585206
rect 67732 585142 67784 585148
rect 67730 578368 67786 578377
rect 67730 578303 67786 578312
rect 67638 558920 67694 558929
rect 67638 558855 67694 558864
rect 67652 557598 67680 558855
rect 67640 557592 67692 557598
rect 67640 557534 67692 557540
rect 67362 556336 67418 556345
rect 67362 556271 67418 556280
rect 67272 442944 67324 442950
rect 67272 442886 67324 442892
rect 66994 439920 67050 439929
rect 66994 439855 67050 439864
rect 67008 439142 67036 439855
rect 66996 439136 67048 439142
rect 66996 439078 67048 439084
rect 67272 439136 67324 439142
rect 67272 439078 67324 439084
rect 66810 437744 66866 437753
rect 66810 437679 66866 437688
rect 66824 437510 66852 437679
rect 66812 437504 66864 437510
rect 66812 437446 66864 437452
rect 66810 435296 66866 435305
rect 66810 435231 66866 435240
rect 66824 434790 66852 435231
rect 66812 434784 66864 434790
rect 66812 434726 66864 434732
rect 66902 433120 66958 433129
rect 66902 433055 66958 433064
rect 66916 432070 66944 433055
rect 66904 432064 66956 432070
rect 66904 432006 66956 432012
rect 66904 431928 66956 431934
rect 66904 431870 66956 431876
rect 66916 430953 66944 431870
rect 66902 430944 66958 430953
rect 66902 430879 66958 430888
rect 66812 429140 66864 429146
rect 66812 429082 66864 429088
rect 66824 428505 66852 429082
rect 66810 428496 66866 428505
rect 66810 428431 66866 428440
rect 66260 426420 66312 426426
rect 66260 426362 66312 426368
rect 66272 426329 66300 426362
rect 66258 426320 66314 426329
rect 66258 426255 66314 426264
rect 66260 425060 66312 425066
rect 66260 425002 66312 425008
rect 66272 424153 66300 425002
rect 66258 424144 66314 424153
rect 66258 424079 66314 424088
rect 66258 421968 66314 421977
rect 66258 421903 66314 421912
rect 66272 421598 66300 421903
rect 66260 421592 66312 421598
rect 66260 421534 66312 421540
rect 66902 417344 66958 417353
rect 66902 417279 66958 417288
rect 66916 416838 66944 417279
rect 66904 416832 66956 416838
rect 66904 416774 66956 416780
rect 66444 415200 66496 415206
rect 66442 415168 66444 415177
rect 66496 415168 66498 415177
rect 66442 415103 66498 415112
rect 66536 408468 66588 408474
rect 66536 408410 66588 408416
rect 66548 408377 66576 408410
rect 66534 408368 66590 408377
rect 66534 408303 66590 408312
rect 66626 406192 66682 406201
rect 66626 406127 66682 406136
rect 66640 405822 66668 406127
rect 66628 405816 66680 405822
rect 66628 405758 66680 405764
rect 66350 403744 66406 403753
rect 66350 403679 66406 403688
rect 66364 403646 66392 403679
rect 66352 403640 66404 403646
rect 66352 403582 66404 403588
rect 66812 401600 66864 401606
rect 66810 401568 66812 401577
rect 66864 401568 66866 401577
rect 66810 401503 66866 401512
rect 66902 399392 66958 399401
rect 66902 399327 66958 399336
rect 66916 398886 66944 399327
rect 66904 398880 66956 398886
rect 66904 398822 66956 398828
rect 66258 396944 66314 396953
rect 66258 396879 66314 396888
rect 66272 396778 66300 396879
rect 66260 396772 66312 396778
rect 66260 396714 66312 396720
rect 66166 389192 66222 389201
rect 66166 389127 66222 389136
rect 66076 389088 66128 389094
rect 66076 389030 66128 389036
rect 66166 356688 66222 356697
rect 66166 356623 66222 356632
rect 66076 336048 66128 336054
rect 66076 335990 66128 335996
rect 65984 334620 66036 334626
rect 65984 334562 66036 334568
rect 65522 314256 65578 314265
rect 65522 314191 65578 314200
rect 65536 313342 65564 314191
rect 65524 313336 65576 313342
rect 65524 313278 65576 313284
rect 64696 306332 64748 306338
rect 64696 306274 64748 306280
rect 65996 301481 66024 334562
rect 65982 301472 66038 301481
rect 65982 301407 66038 301416
rect 64696 287088 64748 287094
rect 64696 287030 64748 287036
rect 64512 269136 64564 269142
rect 64512 269078 64564 269084
rect 64524 241505 64552 269078
rect 64604 262268 64656 262274
rect 64604 262210 64656 262216
rect 64510 241496 64566 241505
rect 64510 241431 64566 241440
rect 64616 232665 64644 262210
rect 64602 232656 64658 232665
rect 64602 232591 64658 232600
rect 64708 213926 64736 287030
rect 66088 276049 66116 335990
rect 66074 276040 66130 276049
rect 66074 275975 66130 275984
rect 66074 272096 66130 272105
rect 66074 272031 66130 272040
rect 65984 264240 66036 264246
rect 65984 264182 66036 264188
rect 65890 250064 65946 250073
rect 65890 249999 65946 250008
rect 65904 237590 65932 249999
rect 65892 237584 65944 237590
rect 65892 237526 65944 237532
rect 65996 235958 66024 264182
rect 65984 235952 66036 235958
rect 65984 235894 66036 235900
rect 66088 227662 66116 272031
rect 66180 267730 66208 356623
rect 67284 341193 67312 439078
rect 67376 419529 67404 556271
rect 67454 552256 67510 552265
rect 67454 552191 67510 552200
rect 67362 419520 67418 419529
rect 67362 419455 67418 419464
rect 67468 412729 67496 552191
rect 67548 540932 67600 540938
rect 67548 540874 67600 540880
rect 67560 539646 67588 540874
rect 67548 539640 67600 539646
rect 67548 539582 67600 539588
rect 67548 539504 67600 539510
rect 67548 539446 67600 539452
rect 67454 412720 67510 412729
rect 67454 412655 67510 412664
rect 67362 396944 67418 396953
rect 67362 396879 67418 396888
rect 67376 349081 67404 396879
rect 67362 349072 67418 349081
rect 67362 349007 67418 349016
rect 67270 341184 67326 341193
rect 67270 341119 67326 341128
rect 67180 335368 67232 335374
rect 67180 335310 67232 335316
rect 66812 326868 66864 326874
rect 66812 326810 66864 326816
rect 66718 323776 66774 323785
rect 66718 323711 66774 323720
rect 66732 322998 66760 323711
rect 66720 322992 66772 322998
rect 66720 322934 66772 322940
rect 66628 321564 66680 321570
rect 66628 321506 66680 321512
rect 66640 320521 66668 321506
rect 66626 320512 66682 320521
rect 66626 320447 66682 320456
rect 66718 318336 66774 318345
rect 66718 318271 66774 318280
rect 66732 317490 66760 318271
rect 66720 317484 66772 317490
rect 66720 317426 66772 317432
rect 66626 309904 66682 309913
rect 66626 309839 66682 309848
rect 66640 309194 66668 309839
rect 66628 309188 66680 309194
rect 66628 309130 66680 309136
rect 66536 307760 66588 307766
rect 66536 307702 66588 307708
rect 66548 306921 66576 307702
rect 66534 306912 66590 306921
rect 66534 306847 66590 306856
rect 66718 293040 66774 293049
rect 66718 292975 66774 292984
rect 66732 292602 66760 292975
rect 66720 292596 66772 292602
rect 66720 292538 66772 292544
rect 66718 287872 66774 287881
rect 66718 287807 66774 287816
rect 66732 287094 66760 287807
rect 66720 287088 66772 287094
rect 66720 287030 66772 287036
rect 66824 287054 66852 326810
rect 66902 324864 66958 324873
rect 66902 324799 66958 324808
rect 66916 324358 66944 324799
rect 66904 324352 66956 324358
rect 66904 324294 66956 324300
rect 67192 322697 67220 335310
rect 67284 327049 67312 341119
rect 67364 332648 67416 332654
rect 67364 332590 67416 332596
rect 67270 327040 67326 327049
rect 67270 326975 67326 326984
rect 67178 322688 67234 322697
rect 67178 322623 67234 322632
rect 66902 319424 66958 319433
rect 66902 319359 66958 319368
rect 66916 318850 66944 319359
rect 66904 318844 66956 318850
rect 66904 318786 66956 318792
rect 66904 317552 66956 317558
rect 66902 317520 66904 317529
rect 66956 317520 66958 317529
rect 66902 317455 66958 317464
rect 66996 315716 67048 315722
rect 66996 315658 67048 315664
rect 66904 313268 66956 313274
rect 66904 313210 66956 313216
rect 66916 313177 66944 313210
rect 66902 313168 66958 313177
rect 66902 313103 66958 313112
rect 66904 311840 66956 311846
rect 66904 311782 66956 311788
rect 66916 311001 66944 311782
rect 66902 310992 66958 311001
rect 66902 310927 66958 310936
rect 67008 306374 67036 315658
rect 67086 309088 67142 309097
rect 67086 309023 67142 309032
rect 67100 308446 67128 309023
rect 67088 308440 67140 308446
rect 67088 308382 67140 308388
rect 67086 308000 67142 308009
rect 67086 307935 67142 307944
rect 67100 307086 67128 307935
rect 67088 307080 67140 307086
rect 67088 307022 67140 307028
rect 67008 306346 67128 306374
rect 66904 306332 66956 306338
rect 66904 306274 66956 306280
rect 66916 305833 66944 306274
rect 66902 305824 66958 305833
rect 66902 305759 66958 305768
rect 66904 303680 66956 303686
rect 66902 303648 66904 303657
rect 66956 303648 66958 303657
rect 66902 303583 66958 303592
rect 66996 303612 67048 303618
rect 66996 303554 67048 303560
rect 67008 302569 67036 303554
rect 66994 302560 67050 302569
rect 66994 302495 67050 302504
rect 66902 300656 66958 300665
rect 66902 300591 66958 300600
rect 66916 299538 66944 300591
rect 67100 299577 67128 306346
rect 67178 304736 67234 304745
rect 67178 304671 67234 304680
rect 67086 299568 67142 299577
rect 66904 299532 66956 299538
rect 67086 299503 67142 299512
rect 66904 299474 66956 299480
rect 66904 296676 66956 296682
rect 66904 296618 66956 296624
rect 66916 296313 66944 296618
rect 66902 296304 66958 296313
rect 66902 296239 66958 296248
rect 67086 294128 67142 294137
rect 67086 294063 67142 294072
rect 66996 293956 67048 293962
rect 66996 293898 67048 293904
rect 66904 292528 66956 292534
rect 66904 292470 66956 292476
rect 66916 292233 66944 292470
rect 66902 292224 66958 292233
rect 66902 292159 66958 292168
rect 67008 291145 67036 293898
rect 66994 291136 67050 291145
rect 66994 291071 67050 291080
rect 66902 290048 66958 290057
rect 66902 289983 66958 289992
rect 66916 289950 66944 289983
rect 66904 289944 66956 289950
rect 66904 289886 66956 289892
rect 66904 289400 66956 289406
rect 66904 289342 66956 289348
rect 66916 288969 66944 289342
rect 66902 288960 66958 288969
rect 66902 288895 66958 288904
rect 66824 287026 67036 287054
rect 66902 286784 66958 286793
rect 66902 286719 66958 286728
rect 66916 285802 66944 286719
rect 66904 285796 66956 285802
rect 66904 285738 66956 285744
rect 66812 285728 66864 285734
rect 66810 285696 66812 285705
rect 66864 285696 66866 285705
rect 66810 285631 66866 285640
rect 67008 284617 67036 287026
rect 66994 284608 67050 284617
rect 66994 284543 67050 284552
rect 66718 283792 66774 283801
rect 66718 283727 66774 283736
rect 66732 282946 66760 283727
rect 66720 282940 66772 282946
rect 66720 282882 66772 282888
rect 66350 282704 66406 282713
rect 66350 282639 66406 282648
rect 66364 281586 66392 282639
rect 66352 281580 66404 281586
rect 66352 281522 66404 281528
rect 66810 280528 66866 280537
rect 66810 280463 66866 280472
rect 66824 280226 66852 280463
rect 66812 280220 66864 280226
rect 66812 280162 66864 280168
rect 66718 278352 66774 278361
rect 66718 278287 66774 278296
rect 66732 277438 66760 278287
rect 66720 277432 66772 277438
rect 67100 277394 67128 294063
rect 67192 289134 67220 304671
rect 67376 298489 67404 332590
rect 67468 309097 67496 412655
rect 67560 394777 67588 539446
rect 67744 467838 67772 578303
rect 67822 577008 67878 577017
rect 67822 576943 67878 576952
rect 67836 539034 67864 576943
rect 88904 576813 88932 596146
rect 89076 590844 89128 590850
rect 89076 590786 89128 590792
rect 88984 588668 89036 588674
rect 88984 588610 89036 588616
rect 88890 576804 88946 576813
rect 88890 576739 88946 576748
rect 88904 575550 88932 576739
rect 88892 575544 88944 575550
rect 88892 575486 88944 575492
rect 68652 540932 68704 540938
rect 68652 540874 68704 540880
rect 68664 540841 68692 540874
rect 68650 540832 68706 540841
rect 68650 540767 68706 540776
rect 69848 539640 69900 539646
rect 69848 539582 69900 539588
rect 76746 539608 76802 539617
rect 69860 539458 69888 539582
rect 76802 539566 77096 539594
rect 76746 539543 76802 539552
rect 69736 539444 69888 539458
rect 69722 539430 69888 539444
rect 68480 539158 68816 539186
rect 67824 539028 67876 539034
rect 67824 538970 67876 538976
rect 68480 535537 68508 539158
rect 69722 539050 69750 539430
rect 70656 539158 70716 539186
rect 69676 539022 69750 539050
rect 69676 535537 69704 539022
rect 70688 538218 70716 539158
rect 71240 539158 71576 539186
rect 72436 539158 72496 539186
rect 73172 539158 73416 539186
rect 74000 539158 74336 539186
rect 74552 539158 75256 539186
rect 76176 539158 76236 539186
rect 70676 538212 70728 538218
rect 70676 538154 70728 538160
rect 70688 535537 70716 538154
rect 68466 535528 68522 535537
rect 68466 535463 68522 535472
rect 69662 535528 69718 535537
rect 69662 535463 69718 535472
rect 70674 535528 70730 535537
rect 70674 535463 70730 535472
rect 71240 528554 71268 539158
rect 72436 537538 72464 539158
rect 72424 537532 72476 537538
rect 72424 537474 72476 537480
rect 70504 528526 71268 528554
rect 67732 467832 67784 467838
rect 67732 467774 67784 467780
rect 70504 458930 70532 528526
rect 70492 458924 70544 458930
rect 70492 458866 70544 458872
rect 69662 458280 69718 458289
rect 69662 458215 69718 458224
rect 67640 453348 67692 453354
rect 67640 453290 67692 453296
rect 67652 444650 67680 453290
rect 69676 449886 69704 458215
rect 72056 454708 72108 454714
rect 72056 454650 72108 454656
rect 72068 452742 72096 454650
rect 72056 452736 72108 452742
rect 72056 452678 72108 452684
rect 69664 449880 69716 449886
rect 69664 449822 69716 449828
rect 68284 447840 68336 447846
rect 68284 447782 68336 447788
rect 68296 447234 68324 447782
rect 68284 447228 68336 447234
rect 68284 447170 68336 447176
rect 68560 447228 68612 447234
rect 68560 447170 68612 447176
rect 67640 444644 67692 444650
rect 67640 444586 67692 444592
rect 67824 444644 67876 444650
rect 67824 444586 67876 444592
rect 67732 442944 67784 442950
rect 67732 442886 67784 442892
rect 67744 442105 67772 442886
rect 67730 442096 67786 442105
rect 67730 442031 67786 442040
rect 67546 394768 67602 394777
rect 67546 394703 67602 394712
rect 67560 332654 67588 394703
rect 67640 380248 67692 380254
rect 67640 380190 67692 380196
rect 67548 332648 67600 332654
rect 67548 332590 67600 332596
rect 67546 315344 67602 315353
rect 67546 315279 67602 315288
rect 67560 314702 67588 315279
rect 67548 314696 67600 314702
rect 67548 314638 67600 314644
rect 67454 309088 67510 309097
rect 67454 309023 67510 309032
rect 67362 298480 67418 298489
rect 67362 298415 67418 298424
rect 67180 289128 67232 289134
rect 67180 289070 67232 289076
rect 67546 281616 67602 281625
rect 67546 281551 67602 281560
rect 67270 279440 67326 279449
rect 67270 279375 67326 279384
rect 67284 278798 67312 279375
rect 67272 278792 67324 278798
rect 67272 278734 67324 278740
rect 66720 277374 66772 277380
rect 66916 277366 67128 277394
rect 66810 275360 66866 275369
rect 66810 275295 66866 275304
rect 66824 274718 66852 275295
rect 66812 274712 66864 274718
rect 66812 274654 66864 274660
rect 66810 274272 66866 274281
rect 66810 274207 66866 274216
rect 66824 273290 66852 274207
rect 66916 273970 66944 277366
rect 67086 277264 67142 277273
rect 67086 277199 67142 277208
rect 66904 273964 66956 273970
rect 66904 273906 66956 273912
rect 66812 273284 66864 273290
rect 66812 273226 66864 273232
rect 66994 273184 67050 273193
rect 66994 273119 67050 273128
rect 66902 271008 66958 271017
rect 66902 270943 66958 270952
rect 66916 270570 66944 270943
rect 66904 270564 66956 270570
rect 66904 270506 66956 270512
rect 67008 270450 67036 273119
rect 66916 270422 67036 270450
rect 66718 269920 66774 269929
rect 66718 269855 66774 269864
rect 66732 269142 66760 269855
rect 66720 269136 66772 269142
rect 66720 269078 66772 269084
rect 66258 267744 66314 267753
rect 66180 267702 66258 267730
rect 66180 228313 66208 267702
rect 66258 267679 66314 267688
rect 66810 265840 66866 265849
rect 66810 265775 66866 265784
rect 66824 264994 66852 265775
rect 66812 264988 66864 264994
rect 66812 264930 66864 264936
rect 66810 264752 66866 264761
rect 66810 264687 66866 264696
rect 66536 264240 66588 264246
rect 66536 264182 66588 264188
rect 66548 263673 66576 264182
rect 66534 263664 66590 263673
rect 66824 263634 66852 264687
rect 66534 263599 66590 263608
rect 66812 263628 66864 263634
rect 66812 263570 66864 263576
rect 66442 262576 66498 262585
rect 66442 262511 66498 262520
rect 66456 262274 66484 262511
rect 66444 262268 66496 262274
rect 66444 262210 66496 262216
rect 66810 261488 66866 261497
rect 66810 261423 66866 261432
rect 66824 260914 66852 261423
rect 66812 260908 66864 260914
rect 66812 260850 66864 260856
rect 66810 260400 66866 260409
rect 66810 260335 66866 260344
rect 66824 259486 66852 260335
rect 66812 259480 66864 259486
rect 66812 259422 66864 259428
rect 66718 258496 66774 258505
rect 66718 258431 66774 258440
rect 66732 258126 66760 258431
rect 66720 258120 66772 258126
rect 66916 258074 66944 270422
rect 67100 258074 67128 277199
rect 66720 258062 66772 258068
rect 66824 258046 66944 258074
rect 67008 258046 67128 258074
rect 67456 258052 67508 258058
rect 66824 252142 66852 258046
rect 67008 255746 67036 258046
rect 67456 257994 67508 258000
rect 66996 255740 67048 255746
rect 66996 255682 67048 255688
rect 66902 254144 66958 254153
rect 66902 254079 66958 254088
rect 66916 253978 66944 254079
rect 66904 253972 66956 253978
rect 66904 253914 66956 253920
rect 66902 253056 66958 253065
rect 66902 252991 66958 253000
rect 66916 252618 66944 252991
rect 66904 252612 66956 252618
rect 66904 252554 66956 252560
rect 66812 252136 66864 252142
rect 66812 252078 66864 252084
rect 66810 248976 66866 248985
rect 66810 248911 66866 248920
rect 66824 248470 66852 248911
rect 66812 248464 66864 248470
rect 67468 248414 67496 257994
rect 66812 248406 66864 248412
rect 67376 248386 67496 248414
rect 66626 247888 66682 247897
rect 66626 247823 66682 247832
rect 66640 247110 66668 247823
rect 66628 247104 66680 247110
rect 66628 247046 66680 247052
rect 67270 246800 67326 246809
rect 67270 246735 67326 246744
rect 66628 245608 66680 245614
rect 66628 245550 66680 245556
rect 66640 245177 66668 245550
rect 66626 245168 66682 245177
rect 66626 245103 66682 245112
rect 67178 242856 67234 242865
rect 67178 242791 67234 242800
rect 66166 228304 66222 228313
rect 66166 228239 66222 228248
rect 66076 227656 66128 227662
rect 66076 227598 66128 227604
rect 67192 217297 67220 242791
rect 67284 222873 67312 246735
rect 67376 239873 67404 248386
rect 67456 248328 67508 248334
rect 67456 248270 67508 248276
rect 67468 242078 67496 248270
rect 67456 242072 67508 242078
rect 67456 242014 67508 242020
rect 67560 240786 67588 281551
rect 67652 268841 67680 380190
rect 67744 374678 67772 442031
rect 67836 376038 67864 444586
rect 68572 441614 68600 447170
rect 68790 444644 68842 444650
rect 68790 444586 68842 444592
rect 68802 444380 68830 444586
rect 69676 444394 69704 449822
rect 72068 444394 72096 452678
rect 72436 445058 72464 537474
rect 73172 536110 73200 539158
rect 73160 536104 73212 536110
rect 73160 536046 73212 536052
rect 74000 535498 74028 539158
rect 73160 535492 73212 535498
rect 73160 535434 73212 535440
rect 73988 535492 74040 535498
rect 73988 535434 74040 535440
rect 73172 454782 73200 535434
rect 73160 454776 73212 454782
rect 73160 454718 73212 454724
rect 73344 447908 73396 447914
rect 73344 447850 73396 447856
rect 72424 445052 72476 445058
rect 72424 444994 72476 445000
rect 73356 444514 73384 447850
rect 74552 446418 74580 539158
rect 74632 539028 74684 539034
rect 74632 538970 74684 538976
rect 74644 449954 74672 538970
rect 76208 536761 76236 539158
rect 76194 536752 76250 536761
rect 76194 536687 76250 536696
rect 76208 536178 76236 536687
rect 76196 536172 76248 536178
rect 76196 536114 76248 536120
rect 76760 535537 76788 539543
rect 77312 539158 78016 539186
rect 78876 539158 78936 539186
rect 79520 539158 79856 539186
rect 80776 539158 81112 539186
rect 76102 535528 76158 535537
rect 76102 535463 76158 535472
rect 76746 535528 76802 535537
rect 76746 535463 76802 535472
rect 76116 456142 76144 535463
rect 76564 467832 76616 467838
rect 76564 467774 76616 467780
rect 76104 456136 76156 456142
rect 76104 456078 76156 456084
rect 74632 449948 74684 449954
rect 74632 449890 74684 449896
rect 74540 446412 74592 446418
rect 74540 446354 74592 446360
rect 73344 444508 73396 444514
rect 73344 444450 73396 444456
rect 73356 444394 73384 444450
rect 69676 444366 70288 444394
rect 71760 444366 72096 444394
rect 73232 444366 73384 444394
rect 74644 444394 74672 449890
rect 76576 446049 76604 467774
rect 77312 458862 77340 539158
rect 78772 535492 78824 535498
rect 78772 535434 78824 535440
rect 77944 532024 77996 532030
rect 77944 531966 77996 531972
rect 77300 458856 77352 458862
rect 77300 458798 77352 458804
rect 77956 448662 77984 531966
rect 78784 464370 78812 535434
rect 78772 464364 78824 464370
rect 78772 464306 78824 464312
rect 78680 460216 78732 460222
rect 78680 460158 78732 460164
rect 77944 448656 77996 448662
rect 77944 448598 77996 448604
rect 76562 446040 76618 446049
rect 76562 445975 76618 445984
rect 76576 444394 76604 445975
rect 77956 444394 77984 448598
rect 78692 446962 78720 460158
rect 78876 451994 78904 539158
rect 79520 535498 79548 539158
rect 81084 538286 81112 539158
rect 81452 539158 81696 539186
rect 82616 539158 82768 539186
rect 83536 539158 84148 539186
rect 84456 539158 84792 539186
rect 85376 539158 85528 539186
rect 86296 539158 86632 539186
rect 81072 538280 81124 538286
rect 81072 538222 81124 538228
rect 79508 535492 79560 535498
rect 79508 535434 79560 535440
rect 81452 462913 81480 539158
rect 82740 536790 82768 539158
rect 82728 536784 82780 536790
rect 82728 536726 82780 536732
rect 81438 462904 81494 462913
rect 81438 462839 81494 462848
rect 82740 453257 82768 536726
rect 83464 457496 83516 457502
rect 83464 457438 83516 457444
rect 82726 453248 82782 453257
rect 82726 453183 82782 453192
rect 82082 452704 82138 452713
rect 82082 452639 82138 452648
rect 78864 451988 78916 451994
rect 78864 451930 78916 451936
rect 80060 449200 80112 449206
rect 80060 449142 80112 449148
rect 80072 448594 80100 449142
rect 80060 448588 80112 448594
rect 80060 448530 80112 448536
rect 80888 448588 80940 448594
rect 80888 448530 80940 448536
rect 78680 446956 78732 446962
rect 78680 446898 78732 446904
rect 79140 446956 79192 446962
rect 79140 446898 79192 446904
rect 79152 445806 79180 446898
rect 79140 445800 79192 445806
rect 79140 445742 79192 445748
rect 74644 444366 74888 444394
rect 76360 444366 76604 444394
rect 77832 444366 77984 444394
rect 79152 444394 79180 445742
rect 80900 444530 80928 448530
rect 80900 444502 80974 444530
rect 79152 444366 79488 444394
rect 80946 444380 80974 444502
rect 82096 444394 82124 452639
rect 83476 451353 83504 457438
rect 84120 454753 84148 539158
rect 84764 536081 84792 539158
rect 85500 536246 85528 539158
rect 86604 538214 86632 539158
rect 86972 539158 87400 539186
rect 88320 539158 88380 539186
rect 86868 538214 86920 538218
rect 86604 538212 86920 538214
rect 86604 538186 86868 538212
rect 86868 538154 86920 538160
rect 85488 536240 85540 536246
rect 85488 536182 85540 536188
rect 86224 536240 86276 536246
rect 86224 536182 86276 536188
rect 84750 536072 84806 536081
rect 84750 536007 84806 536016
rect 85580 461644 85632 461650
rect 85580 461586 85632 461592
rect 84106 454744 84162 454753
rect 84106 454679 84162 454688
rect 83462 451344 83518 451353
rect 83462 451279 83518 451288
rect 83476 444394 83504 451279
rect 85592 445913 85620 461586
rect 86236 447817 86264 536182
rect 86880 457473 86908 538154
rect 86972 458833 87000 539158
rect 87052 465112 87104 465118
rect 87052 465054 87104 465060
rect 86958 458824 87014 458833
rect 86958 458759 87014 458768
rect 86866 457464 86922 457473
rect 86866 457399 86922 457408
rect 86222 447808 86278 447817
rect 86222 447743 86278 447752
rect 85578 445904 85634 445913
rect 85578 445839 85634 445848
rect 85592 444666 85620 445839
rect 87064 444666 87092 465054
rect 88352 456113 88380 539158
rect 88338 456104 88394 456113
rect 88338 456039 88394 456048
rect 88996 451274 89024 588610
rect 89088 585818 89116 590786
rect 89720 590028 89772 590034
rect 89720 589970 89772 589976
rect 89076 585812 89128 585818
rect 89076 585754 89128 585760
rect 88904 451246 89024 451274
rect 88904 445777 88932 451246
rect 88890 445768 88946 445777
rect 88890 445703 88946 445712
rect 85546 444638 85620 444666
rect 87018 444638 87092 444666
rect 82096 444366 82432 444394
rect 83476 444366 83904 444394
rect 85546 444380 85574 444638
rect 87018 444380 87046 444638
rect 88904 444394 88932 445703
rect 88504 444366 88932 444394
rect 89732 444394 89760 589970
rect 89824 560153 89852 702578
rect 91100 598256 91152 598262
rect 91100 598198 91152 598204
rect 90364 593428 90416 593434
rect 90364 593370 90416 593376
rect 90376 590782 90404 593370
rect 90364 590776 90416 590782
rect 90364 590718 90416 590724
rect 90376 585721 90404 590718
rect 89902 585712 89958 585721
rect 89902 585647 89958 585656
rect 90362 585712 90418 585721
rect 90362 585647 90418 585656
rect 89810 560144 89866 560153
rect 89810 560079 89866 560088
rect 89916 538898 89944 585647
rect 91112 573594 91140 598198
rect 92480 595468 92532 595474
rect 92480 595410 92532 595416
rect 91190 587072 91246 587081
rect 91190 587007 91246 587016
rect 91204 586566 91232 587007
rect 91192 586560 91244 586566
rect 91192 586502 91244 586508
rect 92110 584896 92166 584905
rect 92110 584831 92166 584840
rect 92124 584458 92152 584831
rect 92112 584452 92164 584458
rect 92112 584394 92164 584400
rect 91928 583704 91980 583710
rect 91926 583672 91928 583681
rect 91980 583672 91982 583681
rect 91926 583607 91982 583616
rect 91190 581632 91246 581641
rect 91190 581567 91246 581576
rect 91204 581058 91232 581567
rect 91192 581052 91244 581058
rect 91192 580994 91244 581000
rect 91190 578912 91246 578921
rect 91190 578847 91246 578856
rect 91204 578270 91232 578847
rect 91192 578264 91244 578270
rect 91192 578206 91244 578212
rect 91190 577552 91246 577561
rect 91190 577487 91246 577496
rect 91204 576910 91232 577487
rect 91192 576904 91244 576910
rect 91192 576846 91244 576852
rect 91926 574832 91982 574841
rect 91926 574767 91928 574776
rect 91980 574767 91982 574776
rect 91928 574738 91980 574744
rect 91112 573566 91324 573594
rect 91098 573472 91154 573481
rect 91098 573407 91154 573416
rect 91112 572762 91140 573407
rect 91100 572756 91152 572762
rect 91100 572698 91152 572704
rect 91190 572112 91246 572121
rect 91190 572047 91246 572056
rect 91100 571464 91152 571470
rect 91098 571432 91100 571441
rect 91152 571432 91154 571441
rect 91204 571402 91232 572047
rect 91098 571367 91154 571376
rect 91192 571396 91244 571402
rect 91192 571338 91244 571344
rect 91098 570072 91154 570081
rect 91098 570007 91154 570016
rect 91112 569974 91140 570007
rect 91100 569968 91152 569974
rect 91100 569910 91152 569916
rect 91296 567866 91324 573566
rect 91742 568712 91798 568721
rect 91742 568647 91798 568656
rect 91100 567860 91152 567866
rect 91100 567802 91152 567808
rect 91284 567860 91336 567866
rect 91284 567802 91336 567808
rect 91112 567769 91140 567802
rect 91098 567760 91154 567769
rect 91098 567695 91154 567704
rect 91100 565888 91152 565894
rect 91098 565856 91100 565865
rect 91152 565856 91154 565865
rect 91098 565791 91154 565800
rect 91098 564496 91154 564505
rect 91098 564431 91100 564440
rect 91152 564431 91154 564440
rect 91100 564402 91152 564408
rect 91098 563136 91154 563145
rect 91098 563071 91100 563080
rect 91152 563071 91154 563080
rect 91100 563042 91152 563048
rect 91098 560960 91154 560969
rect 91098 560895 91154 560904
rect 89904 538892 89956 538898
rect 89904 538834 89956 538840
rect 91112 530602 91140 560895
rect 91190 558240 91246 558249
rect 91190 558175 91246 558184
rect 91204 557598 91232 558175
rect 91192 557592 91244 557598
rect 91192 557534 91244 557540
rect 91190 556880 91246 556889
rect 91190 556815 91246 556824
rect 91204 556238 91232 556815
rect 91192 556232 91244 556238
rect 91192 556174 91244 556180
rect 91190 555520 91246 555529
rect 91190 555455 91246 555464
rect 91204 554810 91232 555455
rect 91192 554804 91244 554810
rect 91192 554746 91244 554752
rect 91282 552800 91338 552809
rect 91282 552735 91338 552744
rect 91192 552152 91244 552158
rect 91190 552120 91192 552129
rect 91244 552120 91246 552129
rect 91296 552090 91324 552735
rect 91190 552055 91246 552064
rect 91284 552084 91336 552090
rect 91284 552026 91336 552032
rect 91190 549400 91246 549409
rect 91190 549335 91246 549344
rect 91204 549302 91232 549335
rect 91192 549296 91244 549302
rect 91192 549238 91244 549244
rect 91190 547904 91246 547913
rect 91190 547839 91246 547848
rect 91204 533390 91232 547839
rect 91282 546544 91338 546553
rect 91282 546479 91284 546488
rect 91336 546479 91338 546488
rect 91284 546450 91336 546456
rect 91296 544490 91324 546450
rect 91296 544462 91416 544490
rect 91284 544400 91336 544406
rect 91284 544342 91336 544348
rect 91296 544105 91324 544342
rect 91282 544096 91338 544105
rect 91282 544031 91338 544040
rect 91282 542464 91338 542473
rect 91282 542399 91284 542408
rect 91336 542399 91338 542408
rect 91284 542370 91336 542376
rect 91284 541680 91336 541686
rect 91284 541622 91336 541628
rect 91296 541385 91324 541622
rect 91282 541376 91338 541385
rect 91282 541311 91338 541320
rect 91282 539744 91338 539753
rect 91282 539679 91284 539688
rect 91336 539679 91338 539688
rect 91284 539650 91336 539656
rect 91388 534750 91416 544462
rect 91376 534744 91428 534750
rect 91376 534686 91428 534692
rect 91192 533384 91244 533390
rect 91192 533326 91244 533332
rect 91100 530596 91152 530602
rect 91100 530538 91152 530544
rect 91100 456068 91152 456074
rect 91100 456010 91152 456016
rect 91112 454102 91140 456010
rect 91100 454096 91152 454102
rect 91100 454038 91152 454044
rect 91112 451274 91140 454038
rect 91756 453257 91784 568647
rect 91834 560144 91890 560153
rect 91834 560079 91890 560088
rect 91848 548554 91876 560079
rect 91836 548548 91888 548554
rect 91836 548490 91888 548496
rect 91742 453248 91798 453257
rect 91742 453183 91798 453192
rect 91112 451246 91232 451274
rect 90132 444544 90188 444553
rect 90132 444479 90188 444488
rect 90146 444394 90174 444479
rect 89732 444380 90174 444394
rect 91204 444394 91232 451246
rect 92492 444689 92520 595410
rect 93780 584458 93808 703394
rect 101404 703112 101456 703118
rect 101404 703054 101456 703060
rect 97908 702772 97960 702778
rect 97908 702714 97960 702720
rect 94504 702636 94556 702642
rect 94504 702578 94556 702584
rect 93768 584452 93820 584458
rect 93768 584394 93820 584400
rect 94516 583710 94544 702578
rect 95884 594856 95936 594862
rect 95884 594798 95936 594804
rect 93768 583704 93820 583710
rect 93768 583646 93820 583652
rect 94504 583704 94556 583710
rect 94504 583646 94556 583652
rect 93780 581641 93808 583646
rect 93766 581632 93822 581641
rect 93766 581567 93822 581576
rect 93768 574796 93820 574802
rect 93768 574738 93820 574744
rect 93780 569226 93808 574738
rect 93768 569220 93820 569226
rect 93768 569162 93820 569168
rect 92570 545184 92626 545193
rect 92570 545119 92626 545128
rect 92584 543017 92612 545119
rect 92570 543008 92626 543017
rect 92570 542943 92626 542952
rect 94504 542428 94556 542434
rect 94504 542370 94556 542376
rect 93124 539708 93176 539714
rect 93124 539650 93176 539656
rect 93136 464409 93164 539650
rect 93122 464400 93178 464409
rect 93122 464335 93178 464344
rect 94516 462913 94544 542370
rect 94502 462904 94558 462913
rect 94502 462839 94558 462848
rect 95896 449954 95924 594798
rect 96620 592136 96672 592142
rect 96620 592078 96672 592084
rect 96528 544400 96580 544406
rect 96528 544342 96580 544348
rect 96540 465769 96568 544342
rect 96526 465760 96582 465769
rect 96526 465695 96582 465704
rect 95884 449948 95936 449954
rect 95884 449890 95936 449896
rect 94410 445768 94466 445777
rect 94410 445703 94466 445712
rect 92478 444680 92534 444689
rect 92478 444615 92534 444624
rect 93076 444680 93132 444689
rect 93076 444615 93132 444624
rect 89732 444366 90160 444380
rect 91204 444366 91632 444394
rect 93090 444380 93118 444615
rect 94424 444394 94452 445703
rect 95896 444394 95924 449890
rect 96632 445777 96660 592078
rect 97920 580961 97948 702714
rect 97998 592104 98054 592113
rect 97998 592039 98054 592048
rect 97906 580952 97962 580961
rect 97906 580887 97962 580896
rect 97920 580281 97948 580887
rect 97906 580272 97962 580281
rect 97906 580207 97962 580216
rect 97264 571464 97316 571470
rect 97264 571406 97316 571412
rect 97276 456074 97304 571406
rect 97264 456068 97316 456074
rect 97264 456010 97316 456016
rect 98012 445806 98040 592039
rect 100022 590880 100078 590889
rect 100022 590815 100078 590824
rect 98642 588704 98698 588713
rect 98642 588639 98698 588648
rect 98656 447166 98684 588639
rect 100036 551342 100064 590815
rect 100758 588840 100814 588849
rect 100758 588775 100814 588784
rect 100024 551336 100076 551342
rect 100024 551278 100076 551284
rect 100772 460934 100800 588775
rect 101416 574802 101444 703054
rect 105464 700330 105492 703520
rect 130384 703248 130436 703254
rect 130384 703190 130436 703196
rect 124864 703044 124916 703050
rect 124864 702986 124916 702992
rect 105452 700324 105504 700330
rect 105452 700266 105504 700272
rect 106924 597576 106976 597582
rect 106924 597518 106976 597524
rect 105544 587172 105596 587178
rect 105544 587114 105596 587120
rect 103520 585812 103572 585818
rect 103520 585754 103572 585760
rect 102784 581052 102836 581058
rect 102784 580994 102836 581000
rect 101404 574796 101456 574802
rect 101404 574738 101456 574744
rect 101404 565888 101456 565894
rect 101404 565830 101456 565836
rect 100772 460906 100984 460934
rect 98644 447160 98696 447166
rect 98644 447102 98696 447108
rect 98000 445800 98052 445806
rect 96618 445768 96674 445777
rect 96618 445703 96674 445712
rect 97354 445768 97410 445777
rect 97354 445703 97410 445712
rect 97998 445768 98000 445777
rect 98052 445768 98054 445777
rect 97998 445703 98054 445712
rect 97368 444394 97396 445703
rect 98656 444394 98684 447102
rect 100956 444689 100984 460906
rect 101416 456142 101444 565830
rect 102796 458862 102824 580994
rect 102784 458856 102836 458862
rect 102784 458798 102836 458804
rect 101404 456136 101456 456142
rect 101404 456078 101456 456084
rect 103532 447234 103560 585754
rect 104808 577516 104860 577522
rect 104808 577458 104860 577464
rect 104820 576910 104848 577458
rect 104808 576904 104860 576910
rect 104808 576846 104860 576852
rect 104164 546508 104216 546514
rect 104164 546450 104216 546456
rect 104176 462233 104204 546450
rect 104162 462224 104218 462233
rect 104162 462159 104218 462168
rect 104820 447817 104848 576846
rect 104806 447808 104862 447817
rect 104806 447743 104862 447752
rect 103520 447228 103572 447234
rect 103520 447170 103572 447176
rect 102140 445800 102192 445806
rect 102140 445742 102192 445748
rect 100942 444680 100998 444689
rect 100942 444615 100998 444624
rect 100956 444394 100984 444615
rect 94424 444366 94760 444394
rect 95896 444366 96232 444394
rect 97368 444366 97704 444394
rect 98656 444366 99176 444394
rect 100832 444366 100984 444394
rect 102152 444394 102180 445742
rect 103532 444394 103560 447170
rect 105556 445806 105584 587114
rect 105636 575544 105688 575550
rect 105636 575486 105688 575492
rect 105648 457502 105676 575486
rect 105636 457496 105688 457502
rect 105636 457438 105688 457444
rect 106936 445874 106964 597518
rect 108302 595504 108358 595513
rect 108302 595439 108358 595448
rect 107106 591016 107162 591025
rect 107106 590951 107162 590960
rect 107120 553110 107148 590951
rect 107108 553104 107160 553110
rect 107108 553046 107160 553052
rect 107016 552152 107068 552158
rect 107016 552094 107068 552100
rect 107028 462913 107056 552094
rect 108120 545760 108172 545766
rect 108120 545702 108172 545708
rect 108132 543017 108160 545702
rect 108118 543008 108174 543017
rect 108118 542943 108174 542952
rect 107014 462904 107070 462913
rect 107014 462839 107070 462848
rect 108316 448769 108344 595439
rect 110420 593496 110472 593502
rect 110420 593438 110472 593444
rect 108948 554804 109000 554810
rect 108948 554746 109000 554752
rect 108302 448760 108358 448769
rect 108302 448695 108358 448704
rect 106924 445868 106976 445874
rect 106924 445810 106976 445816
rect 105544 445800 105596 445806
rect 105544 445742 105596 445748
rect 105556 444394 105584 445742
rect 106936 444666 106964 445810
rect 102152 444366 102304 444394
rect 103532 444366 103776 444394
rect 105432 444366 105584 444394
rect 106890 444638 106964 444666
rect 108316 444666 108344 448695
rect 108960 447953 108988 554746
rect 109040 553104 109092 553110
rect 109040 553046 109092 553052
rect 108946 447944 109002 447953
rect 108946 447879 109002 447888
rect 108316 444638 108390 444666
rect 106890 444380 106918 444638
rect 108362 444380 108390 444638
rect 109052 444394 109080 553046
rect 110432 445777 110460 593438
rect 112444 592068 112496 592074
rect 112444 592010 112496 592016
rect 111064 549296 111116 549302
rect 111064 549238 111116 549244
rect 111076 448633 111104 549238
rect 112456 452674 112484 592010
rect 113180 588600 113232 588606
rect 113180 588542 113232 588548
rect 112444 452668 112496 452674
rect 112444 452610 112496 452616
rect 112456 451246 112484 452610
rect 112444 451240 112496 451246
rect 112444 451182 112496 451188
rect 111062 448624 111118 448633
rect 111062 448559 111118 448568
rect 110418 445768 110474 445777
rect 110418 445703 110474 445712
rect 111154 445768 111210 445777
rect 111154 445703 111210 445712
rect 109498 444816 109554 444825
rect 109498 444751 109554 444760
rect 109512 444394 109540 444751
rect 111168 444394 111196 445703
rect 112456 444394 112484 451182
rect 113192 445777 113220 588542
rect 116582 585712 116638 585721
rect 116582 585647 116638 585656
rect 115204 584452 115256 584458
rect 115204 584394 115256 584400
rect 115216 447846 115244 584394
rect 115388 539572 115440 539578
rect 115388 539514 115440 539520
rect 115400 538665 115428 539514
rect 115386 538656 115442 538665
rect 115386 538591 115442 538600
rect 115400 538286 115428 538591
rect 115388 538280 115440 538286
rect 115388 538222 115440 538228
rect 116596 450022 116624 585647
rect 121552 578264 121604 578270
rect 121552 578206 121604 578212
rect 120816 572756 120868 572762
rect 120816 572698 120868 572704
rect 120632 564460 120684 564466
rect 120632 564402 120684 564408
rect 117320 551336 117372 551342
rect 117320 551278 117372 551284
rect 116584 450016 116636 450022
rect 116584 449958 116636 449964
rect 115204 447840 115256 447846
rect 115204 447782 115256 447788
rect 113178 445768 113234 445777
rect 113178 445703 113234 445712
rect 114098 445768 114154 445777
rect 114098 445703 114154 445712
rect 114112 444394 114140 445703
rect 116596 444394 116624 449958
rect 117332 445777 117360 551278
rect 118698 460184 118754 460193
rect 118698 460119 118754 460128
rect 117318 445768 117374 445777
rect 117318 445703 117374 445712
rect 109052 444366 109848 444394
rect 111168 444366 111504 444394
rect 112456 444366 112976 444394
rect 114112 444366 114448 444394
rect 116104 444366 116624 444394
rect 117332 444394 117360 445703
rect 118712 444394 118740 460119
rect 119160 444440 119212 444446
rect 117332 444366 117576 444394
rect 118712 444388 119160 444394
rect 118712 444382 119212 444388
rect 118712 444366 119200 444382
rect 68572 441586 68692 441614
rect 68664 389065 68692 441586
rect 120644 404297 120672 564402
rect 120724 451920 120776 451926
rect 120724 451862 120776 451868
rect 120736 440201 120764 451862
rect 120722 440192 120778 440201
rect 120722 440127 120778 440136
rect 120722 434752 120778 434761
rect 120722 434687 120778 434696
rect 120630 404288 120686 404297
rect 120630 404223 120686 404232
rect 120644 403034 120672 404223
rect 120632 403028 120684 403034
rect 120632 402970 120684 402976
rect 86222 390960 86278 390969
rect 86222 390895 86278 390904
rect 92754 390960 92810 390969
rect 102138 390960 102194 390969
rect 92810 390918 93440 390946
rect 92754 390895 92810 390904
rect 70030 390688 70086 390697
rect 70086 390646 70288 390674
rect 73232 390646 73384 390674
rect 70030 390623 70086 390632
rect 68802 390130 68830 390388
rect 68802 390102 68876 390130
rect 68650 389056 68706 389065
rect 68650 388991 68706 389000
rect 68848 388793 68876 390102
rect 68834 388784 68890 388793
rect 68834 388719 68890 388728
rect 70136 386414 70164 390646
rect 71870 390416 71926 390425
rect 71760 390374 71870 390402
rect 71926 390374 72188 390402
rect 71870 390351 71926 390360
rect 71884 390291 71912 390351
rect 70136 386386 70348 386414
rect 67824 376032 67876 376038
rect 67824 375974 67876 375980
rect 67732 374672 67784 374678
rect 67732 374614 67784 374620
rect 70320 371890 70348 386386
rect 72160 383654 72188 390374
rect 73356 389162 73384 390646
rect 80058 390416 80114 390425
rect 74552 390374 74888 390402
rect 75932 390374 76360 390402
rect 77404 390374 77832 390402
rect 79152 390374 79488 390402
rect 73160 389156 73212 389162
rect 73160 389098 73212 389104
rect 73344 389156 73396 389162
rect 73344 389098 73396 389104
rect 72160 383626 72464 383654
rect 70308 371884 70360 371890
rect 70308 371826 70360 371832
rect 71688 365288 71740 365294
rect 71688 365230 71740 365236
rect 71042 355328 71098 355337
rect 71042 355263 71098 355272
rect 70398 351928 70454 351937
rect 70398 351863 70454 351872
rect 67824 351212 67876 351218
rect 67824 351154 67876 351160
rect 67730 347032 67786 347041
rect 67730 346967 67786 346976
rect 67744 312089 67772 346967
rect 67836 321609 67864 351154
rect 70412 345014 70440 351863
rect 70412 344986 70808 345014
rect 70122 342272 70178 342281
rect 70122 342207 70178 342216
rect 69112 329860 69164 329866
rect 69112 329802 69164 329808
rect 68006 328672 68062 328681
rect 68006 328607 68062 328616
rect 68020 326874 68048 328607
rect 69124 327434 69152 329802
rect 70136 327570 70164 342207
rect 70674 332752 70730 332761
rect 70674 332687 70730 332696
rect 70688 327570 70716 332687
rect 69736 327542 70164 327570
rect 70472 327542 70716 327570
rect 69000 327406 69152 327434
rect 70780 327162 70808 344986
rect 70780 327134 70992 327162
rect 70032 327072 70084 327078
rect 70030 327040 70032 327049
rect 70084 327040 70086 327049
rect 70030 326975 70086 326984
rect 68652 326936 68704 326942
rect 68652 326878 68704 326884
rect 70964 326890 70992 327134
rect 71056 327078 71084 355263
rect 71700 351937 71728 365230
rect 71686 351928 71742 351937
rect 71686 351863 71742 351872
rect 72436 340202 72464 383626
rect 73172 365294 73200 389098
rect 74552 389094 74580 390374
rect 74540 389088 74592 389094
rect 74540 389030 74592 389036
rect 73160 365288 73212 365294
rect 73160 365230 73212 365236
rect 74448 345704 74500 345710
rect 74448 345646 74500 345652
rect 72424 340196 72476 340202
rect 72424 340138 72476 340144
rect 73066 339688 73122 339697
rect 73066 339623 73122 339632
rect 71410 334248 71466 334257
rect 71410 334183 71466 334192
rect 71044 327072 71096 327078
rect 71044 327014 71096 327020
rect 71424 326942 71452 334183
rect 72240 330540 72292 330546
rect 72240 330482 72292 330488
rect 72252 327570 72280 330482
rect 73080 327570 73108 339623
rect 74460 335354 74488 345646
rect 74552 336054 74580 389030
rect 75932 379506 75960 390374
rect 77404 389298 77432 390374
rect 77392 389292 77444 389298
rect 77392 389234 77444 389240
rect 75920 379500 75972 379506
rect 75920 379442 75972 379448
rect 76564 379500 76616 379506
rect 76564 379442 76616 379448
rect 76576 362273 76604 379442
rect 77404 373994 77432 389234
rect 79152 387802 79180 390374
rect 80058 390351 80114 390360
rect 80610 390416 80666 390425
rect 80666 390374 80960 390402
rect 82096 390374 82432 390402
rect 83568 390374 83904 390402
rect 80610 390351 80666 390360
rect 80072 389201 80100 390351
rect 80058 389192 80114 389201
rect 80058 389127 80114 389136
rect 79140 387796 79192 387802
rect 79140 387738 79192 387744
rect 79152 387326 79180 387738
rect 78680 387320 78732 387326
rect 78680 387262 78732 387268
rect 79140 387320 79192 387326
rect 79140 387262 79192 387268
rect 77312 373966 77432 373994
rect 76562 362264 76618 362273
rect 76562 362199 76618 362208
rect 77312 358057 77340 373966
rect 77298 358048 77354 358057
rect 77298 357983 77354 357992
rect 78692 347070 78720 387262
rect 80072 364993 80100 389127
rect 82096 386374 82124 390374
rect 83568 387705 83596 390374
rect 85546 390130 85574 390388
rect 85546 390102 85620 390130
rect 83554 387696 83610 387705
rect 83554 387631 83610 387640
rect 83568 387297 83596 387631
rect 83554 387288 83610 387297
rect 83554 387223 83610 387232
rect 82084 386368 82136 386374
rect 82084 386310 82136 386316
rect 82096 365702 82124 386310
rect 85486 378856 85542 378865
rect 85486 378791 85542 378800
rect 81440 365696 81492 365702
rect 81440 365638 81492 365644
rect 82084 365696 82136 365702
rect 82084 365638 82136 365644
rect 80058 364984 80114 364993
rect 80058 364919 80114 364928
rect 81452 364410 81480 365638
rect 81440 364404 81492 364410
rect 81440 364346 81492 364352
rect 80058 357504 80114 357513
rect 80058 357439 80114 357448
rect 79968 351280 80020 351286
rect 79968 351222 80020 351228
rect 78680 347064 78732 347070
rect 78680 347006 78732 347012
rect 77208 343664 77260 343670
rect 77208 343606 77260 343612
rect 75828 341556 75880 341562
rect 75828 341498 75880 341504
rect 74630 336832 74686 336841
rect 74630 336767 74686 336776
rect 74540 336048 74592 336054
rect 74540 335990 74592 335996
rect 74368 335326 74488 335354
rect 73710 334384 73766 334393
rect 73710 334319 73766 334328
rect 73724 327570 73752 334319
rect 74368 327570 74396 335326
rect 74644 327842 74672 336767
rect 74644 327814 74718 327842
rect 71944 327542 72280 327570
rect 72680 327542 73108 327570
rect 73416 327542 73752 327570
rect 73968 327542 74396 327570
rect 74690 327556 74718 327814
rect 75840 327570 75868 341498
rect 77116 338768 77168 338774
rect 77116 338710 77168 338716
rect 77128 331158 77156 338710
rect 76472 331152 76524 331158
rect 76472 331094 76524 331100
rect 77116 331152 77168 331158
rect 77116 331094 77168 331100
rect 76484 327570 76512 331094
rect 77220 327570 77248 343606
rect 79876 342916 79928 342922
rect 79876 342858 79928 342864
rect 77300 340264 77352 340270
rect 77300 340206 77352 340212
rect 77312 327593 77340 340206
rect 77942 332616 77998 332625
rect 77942 332551 77998 332560
rect 75440 327542 75868 327570
rect 76176 327542 76512 327570
rect 76912 327542 77248 327570
rect 77298 327584 77354 327593
rect 77956 327570 77984 332551
rect 79416 329996 79468 330002
rect 79416 329938 79468 329944
rect 77648 327542 77984 327570
rect 78218 327584 78274 327593
rect 77298 327519 77354 327528
rect 79428 327570 79456 329938
rect 79888 327570 79916 342858
rect 79980 330002 80008 351222
rect 79968 329996 80020 330002
rect 79968 329938 80020 329944
rect 78274 327556 78384 327570
rect 78274 327542 78398 327556
rect 79120 327542 79456 327570
rect 79672 327542 79916 327570
rect 80072 327570 80100 357439
rect 80702 341048 80758 341057
rect 80702 340983 80758 340992
rect 80716 327570 80744 340983
rect 81452 327570 81480 364346
rect 83464 352572 83516 352578
rect 83464 352514 83516 352520
rect 82726 338736 82782 338745
rect 82726 338671 82782 338680
rect 82740 327570 82768 338671
rect 80072 327542 80408 327570
rect 80716 327542 81144 327570
rect 81452 327542 81880 327570
rect 82616 327542 82768 327570
rect 83002 327584 83058 327593
rect 78218 327519 78274 327528
rect 78370 327298 78398 327542
rect 83476 327570 83504 352514
rect 85500 345098 85528 378791
rect 85592 368626 85620 390102
rect 85580 368620 85632 368626
rect 85580 368562 85632 368568
rect 85592 366353 85620 368562
rect 85578 366344 85634 366353
rect 85578 366279 85634 366288
rect 86236 354674 86264 390895
rect 91374 390416 91430 390425
rect 87018 390130 87046 390388
rect 88352 390374 88504 390402
rect 89824 390374 90160 390402
rect 87018 390102 87092 390130
rect 87064 385014 87092 390102
rect 87052 385008 87104 385014
rect 87052 384950 87104 384956
rect 87064 384402 87092 384950
rect 87052 384396 87104 384402
rect 87052 384338 87104 384344
rect 88248 384396 88300 384402
rect 88248 384338 88300 384344
rect 87604 378820 87656 378826
rect 87604 378762 87656 378768
rect 86960 366376 87012 366382
rect 86960 366318 87012 366324
rect 86972 357513 87000 366318
rect 87616 363089 87644 378762
rect 88260 378729 88288 384338
rect 88352 382226 88380 390374
rect 89824 389065 89852 390374
rect 91430 390374 91968 390402
rect 91374 390351 91430 390360
rect 91940 389162 91968 390374
rect 91928 389156 91980 389162
rect 91928 389098 91980 389104
rect 93216 389156 93268 389162
rect 93216 389098 93268 389104
rect 89810 389056 89866 389065
rect 89810 388991 89866 389000
rect 91006 388376 91062 388385
rect 91006 388311 91062 388320
rect 88340 382220 88392 382226
rect 88340 382162 88392 382168
rect 88246 378720 88302 378729
rect 88246 378655 88302 378664
rect 87602 363080 87658 363089
rect 87602 363015 87658 363024
rect 86958 357504 87014 357513
rect 86958 357439 87014 357448
rect 85776 354646 86264 354674
rect 85776 349353 85804 354646
rect 85762 349344 85818 349353
rect 85762 349279 85818 349288
rect 84200 345092 84252 345098
rect 84200 345034 84252 345040
rect 85488 345092 85540 345098
rect 85488 345034 85540 345040
rect 84212 335354 84240 345034
rect 85776 345014 85804 349279
rect 85776 344986 86448 345014
rect 85672 338156 85724 338162
rect 85672 338098 85724 338104
rect 84212 335326 84424 335354
rect 83740 331288 83792 331294
rect 83740 331230 83792 331236
rect 83058 327542 83504 327570
rect 83752 327570 83780 331230
rect 84396 327570 84424 335326
rect 85684 327570 85712 338098
rect 86316 331900 86368 331906
rect 86316 331842 86368 331848
rect 86328 327570 86356 331842
rect 83752 327542 84088 327570
rect 84396 327542 84824 327570
rect 85560 327542 85712 327570
rect 86112 327542 86356 327570
rect 86420 327570 86448 344986
rect 87616 338774 87644 363015
rect 88984 358828 89036 358834
rect 88984 358770 89036 358776
rect 88996 342922 89024 358770
rect 91020 347818 91048 388311
rect 93124 387796 93176 387802
rect 93124 387738 93176 387744
rect 91190 359272 91246 359281
rect 91190 359207 91246 359216
rect 91204 358834 91232 359207
rect 91192 358828 91244 358834
rect 91192 358770 91244 358776
rect 92388 356720 92440 356726
rect 92388 356662 92440 356668
rect 89720 347812 89772 347818
rect 89720 347754 89772 347760
rect 91008 347812 91060 347818
rect 91008 347754 91060 347760
rect 89732 345710 89760 347754
rect 89720 345704 89772 345710
rect 89720 345646 89772 345652
rect 90916 343732 90968 343738
rect 90916 343674 90968 343680
rect 88984 342916 89036 342922
rect 88984 342858 89036 342864
rect 87604 338768 87656 338774
rect 87604 338710 87656 338716
rect 87142 337104 87198 337113
rect 87142 337039 87198 337048
rect 87156 327570 87184 337039
rect 88614 336968 88670 336977
rect 88614 336903 88670 336912
rect 88430 330032 88486 330041
rect 88430 329967 88486 329976
rect 86420 327542 86848 327570
rect 87156 327542 87584 327570
rect 83002 327519 83058 327528
rect 88444 327434 88472 329967
rect 88628 327570 88656 336903
rect 89810 335608 89866 335617
rect 89810 335543 89866 335552
rect 89824 327842 89852 335543
rect 89778 327814 89852 327842
rect 88628 327542 89056 327570
rect 89778 327556 89806 327814
rect 90928 327570 90956 343674
rect 92400 335354 92428 356662
rect 93136 340270 93164 387738
rect 93228 354006 93256 389098
rect 93412 388482 93440 390918
rect 107934 390960 107990 390969
rect 102194 390918 102640 390946
rect 102138 390895 102194 390904
rect 94576 390646 94728 390674
rect 93400 388476 93452 388482
rect 93400 388418 93452 388424
rect 94700 387870 94728 390646
rect 95882 390416 95938 390425
rect 97354 390416 97410 390425
rect 95938 390374 96232 390402
rect 95882 390351 95938 390360
rect 98826 390416 98882 390425
rect 97410 390374 97856 390402
rect 97354 390351 97410 390360
rect 95238 388512 95294 388521
rect 95238 388447 95294 388456
rect 94688 387864 94740 387870
rect 94688 387806 94740 387812
rect 95252 366382 95280 388447
rect 95896 387025 95924 390351
rect 95882 387016 95938 387025
rect 95882 386951 95938 386960
rect 97262 369880 97318 369889
rect 97262 369815 97318 369824
rect 95240 366376 95292 366382
rect 95240 366318 95292 366324
rect 96526 361040 96582 361049
rect 96526 360975 96582 360984
rect 95146 356280 95202 356289
rect 95146 356215 95202 356224
rect 95160 355366 95188 356215
rect 93860 355360 93912 355366
rect 93860 355302 93912 355308
rect 95148 355360 95200 355366
rect 95148 355302 95200 355308
rect 93216 354000 93268 354006
rect 93216 353942 93268 353948
rect 93676 342304 93728 342310
rect 93676 342246 93728 342252
rect 93124 340264 93176 340270
rect 93124 340206 93176 340212
rect 92216 335326 92428 335354
rect 91100 329860 91152 329866
rect 91100 329802 91152 329808
rect 91112 327758 91140 329802
rect 91100 327752 91152 327758
rect 91100 327694 91152 327700
rect 92216 327570 92244 335326
rect 92386 332480 92442 332489
rect 92386 332415 92442 332424
rect 90528 327542 90956 327570
rect 91816 327542 92244 327570
rect 88320 327406 88472 327434
rect 78586 327312 78642 327321
rect 78370 327284 78586 327298
rect 78384 327270 78586 327284
rect 78586 327247 78642 327256
rect 91264 327146 91600 327162
rect 92400 327146 92428 332415
rect 92846 331256 92902 331265
rect 92846 331191 92902 331200
rect 92860 327570 92888 331191
rect 93688 327570 93716 342246
rect 92552 327542 92888 327570
rect 93288 327542 93716 327570
rect 93872 327570 93900 355302
rect 95146 351112 95202 351121
rect 95146 351047 95202 351056
rect 95160 349194 95188 351047
rect 95160 349166 95372 349194
rect 95344 331158 95372 349166
rect 95332 331152 95384 331158
rect 95332 331094 95384 331100
rect 95884 331152 95936 331158
rect 95884 331094 95936 331100
rect 95792 331084 95844 331090
rect 95792 331026 95844 331032
rect 95054 330712 95110 330721
rect 95054 330647 95110 330656
rect 95068 327570 95096 330647
rect 95804 327570 95832 331026
rect 93872 327542 94024 327570
rect 94760 327542 95096 327570
rect 95496 327542 95832 327570
rect 95896 327570 95924 331094
rect 96540 331090 96568 360975
rect 97170 332888 97226 332897
rect 97170 332823 97226 332832
rect 96528 331084 96580 331090
rect 96528 331026 96580 331032
rect 97184 327570 97212 332823
rect 97276 331906 97304 369815
rect 97828 355366 97856 390374
rect 100666 390416 100722 390425
rect 98882 390374 99328 390402
rect 98826 390351 98882 390360
rect 99300 366382 99328 390374
rect 100722 390374 101168 390402
rect 100666 390351 100722 390360
rect 101140 389065 101168 390374
rect 102612 389162 102640 390918
rect 107934 390895 107990 390904
rect 114098 390960 114154 390969
rect 114154 390918 114448 390946
rect 114098 390895 114154 390904
rect 104990 390416 105046 390425
rect 103776 390374 104112 390402
rect 102600 389156 102652 389162
rect 102600 389098 102652 389104
rect 101126 389056 101182 389065
rect 101126 388991 101182 389000
rect 101954 389056 102010 389065
rect 101954 388991 102010 389000
rect 100116 388476 100168 388482
rect 100116 388418 100168 388424
rect 101404 388476 101456 388482
rect 101404 388418 101456 388424
rect 99288 366376 99340 366382
rect 99288 366318 99340 366324
rect 100128 364313 100156 388418
rect 100114 364304 100170 364313
rect 100114 364239 100170 364248
rect 100024 362976 100076 362982
rect 100024 362918 100076 362924
rect 97816 355360 97868 355366
rect 97816 355302 97868 355308
rect 100036 345014 100064 362918
rect 101416 352578 101444 388418
rect 101968 360233 101996 388991
rect 104084 385014 104112 390374
rect 106554 390416 106610 390425
rect 105046 390374 105432 390402
rect 104990 390351 105046 390360
rect 106610 390374 107332 390402
rect 106554 390351 106610 390360
rect 104072 385008 104124 385014
rect 104072 384950 104124 384956
rect 105004 381585 105032 390351
rect 105544 389156 105596 389162
rect 105544 389098 105596 389104
rect 104990 381576 105046 381585
rect 104990 381511 105046 381520
rect 102046 367160 102102 367169
rect 102046 367095 102102 367104
rect 101494 360224 101550 360233
rect 101494 360159 101550 360168
rect 101954 360224 102010 360233
rect 101954 360159 102010 360168
rect 101404 352572 101456 352578
rect 101404 352514 101456 352520
rect 100036 344986 100156 345014
rect 98642 339552 98698 339561
rect 98642 339487 98698 339496
rect 97264 331900 97316 331906
rect 97264 331842 97316 331848
rect 97908 331288 97960 331294
rect 97908 331230 97960 331236
rect 97920 330546 97948 331230
rect 97908 330540 97960 330546
rect 97908 330482 97960 330488
rect 98656 330449 98684 339487
rect 100128 331129 100156 344986
rect 101508 341562 101536 360159
rect 101956 346452 102008 346458
rect 101956 346394 102008 346400
rect 101496 341556 101548 341562
rect 101496 341498 101548 341504
rect 101968 331158 101996 346394
rect 101496 331152 101548 331158
rect 100114 331120 100170 331129
rect 101496 331094 101548 331100
rect 101956 331152 102008 331158
rect 101956 331094 102008 331100
rect 100114 331055 100170 331064
rect 99286 330576 99342 330585
rect 99286 330511 99342 330520
rect 97814 330440 97870 330449
rect 97814 330375 97870 330384
rect 98642 330440 98698 330449
rect 98642 330375 98698 330384
rect 97828 327570 97856 330375
rect 98550 330304 98606 330313
rect 98550 330239 98606 330248
rect 98564 327570 98592 330239
rect 99300 327570 99328 330511
rect 100024 330064 100076 330070
rect 100024 330006 100076 330012
rect 100036 327570 100064 330006
rect 95896 327542 96232 327570
rect 96968 327542 97212 327570
rect 97520 327542 97856 327570
rect 98256 327542 98592 327570
rect 98992 327542 99328 327570
rect 99728 327542 100064 327570
rect 100128 327570 100156 331055
rect 101508 327570 101536 331094
rect 102060 327570 102088 367095
rect 102784 365764 102836 365770
rect 102784 365706 102836 365712
rect 102692 340944 102744 340950
rect 102692 340886 102744 340892
rect 102508 331356 102560 331362
rect 102508 331298 102560 331304
rect 100128 327542 100464 327570
rect 101200 327542 101536 327570
rect 101936 327542 102088 327570
rect 102520 327434 102548 331298
rect 102704 329202 102732 340886
rect 102796 330070 102824 365706
rect 104808 352640 104860 352646
rect 104808 352582 104860 352588
rect 104256 330132 104308 330138
rect 104256 330074 104308 330080
rect 102784 330064 102836 330070
rect 102784 330006 102836 330012
rect 102704 329174 102824 329202
rect 102796 327570 102824 329174
rect 104268 327570 104296 330074
rect 104820 327570 104848 352582
rect 105556 345681 105584 389098
rect 107304 383654 107332 390374
rect 107948 388385 107976 390895
rect 115754 390688 115810 390697
rect 115810 390646 115888 390674
rect 115754 390623 115810 390632
rect 111504 390510 111656 390538
rect 108026 390416 108082 390425
rect 109498 390416 109554 390425
rect 108082 390374 108804 390402
rect 108026 390351 108082 390360
rect 107934 388376 107990 388385
rect 107934 388311 107990 388320
rect 108776 383654 108804 390374
rect 109554 390374 110184 390402
rect 109498 390351 109554 390360
rect 110156 385694 110184 390374
rect 111628 389230 111656 390510
rect 112640 390374 112976 390402
rect 111708 389836 111760 389842
rect 111708 389778 111760 389784
rect 111616 389224 111668 389230
rect 111616 389166 111668 389172
rect 111628 388686 111656 389166
rect 111616 388680 111668 388686
rect 111616 388622 111668 388628
rect 110144 385688 110196 385694
rect 110144 385630 110196 385636
rect 107304 383626 107516 383654
rect 108776 383626 108896 383654
rect 105634 381576 105690 381585
rect 105634 381511 105690 381520
rect 105648 352578 105676 381511
rect 107488 373318 107516 383626
rect 107476 373312 107528 373318
rect 107476 373254 107528 373260
rect 108868 370530 108896 383626
rect 108304 370524 108356 370530
rect 108304 370466 108356 370472
rect 108856 370524 108908 370530
rect 108856 370466 108908 370472
rect 107568 361616 107620 361622
rect 107568 361558 107620 361564
rect 105636 352572 105688 352578
rect 105636 352514 105688 352520
rect 105542 345672 105598 345681
rect 105542 345607 105598 345616
rect 105544 342372 105596 342378
rect 105544 342314 105596 342320
rect 104900 335436 104952 335442
rect 104900 335378 104952 335384
rect 102796 327542 103224 327570
rect 103960 327542 104296 327570
rect 104696 327542 104848 327570
rect 104912 327570 104940 335378
rect 105556 330138 105584 342314
rect 106464 338224 106516 338230
rect 106186 338192 106242 338201
rect 106464 338166 106516 338172
rect 106186 338127 106242 338136
rect 105544 330132 105596 330138
rect 105544 330074 105596 330080
rect 106200 327842 106228 338127
rect 106154 327814 106228 327842
rect 104912 327542 105432 327570
rect 106154 327556 106182 327814
rect 106476 327570 106504 338166
rect 107580 331158 107608 361558
rect 108316 358766 108344 370466
rect 111062 361856 111118 361865
rect 111062 361791 111118 361800
rect 109682 359000 109738 359009
rect 109682 358935 109738 358944
rect 107844 358760 107896 358766
rect 107844 358702 107896 358708
rect 108304 358760 108356 358766
rect 108304 358702 108356 358708
rect 107856 357474 107884 358702
rect 107844 357468 107896 357474
rect 107844 357410 107896 357416
rect 107568 331152 107620 331158
rect 107568 331094 107620 331100
rect 107856 327570 107884 357410
rect 108946 343768 109002 343777
rect 108946 343703 109002 343712
rect 108028 331152 108080 331158
rect 108028 331094 108080 331100
rect 106476 327542 106904 327570
rect 107640 327542 107884 327570
rect 108040 327570 108068 331094
rect 108304 330880 108356 330886
rect 108304 330822 108356 330828
rect 108316 330721 108344 330822
rect 108302 330712 108358 330721
rect 108302 330647 108358 330656
rect 108960 327842 108988 343703
rect 109696 338745 109724 358935
rect 110418 353424 110474 353433
rect 110418 353359 110474 353368
rect 110326 346624 110382 346633
rect 110326 346559 110382 346568
rect 109682 338736 109738 338745
rect 109682 338671 109738 338680
rect 110340 335354 110368 346559
rect 110432 345014 110460 353359
rect 111076 351286 111104 361791
rect 111720 353433 111748 389778
rect 112640 389065 112668 390374
rect 112626 389056 112682 389065
rect 112626 388991 112682 389000
rect 112444 388680 112496 388686
rect 112444 388622 112496 388628
rect 111798 354920 111854 354929
rect 111798 354855 111854 354864
rect 111706 353424 111762 353433
rect 111706 353359 111762 353368
rect 111064 351280 111116 351286
rect 111064 351222 111116 351228
rect 111812 345014 111840 354855
rect 112456 349858 112484 388622
rect 115110 382256 115166 382265
rect 115110 382191 115112 382200
rect 115164 382191 115166 382200
rect 115756 382220 115808 382226
rect 115112 382162 115164 382168
rect 115756 382162 115808 382168
rect 115768 380934 115796 382162
rect 115756 380928 115808 380934
rect 115756 380870 115808 380876
rect 115860 364449 115888 390646
rect 115938 390416 115994 390425
rect 120170 390416 120226 390425
rect 115994 390374 116104 390402
rect 117576 390374 117912 390402
rect 115938 390351 115994 390360
rect 114558 364440 114614 364449
rect 114558 364375 114614 364384
rect 115846 364440 115902 364449
rect 115846 364375 115902 364384
rect 112444 349852 112496 349858
rect 112444 349794 112496 349800
rect 110432 344986 110736 345014
rect 111812 344986 112024 345014
rect 108914 327814 108988 327842
rect 110064 335326 110368 335354
rect 108040 327542 108376 327570
rect 108914 327556 108942 327814
rect 110064 327570 110092 335326
rect 110604 330404 110656 330410
rect 110604 330346 110656 330352
rect 110616 327570 110644 330346
rect 109664 327542 110092 327570
rect 110400 327542 110644 327570
rect 110708 327570 110736 344986
rect 111706 340912 111762 340921
rect 111706 340847 111762 340856
rect 111720 330410 111748 340847
rect 111708 330404 111760 330410
rect 111708 330346 111760 330352
rect 111892 329860 111944 329866
rect 111892 329802 111944 329808
rect 111904 327729 111932 329802
rect 111890 327720 111946 327729
rect 111890 327655 111946 327664
rect 110708 327542 111136 327570
rect 111996 327434 112024 344986
rect 114468 339584 114520 339590
rect 114468 339526 114520 339532
rect 114376 331152 114428 331158
rect 114376 331094 114428 331100
rect 112810 330032 112866 330041
rect 112810 329967 112866 329976
rect 113640 329996 113692 330002
rect 112824 327570 112852 329967
rect 113640 329938 113692 329944
rect 113652 327570 113680 329938
rect 114388 327570 114416 331094
rect 114480 330002 114508 339526
rect 114468 329996 114520 330002
rect 114468 329938 114520 329944
rect 114572 327842 114600 364375
rect 115202 347984 115258 347993
rect 115202 347919 115258 347928
rect 115020 332716 115072 332722
rect 115020 332658 115072 332664
rect 115032 330546 115060 332658
rect 115216 330886 115244 347919
rect 115952 345817 115980 390351
rect 117884 389162 117912 390374
rect 118712 390374 119048 390402
rect 118712 389201 118740 390374
rect 120226 390374 120520 390402
rect 120170 390351 120226 390360
rect 118698 389192 118754 389201
rect 117872 389156 117924 389162
rect 118698 389127 118754 389136
rect 117872 389098 117924 389104
rect 118712 382294 118740 389127
rect 120184 388482 120212 390351
rect 120172 388476 120224 388482
rect 120172 388418 120224 388424
rect 118700 382288 118752 382294
rect 118700 382230 118752 382236
rect 119436 382288 119488 382294
rect 119436 382230 119488 382236
rect 119342 370016 119398 370025
rect 119342 369951 119398 369960
rect 118792 354000 118844 354006
rect 118792 353942 118844 353948
rect 118804 350606 118832 353942
rect 118792 350600 118844 350606
rect 118698 350568 118754 350577
rect 119356 350577 119384 369951
rect 119448 367810 119476 382230
rect 120736 371385 120764 434687
rect 120828 419529 120856 572698
rect 121460 548548 121512 548554
rect 121460 548490 121512 548496
rect 120908 444440 120960 444446
rect 120908 444382 120960 444388
rect 120920 442785 120948 444382
rect 120906 442776 120962 442785
rect 120906 442711 120962 442720
rect 121182 439920 121238 439929
rect 121182 439855 121238 439864
rect 121196 438938 121224 439855
rect 121184 438932 121236 438938
rect 121184 438874 121236 438880
rect 120814 419520 120870 419529
rect 120814 419455 120870 419464
rect 120828 390697 120856 419455
rect 121472 396953 121500 548490
rect 121564 428505 121592 578206
rect 123392 569220 123444 569226
rect 123392 569162 123444 569168
rect 122104 556232 122156 556238
rect 122104 556174 122156 556180
rect 121642 453248 121698 453257
rect 121642 453183 121698 453192
rect 121550 428496 121606 428505
rect 121550 428431 121606 428440
rect 121552 418124 121604 418130
rect 121552 418066 121604 418072
rect 121564 417353 121592 418066
rect 121550 417344 121606 417353
rect 121550 417279 121606 417288
rect 121458 396944 121514 396953
rect 121458 396879 121514 396888
rect 121472 396098 121500 396879
rect 121460 396092 121512 396098
rect 121460 396034 121512 396040
rect 121458 392592 121514 392601
rect 121458 392527 121514 392536
rect 120814 390688 120870 390697
rect 120814 390623 120870 390632
rect 120722 371376 120778 371385
rect 120722 371311 120778 371320
rect 119436 367804 119488 367810
rect 119436 367746 119488 367752
rect 120080 360256 120132 360262
rect 120080 360198 120132 360204
rect 118792 350542 118844 350548
rect 119342 350568 119398 350577
rect 118698 350503 118754 350512
rect 117228 347880 117280 347886
rect 117228 347822 117280 347828
rect 115938 345808 115994 345817
rect 115938 345743 115994 345752
rect 116582 342408 116638 342417
rect 116582 342343 116638 342352
rect 115940 336796 115992 336802
rect 115940 336738 115992 336744
rect 115664 332648 115716 332654
rect 115664 332590 115716 332596
rect 115204 330880 115256 330886
rect 115204 330822 115256 330828
rect 115020 330540 115072 330546
rect 115020 330482 115072 330488
rect 114572 327814 114646 327842
rect 112608 327542 112852 327570
rect 113344 327542 113680 327570
rect 114080 327542 114416 327570
rect 114618 327570 114646 327814
rect 115676 327570 115704 332590
rect 114618 327556 114784 327570
rect 114632 327542 114784 327556
rect 115368 327542 115704 327570
rect 115952 327570 115980 336738
rect 116596 331158 116624 342343
rect 116584 331152 116636 331158
rect 116584 331094 116636 331100
rect 117240 327570 117268 347822
rect 117318 347712 117374 347721
rect 117318 347647 117374 347656
rect 117332 346497 117360 347647
rect 117318 346488 117374 346497
rect 117318 346423 117374 346432
rect 117332 345014 117360 346423
rect 118606 345128 118662 345137
rect 118606 345063 118662 345072
rect 117332 344986 117912 345014
rect 117780 331152 117832 331158
rect 117780 331094 117832 331100
rect 117792 327570 117820 331094
rect 115952 327542 116104 327570
rect 116840 327542 117268 327570
rect 117576 327542 117820 327570
rect 117884 327570 117912 344986
rect 118620 331158 118648 345063
rect 118712 331158 118740 350503
rect 118608 331152 118660 331158
rect 118608 331094 118660 331100
rect 118700 331152 118752 331158
rect 118700 331094 118752 331100
rect 118804 327570 118832 350542
rect 119342 350503 119398 350512
rect 119436 331152 119488 331158
rect 119436 331094 119488 331100
rect 119448 327570 119476 331094
rect 120092 327570 120120 360198
rect 120736 352646 120764 371311
rect 121472 368966 121500 392527
rect 121564 389842 121592 417279
rect 121656 410553 121684 453183
rect 121642 410544 121698 410553
rect 121642 410479 121698 410488
rect 121656 409902 121684 410479
rect 121644 409896 121696 409902
rect 121644 409838 121696 409844
rect 122116 407114 122144 556174
rect 123116 458856 123168 458862
rect 123116 458798 123168 458804
rect 122932 457496 122984 457502
rect 122932 457438 122984 457444
rect 122944 424153 122972 457438
rect 123128 433129 123156 458798
rect 123114 433120 123170 433129
rect 123114 433055 123170 433064
rect 123298 428496 123354 428505
rect 123298 428431 123354 428440
rect 122930 424144 122986 424153
rect 122930 424079 122986 424088
rect 123206 424144 123262 424153
rect 123206 424079 123262 424088
rect 122746 422240 122802 422249
rect 122746 422175 122802 422184
rect 122760 412865 122788 422175
rect 123114 415168 123170 415177
rect 123114 415103 123116 415112
rect 123168 415103 123170 415112
rect 123116 415074 123168 415080
rect 123116 413976 123168 413982
rect 123116 413918 123168 413924
rect 122746 412856 122802 412865
rect 122746 412791 122802 412800
rect 123128 412729 123156 413918
rect 123114 412720 123170 412729
rect 123114 412655 123170 412664
rect 122746 412584 122802 412593
rect 122746 412519 122802 412528
rect 122104 407108 122156 407114
rect 122104 407050 122156 407056
rect 122760 403073 122788 412519
rect 123024 407108 123076 407114
rect 123024 407050 123076 407056
rect 122746 403064 122802 403073
rect 122746 402999 122802 403008
rect 122746 402928 122802 402937
rect 122746 402863 122802 402872
rect 122760 393417 122788 402863
rect 122746 393408 122802 393417
rect 122746 393343 122802 393352
rect 122746 393272 122802 393281
rect 122746 393207 122802 393216
rect 121552 389836 121604 389842
rect 121552 389778 121604 389784
rect 122760 383761 122788 393207
rect 123036 392601 123064 407050
rect 123022 392592 123078 392601
rect 123022 392527 123078 392536
rect 123128 384334 123156 412655
rect 123116 384328 123168 384334
rect 123116 384270 123168 384276
rect 122746 383752 122802 383761
rect 122746 383687 122802 383696
rect 122746 383616 122802 383625
rect 122746 383551 122802 383560
rect 122760 374105 122788 383551
rect 123220 380254 123248 424079
rect 123208 380248 123260 380254
rect 123208 380190 123260 380196
rect 122746 374096 122802 374105
rect 122746 374031 122802 374040
rect 122746 373960 122802 373969
rect 122746 373895 122802 373904
rect 121460 368960 121512 368966
rect 121460 368902 121512 368908
rect 122104 368960 122156 368966
rect 122104 368902 122156 368908
rect 121472 368558 121500 368902
rect 121460 368552 121512 368558
rect 121460 368494 121512 368500
rect 122116 363662 122144 368902
rect 122760 364585 122788 373895
rect 122746 364576 122802 364585
rect 122746 364511 122802 364520
rect 122746 364168 122802 364177
rect 122746 364103 122802 364112
rect 122104 363656 122156 363662
rect 122104 363598 122156 363604
rect 121458 361720 121514 361729
rect 121458 361655 121514 361664
rect 121472 356726 121500 361655
rect 121460 356720 121512 356726
rect 121460 356662 121512 356668
rect 122760 355337 122788 364103
rect 123312 360913 123340 428431
rect 123404 421977 123432 569162
rect 124220 557592 124272 557598
rect 124220 557534 124272 557540
rect 123576 456136 123628 456142
rect 123576 456078 123628 456084
rect 123390 421968 123446 421977
rect 123390 421903 123446 421912
rect 123404 421598 123432 421903
rect 123392 421592 123444 421598
rect 123392 421534 123444 421540
rect 123588 406201 123616 456078
rect 124128 444372 124180 444378
rect 124128 444314 124180 444320
rect 124140 444281 124168 444314
rect 124126 444272 124182 444281
rect 124126 444207 124182 444216
rect 124126 442096 124182 442105
rect 124126 442031 124182 442040
rect 124140 441658 124168 442031
rect 124128 441652 124180 441658
rect 124128 441594 124180 441600
rect 123852 438184 123904 438190
rect 123852 438126 123904 438132
rect 123864 437753 123892 438126
rect 123850 437744 123906 437753
rect 123850 437679 123906 437688
rect 124126 433120 124182 433129
rect 124126 433055 124182 433064
rect 124140 432614 124168 433055
rect 124128 432608 124180 432614
rect 124128 432550 124180 432556
rect 124128 408400 124180 408406
rect 124126 408368 124128 408377
rect 124180 408368 124182 408377
rect 124126 408303 124182 408312
rect 123574 406192 123630 406201
rect 123574 406127 123630 406136
rect 123588 405890 123616 406127
rect 123576 405884 123628 405890
rect 123576 405826 123628 405832
rect 124128 401600 124180 401606
rect 124126 401568 124128 401577
rect 124180 401568 124182 401577
rect 124126 401503 124182 401512
rect 123666 399392 123722 399401
rect 123666 399327 123722 399336
rect 123680 398886 123708 399327
rect 123668 398880 123720 398886
rect 123668 398822 123720 398828
rect 124126 394768 124182 394777
rect 124232 394754 124260 557534
rect 124876 536761 124904 702986
rect 126244 702908 126296 702914
rect 126244 702850 126296 702856
rect 125600 569968 125652 569974
rect 125600 569910 125652 569916
rect 124862 536752 124918 536761
rect 124862 536687 124918 536696
rect 124404 456068 124456 456074
rect 124404 456010 124456 456016
rect 124312 448656 124364 448662
rect 124312 448598 124364 448604
rect 124182 394726 124260 394754
rect 124126 394703 124182 394712
rect 123482 367704 123538 367713
rect 123482 367639 123538 367648
rect 123298 360904 123354 360913
rect 123298 360839 123354 360848
rect 122840 356108 122892 356114
rect 122840 356050 122892 356056
rect 122746 355328 122802 355337
rect 122746 355263 122802 355272
rect 122748 354000 122800 354006
rect 122748 353942 122800 353948
rect 120724 352640 120776 352646
rect 120724 352582 120776 352588
rect 121366 343904 121422 343913
rect 121366 343839 121422 343848
rect 120722 338464 120778 338473
rect 120722 338399 120778 338408
rect 120736 330585 120764 338399
rect 120722 330576 120778 330585
rect 120722 330511 120778 330520
rect 121380 327570 121408 343839
rect 122102 328808 122158 328817
rect 122102 328743 122158 328752
rect 122116 327570 122144 328743
rect 122760 327570 122788 353942
rect 122852 351218 122880 356050
rect 123496 354754 123524 367639
rect 123484 354748 123536 354754
rect 123484 354690 123536 354696
rect 122840 351212 122892 351218
rect 122840 351154 122892 351160
rect 122932 346996 122984 347002
rect 122932 346938 122984 346944
rect 122944 345273 122972 346938
rect 122930 345264 122986 345273
rect 122930 345199 122986 345208
rect 122944 335354 122972 345199
rect 122852 335326 122972 335354
rect 122852 331158 122880 335326
rect 122840 331152 122892 331158
rect 122840 331094 122892 331100
rect 123496 328545 123524 354690
rect 124324 351121 124352 448598
rect 124416 415138 124444 456010
rect 124864 445868 124916 445874
rect 124864 445810 124916 445816
rect 124876 435305 124904 445810
rect 124862 435296 124918 435305
rect 124862 435231 124918 435240
rect 124404 415132 124456 415138
rect 124404 415074 124456 415080
rect 125612 413982 125640 569910
rect 126256 545766 126284 702850
rect 129004 702704 129056 702710
rect 129004 702646 129056 702652
rect 126980 571396 127032 571402
rect 126980 571338 127032 571344
rect 126244 545760 126296 545766
rect 126244 545702 126296 545708
rect 126336 452736 126388 452742
rect 126336 452678 126388 452684
rect 125692 447840 125744 447846
rect 125692 447782 125744 447788
rect 125704 438190 125732 447782
rect 126242 444680 126298 444689
rect 126242 444615 126298 444624
rect 125692 438184 125744 438190
rect 125692 438126 125744 438132
rect 125600 413976 125652 413982
rect 125600 413918 125652 413924
rect 124864 405884 124916 405890
rect 124864 405826 124916 405832
rect 124876 360330 124904 405826
rect 124956 398880 125008 398886
rect 124956 398822 125008 398828
rect 124968 392018 124996 398822
rect 124956 392012 125008 392018
rect 124956 391954 125008 391960
rect 124968 391406 124996 391954
rect 124956 391400 125008 391406
rect 124956 391342 125008 391348
rect 124956 374672 125008 374678
rect 124956 374614 125008 374620
rect 124864 360324 124916 360330
rect 124864 360266 124916 360272
rect 124968 354674 124996 374614
rect 125600 360324 125652 360330
rect 125600 360266 125652 360272
rect 125612 358873 125640 360266
rect 125598 358864 125654 358873
rect 125598 358799 125654 358808
rect 124876 354646 124996 354674
rect 124310 351112 124366 351121
rect 124310 351047 124366 351056
rect 124876 350713 124904 354646
rect 124862 350704 124918 350713
rect 124862 350639 124918 350648
rect 124128 347064 124180 347070
rect 124128 347006 124180 347012
rect 124140 346633 124168 347006
rect 124126 346624 124182 346633
rect 124126 346559 124182 346568
rect 123668 331152 123720 331158
rect 123668 331094 123720 331100
rect 123482 328536 123538 328545
rect 123482 328471 123538 328480
rect 123496 327570 123524 328471
rect 117884 327542 118312 327570
rect 118804 327542 119048 327570
rect 119448 327542 119784 327570
rect 120092 327542 120336 327570
rect 121072 327542 121408 327570
rect 121808 327542 122144 327570
rect 122544 327542 122788 327570
rect 123280 327542 123524 327570
rect 123680 327570 123708 331094
rect 124876 328506 124904 350639
rect 125322 334112 125378 334121
rect 125322 334047 125378 334056
rect 124864 328500 124916 328506
rect 124864 328442 124916 328448
rect 124876 327570 124904 328442
rect 123680 327542 124016 327570
rect 124752 327542 124904 327570
rect 102520 327406 102672 327434
rect 111872 327406 112024 327434
rect 114756 327214 114784 327542
rect 125336 327298 125364 334047
rect 125612 331158 125640 358799
rect 126256 357377 126284 444615
rect 126348 367130 126376 452678
rect 126992 418130 127020 571338
rect 128360 567860 128412 567866
rect 128360 567802 128412 567808
rect 126980 418124 127032 418130
rect 126980 418066 127032 418072
rect 126980 415132 127032 415138
rect 126980 415074 127032 415080
rect 126336 367124 126388 367130
rect 126336 367066 126388 367072
rect 125690 357368 125746 357377
rect 125690 357303 125746 357312
rect 126242 357368 126298 357377
rect 126242 357303 126298 357312
rect 125704 356153 125732 357303
rect 125690 356144 125746 356153
rect 125690 356079 125746 356088
rect 125600 331152 125652 331158
rect 125600 331094 125652 331100
rect 125704 327570 125732 356079
rect 126348 354006 126376 367066
rect 126992 360913 127020 415074
rect 128372 408406 128400 567802
rect 129016 544406 129044 702646
rect 129004 544400 129056 544406
rect 129004 544342 129056 544348
rect 130396 536790 130424 703190
rect 133144 700324 133196 700330
rect 133144 700266 133196 700272
rect 132500 590708 132552 590714
rect 132500 590650 132552 590656
rect 130476 552084 130528 552090
rect 130476 552026 130528 552032
rect 130384 536784 130436 536790
rect 130384 536726 130436 536732
rect 128450 536072 128506 536081
rect 128450 536007 128506 536016
rect 128360 408400 128412 408406
rect 128360 408342 128412 408348
rect 128372 407794 128400 408342
rect 128360 407788 128412 407794
rect 128360 407730 128412 407736
rect 128464 387802 128492 536007
rect 130382 448624 130438 448633
rect 130382 448559 130438 448568
rect 128452 387796 128504 387802
rect 128452 387738 128504 387744
rect 126978 360904 127034 360913
rect 126978 360839 127034 360848
rect 128360 360324 128412 360330
rect 128360 360266 128412 360272
rect 126978 359408 127034 359417
rect 126978 359343 127034 359352
rect 126992 357649 127020 359343
rect 126978 357640 127034 357649
rect 126978 357575 127034 357584
rect 126336 354000 126388 354006
rect 126336 353942 126388 353948
rect 126992 345014 127020 357575
rect 128372 345014 128400 360266
rect 129738 356008 129794 356017
rect 129738 355943 129794 355952
rect 129752 354793 129780 355943
rect 129738 354784 129794 354793
rect 129738 354719 129794 354728
rect 129004 349172 129056 349178
rect 129004 349114 129056 349120
rect 126992 344986 127848 345014
rect 128372 344986 128584 345014
rect 126428 331152 126480 331158
rect 126428 331094 126480 331100
rect 126440 327570 126468 331094
rect 127716 330132 127768 330138
rect 127716 330074 127768 330080
rect 127728 327570 127756 330074
rect 125704 327542 126040 327570
rect 126440 327542 126776 327570
rect 127512 327542 127756 327570
rect 127820 327570 127848 344986
rect 128556 327570 128584 344986
rect 129016 330138 129044 349114
rect 129004 330132 129056 330138
rect 129004 330074 129056 330080
rect 129752 327842 129780 354719
rect 130396 352617 130424 448559
rect 130488 389230 130516 552026
rect 132512 444378 132540 590650
rect 133156 538218 133184 700266
rect 133880 563100 133932 563106
rect 133880 563042 133932 563048
rect 133144 538212 133196 538218
rect 133144 538154 133196 538160
rect 132500 444372 132552 444378
rect 132500 444314 132552 444320
rect 133788 444372 133840 444378
rect 133788 444314 133840 444320
rect 133800 443698 133828 444314
rect 133788 443692 133840 443698
rect 133788 443634 133840 443640
rect 133144 441652 133196 441658
rect 133144 441594 133196 441600
rect 130476 389224 130528 389230
rect 130476 389166 130528 389172
rect 130476 380928 130528 380934
rect 130476 380870 130528 380876
rect 130488 356017 130516 380870
rect 133156 370598 133184 441594
rect 133892 401606 133920 563042
rect 136652 541686 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202604 703656 202656 703662
rect 202604 703598 202656 703604
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702545 154160 703520
rect 154118 702536 154174 702545
rect 154118 702471 154174 702480
rect 170324 702434 170352 703520
rect 202616 703474 202644 703598
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234988 703588 235040 703594
rect 234988 703530 235040 703536
rect 202800 703474 202828 703520
rect 202616 703446 202828 703474
rect 169772 702406 170352 702434
rect 169772 596834 169800 702406
rect 218992 700330 219020 703520
rect 235000 703474 235028 703530
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267464 703520 267516 703526
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 703474 267688 703520
rect 267516 703468 267688 703474
rect 267464 703462 267688 703468
rect 267476 703446 267688 703462
rect 283852 703390 283880 703520
rect 300136 703458 300164 703520
rect 300124 703452 300176 703458
rect 300124 703394 300176 703400
rect 283840 703384 283892 703390
rect 283840 703326 283892 703332
rect 332520 703322 332548 703520
rect 332508 703316 332560 703322
rect 332508 703258 332560 703264
rect 348804 703186 348832 703520
rect 348792 703180 348844 703186
rect 348792 703122 348844 703128
rect 364996 702982 365024 703520
rect 397472 703118 397500 703520
rect 413664 703254 413692 703520
rect 413652 703248 413704 703254
rect 413652 703190 413704 703196
rect 397460 703112 397512 703118
rect 397460 703054 397512 703060
rect 429856 703050 429884 703520
rect 429844 703044 429896 703050
rect 429844 702986 429896 702992
rect 364984 702976 365036 702982
rect 364984 702918 365036 702924
rect 462332 702914 462360 703520
rect 462320 702908 462372 702914
rect 462320 702850 462372 702856
rect 478524 702778 478552 703520
rect 494808 702846 494836 703520
rect 494796 702840 494848 702846
rect 494796 702782 494848 702788
rect 478512 702772 478564 702778
rect 478512 702714 478564 702720
rect 527192 702642 527220 703520
rect 543476 702710 543504 703520
rect 543464 702704 543516 702710
rect 543464 702646 543516 702652
rect 527180 702636 527232 702642
rect 527180 702578 527232 702584
rect 559668 702506 559696 703520
rect 580264 702568 580316 702574
rect 580264 702510 580316 702516
rect 559656 702500 559708 702506
rect 559656 702442 559708 702448
rect 218980 700324 219032 700330
rect 218980 700266 219032 700272
rect 580276 670721 580304 702510
rect 582378 697232 582434 697241
rect 582378 697167 582434 697176
rect 580262 670712 580318 670721
rect 580262 670647 580318 670656
rect 169760 596828 169812 596834
rect 169760 596770 169812 596776
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 589966 580212 590951
rect 580172 589960 580224 589966
rect 580172 589902 580224 589908
rect 141424 586560 141476 586566
rect 141424 586502 141476 586508
rect 136640 541680 136692 541686
rect 136640 541622 136692 541628
rect 135168 432608 135220 432614
rect 135168 432550 135220 432556
rect 133880 401600 133932 401606
rect 133880 401542 133932 401548
rect 135076 401600 135128 401606
rect 135076 401542 135128 401548
rect 135088 400926 135116 401542
rect 135076 400920 135128 400926
rect 135076 400862 135128 400868
rect 133144 370592 133196 370598
rect 133144 370534 133196 370540
rect 135074 367296 135130 367305
rect 135074 367231 135130 367240
rect 132500 358896 132552 358902
rect 132500 358838 132552 358844
rect 132408 356176 132460 356182
rect 132408 356118 132460 356124
rect 130474 356008 130530 356017
rect 130474 355943 130530 355952
rect 130382 352608 130438 352617
rect 130382 352543 130438 352552
rect 129832 345160 129884 345166
rect 129832 345102 129884 345108
rect 129844 345014 129872 345102
rect 129844 344986 130056 345014
rect 129706 327814 129780 327842
rect 127820 327542 128248 327570
rect 128556 327542 128984 327570
rect 129706 327556 129734 327814
rect 130028 327570 130056 344986
rect 132420 335354 132448 356118
rect 132144 335326 132448 335354
rect 131486 329896 131542 329905
rect 131486 329831 131542 329840
rect 131500 327570 131528 329831
rect 132144 327570 132172 335326
rect 132512 327842 132540 358838
rect 132592 353388 132644 353394
rect 132592 353330 132644 353336
rect 132604 345014 132632 353330
rect 132604 344986 132816 345014
rect 130028 327542 130456 327570
rect 131192 327542 131528 327570
rect 131744 327542 132172 327570
rect 132466 327814 132540 327842
rect 132466 327556 132494 327814
rect 132788 327570 132816 344986
rect 134524 340196 134576 340202
rect 134524 340138 134576 340144
rect 134248 339516 134300 339522
rect 134248 339458 134300 339464
rect 134156 329860 134208 329866
rect 134156 329802 134208 329808
rect 134168 327570 134196 329802
rect 132788 327542 133216 327570
rect 133952 327542 134196 327570
rect 134260 327570 134288 339458
rect 134536 329186 134564 340138
rect 135088 329866 135116 367231
rect 135180 347177 135208 432550
rect 135904 407788 135956 407794
rect 135904 407730 135956 407736
rect 135916 367033 135944 407730
rect 136652 385014 136680 541622
rect 137282 444544 137338 444553
rect 137282 444479 137338 444488
rect 136640 385008 136692 385014
rect 136640 384950 136692 384956
rect 137100 385008 137152 385014
rect 137100 384950 137152 384956
rect 137112 384334 137140 384950
rect 137100 384328 137152 384334
rect 137100 384270 137152 384276
rect 137296 372230 137324 444479
rect 137284 372224 137336 372230
rect 137284 372166 137336 372172
rect 137928 372224 137980 372230
rect 137928 372166 137980 372172
rect 137940 371278 137968 372166
rect 137928 371272 137980 371278
rect 137928 371214 137980 371220
rect 135902 367024 135958 367033
rect 135902 366959 135958 366968
rect 136640 364472 136692 364478
rect 136640 364414 136692 364420
rect 135904 357536 135956 357542
rect 135904 357478 135956 357484
rect 135166 347168 135222 347177
rect 135166 347103 135222 347112
rect 135258 335744 135314 335753
rect 135258 335679 135314 335688
rect 135272 329866 135300 335679
rect 135916 331809 135944 357478
rect 136652 345014 136680 364414
rect 136652 344986 137048 345014
rect 135902 331800 135958 331809
rect 135902 331735 135958 331744
rect 136914 331528 136970 331537
rect 136914 331463 136970 331472
rect 135076 329860 135128 329866
rect 135076 329802 135128 329808
rect 135260 329860 135312 329866
rect 135260 329802 135312 329808
rect 135812 329860 135864 329866
rect 135812 329802 135864 329808
rect 134524 329180 134576 329186
rect 134524 329122 134576 329128
rect 135260 329112 135312 329118
rect 135260 329054 135312 329060
rect 135272 328953 135300 329054
rect 135258 328944 135314 328953
rect 135258 328879 135314 328888
rect 135272 327570 135300 328879
rect 135824 327570 135852 329802
rect 136928 327842 136956 331463
rect 136882 327814 136956 327842
rect 134260 327542 134688 327570
rect 135272 327542 135424 327570
rect 135824 327542 136160 327570
rect 136882 327556 136910 327814
rect 137020 327570 137048 344986
rect 137940 331158 137968 371214
rect 141436 369073 141464 586502
rect 580262 577688 580318 577697
rect 580262 577623 580318 577632
rect 579802 537840 579858 537849
rect 579802 537775 579858 537784
rect 579816 537538 579844 537775
rect 579804 537532 579856 537538
rect 579804 537474 579856 537480
rect 580276 534070 580304 577623
rect 582392 536081 582420 697167
rect 582470 683904 582526 683913
rect 582470 683839 582526 683848
rect 582484 577522 582512 683839
rect 582562 644056 582618 644065
rect 582562 643991 582618 644000
rect 582472 577516 582524 577522
rect 582472 577458 582524 577464
rect 582472 554804 582524 554810
rect 582472 554746 582524 554752
rect 582378 536072 582434 536081
rect 582378 536007 582434 536016
rect 580264 534064 580316 534070
rect 580264 534006 580316 534012
rect 582484 524521 582512 554746
rect 582576 539578 582604 643991
rect 582654 630864 582710 630873
rect 582654 630799 582710 630808
rect 582668 540938 582696 630799
rect 582746 617536 582802 617545
rect 582746 617471 582802 617480
rect 582760 595513 582788 617471
rect 582746 595504 582802 595513
rect 582746 595439 582802 595448
rect 582748 593428 582800 593434
rect 582748 593370 582800 593376
rect 582760 564369 582788 593370
rect 582746 564360 582802 564369
rect 582746 564295 582802 564304
rect 582656 540932 582708 540938
rect 582656 540874 582708 540880
rect 582564 539572 582616 539578
rect 582564 539514 582616 539520
rect 582470 524512 582526 524521
rect 582470 524447 582526 524456
rect 580170 511320 580226 511329
rect 580170 511255 580172 511264
rect 580224 511255 580226 511264
rect 580172 511226 580224 511232
rect 582378 484664 582434 484673
rect 582378 484599 582434 484608
rect 169022 458280 169078 458289
rect 169022 458215 169078 458224
rect 161480 454096 161532 454102
rect 161480 454038 161532 454044
rect 160100 450016 160152 450022
rect 160100 449958 160152 449964
rect 144184 444508 144236 444514
rect 144184 444450 144236 444456
rect 141422 369064 141478 369073
rect 141422 368999 141478 369008
rect 138018 367024 138074 367033
rect 138018 366959 138074 366968
rect 138032 365809 138060 366959
rect 138018 365800 138074 365809
rect 138018 365735 138074 365744
rect 137928 331152 137980 331158
rect 137928 331094 137980 331100
rect 138032 327570 138060 365735
rect 144196 352306 144224 444450
rect 157984 438184 158036 438190
rect 157984 438126 158036 438132
rect 148324 421592 148376 421598
rect 148324 421534 148376 421540
rect 145564 376032 145616 376038
rect 145564 375974 145616 375980
rect 144828 368552 144880 368558
rect 144828 368494 144880 368500
rect 144184 352300 144236 352306
rect 144184 352242 144236 352248
rect 144736 352300 144788 352306
rect 144736 352242 144788 352248
rect 144748 351966 144776 352242
rect 144736 351960 144788 351966
rect 144736 351902 144788 351908
rect 140870 349480 140926 349489
rect 140870 349415 140926 349424
rect 140780 347064 140832 347070
rect 140884 347041 140912 349415
rect 140780 347006 140832 347012
rect 140870 347032 140926 347041
rect 140792 346633 140820 347006
rect 140870 346967 140926 346976
rect 140778 346624 140834 346633
rect 140778 346559 140834 346568
rect 142804 346520 142856 346526
rect 142804 346462 142856 346468
rect 139306 342544 139362 342553
rect 139306 342479 139362 342488
rect 139320 327570 139348 342479
rect 142066 339824 142122 339833
rect 142066 339759 142122 339768
rect 141424 332716 141476 332722
rect 141424 332658 141476 332664
rect 140870 331392 140926 331401
rect 140870 331327 140926 331336
rect 139400 331152 139452 331158
rect 139400 331094 139452 331100
rect 137020 327542 137448 327570
rect 138032 327542 138184 327570
rect 138920 327542 139348 327570
rect 139412 327570 139440 331094
rect 140688 331084 140740 331090
rect 140688 331026 140740 331032
rect 139766 328672 139822 328681
rect 139766 328607 139822 328616
rect 139412 327542 139656 327570
rect 125336 327270 125488 327298
rect 114744 327208 114796 327214
rect 114744 327150 114796 327156
rect 91264 327140 91612 327146
rect 91264 327134 91560 327140
rect 91560 327082 91612 327088
rect 92388 327140 92440 327146
rect 92388 327082 92440 327088
rect 139780 327078 139808 328607
rect 140700 327570 140728 331026
rect 140780 330540 140832 330546
rect 140780 330482 140832 330488
rect 140792 329089 140820 330482
rect 140884 330449 140912 331327
rect 140870 330440 140926 330449
rect 140870 330375 140926 330384
rect 140778 329080 140834 329089
rect 140778 329015 140834 329024
rect 140778 328808 140834 328817
rect 140778 328743 140834 328752
rect 140792 327865 140820 328743
rect 140778 327856 140834 327865
rect 140778 327791 140834 327800
rect 141436 327570 141464 332658
rect 142080 327570 142108 339759
rect 142816 331090 142844 346462
rect 142896 341012 142948 341018
rect 142896 340954 142948 340960
rect 142908 334626 142936 340954
rect 142896 334620 142948 334626
rect 142896 334562 142948 334568
rect 144460 334076 144512 334082
rect 144460 334018 144512 334024
rect 144184 331152 144236 331158
rect 144184 331094 144236 331100
rect 142804 331084 142856 331090
rect 142804 331026 142856 331032
rect 142894 330168 142950 330177
rect 142894 330103 142950 330112
rect 142908 327570 142936 330103
rect 144196 327570 144224 331094
rect 140392 327542 140728 327570
rect 141128 327542 141464 327570
rect 141864 327542 142108 327570
rect 142600 327542 142936 327570
rect 143888 327542 144224 327570
rect 144472 327298 144500 334018
rect 144748 331090 144776 351902
rect 144840 331158 144868 368494
rect 145576 352209 145604 375974
rect 147680 361684 147732 361690
rect 147680 361626 147732 361632
rect 144918 352200 144974 352209
rect 144918 352135 144974 352144
rect 145562 352200 145618 352209
rect 145562 352135 145618 352144
rect 144828 331152 144880 331158
rect 144828 331094 144880 331100
rect 144736 331084 144788 331090
rect 144736 331026 144788 331032
rect 144932 327570 144960 352135
rect 147692 345014 147720 361626
rect 147692 344986 147904 345014
rect 146208 334008 146260 334014
rect 146208 333950 146260 333956
rect 146220 327570 146248 333950
rect 146484 331084 146536 331090
rect 146484 331026 146536 331032
rect 144932 327542 145360 327570
rect 146096 327542 146248 327570
rect 146496 327570 146524 331026
rect 147876 327570 147904 344986
rect 148336 328545 148364 421534
rect 155224 385688 155276 385694
rect 155224 385630 155276 385636
rect 150256 374128 150308 374134
rect 150256 374070 150308 374076
rect 150268 364313 150296 374070
rect 150348 372632 150400 372638
rect 150348 372574 150400 372580
rect 150254 364304 150310 364313
rect 150254 364239 150310 364248
rect 150268 363225 150296 364239
rect 150254 363216 150310 363225
rect 150254 363151 150310 363160
rect 148322 328536 148378 328545
rect 148322 328471 148378 328480
rect 150360 327842 150388 372574
rect 150438 363216 150494 363225
rect 150438 363151 150494 363160
rect 150452 345014 150480 363151
rect 154672 355360 154724 355366
rect 154672 355302 154724 355308
rect 153842 345672 153898 345681
rect 153842 345607 153898 345616
rect 150452 344986 150664 345014
rect 150636 331214 150664 344986
rect 153856 335354 153884 345607
rect 154684 345014 154712 355302
rect 154684 344986 154804 345014
rect 153672 335326 153884 335354
rect 150636 331186 150756 331214
rect 150314 327814 150388 327842
rect 146496 327542 146832 327570
rect 147876 327542 148304 327570
rect 150314 327556 150342 327814
rect 144472 327270 144624 327298
rect 149888 327208 149940 327214
rect 147218 327176 147274 327185
rect 147274 327134 147568 327162
rect 149592 327156 149888 327162
rect 150728 327185 150756 331186
rect 153672 329934 153700 335326
rect 153660 329928 153712 329934
rect 153660 329870 153712 329876
rect 151636 329860 151688 329866
rect 151636 329802 151688 329808
rect 149592 327150 149940 327156
rect 150714 327176 150770 327185
rect 149592 327134 149928 327150
rect 147218 327111 147274 327120
rect 150770 327134 151064 327162
rect 150714 327111 150770 327120
rect 151648 327078 151676 329802
rect 152096 328500 152148 328506
rect 152096 328442 152148 328448
rect 152108 327570 152136 328442
rect 153672 327570 153700 329870
rect 154776 328454 154804 344986
rect 154776 328426 154988 328454
rect 151800 327542 152136 327570
rect 153272 327542 153700 327570
rect 153660 327208 153712 327214
rect 153658 327176 153660 327185
rect 154304 327208 154356 327214
rect 153712 327176 153714 327185
rect 154008 327156 154304 327162
rect 154008 327150 154356 327156
rect 154008 327134 154344 327150
rect 153658 327111 153714 327120
rect 139768 327072 139820 327078
rect 139768 327014 139820 327020
rect 151636 327072 151688 327078
rect 154210 327040 154266 327049
rect 151636 327014 151688 327020
rect 152536 327010 152872 327026
rect 152536 327004 152884 327010
rect 152536 326998 152832 327004
rect 154560 326998 154896 327026
rect 154210 326975 154212 326984
rect 152832 326946 152884 326952
rect 154264 326975 154266 326984
rect 154212 326946 154264 326952
rect 71412 326936 71464 326942
rect 68008 326868 68060 326874
rect 68008 326810 68060 326816
rect 68098 326768 68154 326777
rect 68098 326703 68154 326712
rect 68112 325718 68140 326703
rect 68664 326505 68692 326878
rect 70964 326862 71208 326890
rect 143448 326936 143500 326942
rect 71412 326878 71464 326884
rect 143152 326884 143448 326890
rect 149152 326936 149204 326942
rect 143152 326878 143500 326884
rect 148856 326884 149152 326890
rect 148856 326878 149204 326884
rect 143152 326862 143488 326878
rect 148856 326862 149192 326878
rect 68650 326496 68706 326505
rect 68650 326431 68706 326440
rect 68100 325712 68152 325718
rect 68100 325654 68152 325660
rect 154868 325009 154896 326998
rect 154854 325000 154910 325009
rect 154854 324935 154910 324944
rect 154960 323626 154988 328426
rect 154684 323598 154988 323626
rect 67822 321600 67878 321609
rect 67822 321535 67878 321544
rect 67730 312080 67786 312089
rect 67730 312015 67786 312024
rect 154684 277001 154712 323598
rect 154764 322584 154816 322590
rect 154764 322526 154816 322532
rect 154776 321638 154804 322526
rect 154764 321632 154816 321638
rect 154764 321574 154816 321580
rect 154670 276992 154726 277001
rect 154670 276927 154726 276936
rect 67638 268832 67694 268841
rect 67638 268767 67694 268776
rect 67652 267734 67680 268767
rect 67652 267706 67864 267734
rect 67638 255232 67694 255241
rect 67638 255167 67694 255176
rect 67548 240780 67600 240786
rect 67548 240722 67600 240728
rect 67362 239864 67418 239873
rect 67362 239799 67418 239808
rect 67270 222864 67326 222873
rect 67270 222799 67326 222808
rect 67178 217288 67234 217297
rect 67178 217223 67234 217232
rect 64696 213920 64748 213926
rect 64696 213862 64748 213868
rect 67652 205601 67680 255167
rect 67730 245712 67786 245721
rect 67730 245647 67786 245656
rect 67744 215286 67772 245647
rect 67836 237153 67864 267706
rect 154776 264761 154804 321574
rect 155236 296714 155264 385630
rect 155960 371884 156012 371890
rect 155960 371826 156012 371832
rect 155592 361684 155644 361690
rect 155592 361626 155644 361632
rect 155604 356046 155632 361626
rect 155592 356040 155644 356046
rect 155592 355982 155644 355988
rect 155316 352572 155368 352578
rect 155316 352514 155368 352520
rect 155328 322590 155356 352514
rect 155316 322584 155368 322590
rect 155316 322526 155368 322532
rect 155972 315382 156000 371826
rect 157338 364984 157394 364993
rect 157338 364919 157394 364928
rect 156694 353968 156750 353977
rect 156694 353903 156750 353912
rect 156052 349852 156104 349858
rect 156052 349794 156104 349800
rect 156064 325417 156092 349794
rect 156234 328536 156290 328545
rect 156234 328471 156290 328480
rect 156050 325408 156106 325417
rect 156050 325343 156106 325352
rect 156064 324970 156092 325343
rect 156052 324964 156104 324970
rect 156052 324906 156104 324912
rect 156050 324320 156106 324329
rect 156050 324255 156106 324264
rect 156144 324284 156196 324290
rect 156064 323474 156092 324255
rect 156144 324226 156196 324232
rect 156052 323468 156104 323474
rect 156052 323410 156104 323416
rect 156156 323241 156184 324226
rect 156142 323232 156198 323241
rect 156142 323167 156198 323176
rect 156050 322144 156106 322153
rect 156050 322079 156106 322088
rect 156064 321978 156092 322079
rect 156052 321972 156104 321978
rect 156052 321914 156104 321920
rect 156248 321554 156276 328471
rect 156156 321526 156276 321554
rect 155960 315376 156012 315382
rect 155960 315318 156012 315324
rect 155972 314809 156000 315318
rect 155958 314800 156014 314809
rect 155958 314735 156014 314744
rect 156156 308553 156184 321526
rect 156602 321056 156658 321065
rect 156602 320991 156658 321000
rect 156616 320210 156644 320991
rect 156604 320204 156656 320210
rect 156604 320146 156656 320152
rect 156602 318608 156658 318617
rect 156602 318543 156658 318552
rect 156142 308544 156198 308553
rect 156142 308479 156198 308488
rect 156510 307456 156566 307465
rect 156510 307391 156566 307400
rect 156524 306406 156552 307391
rect 156512 306400 156564 306406
rect 156512 306342 156564 306348
rect 156050 304192 156106 304201
rect 156050 304127 156106 304136
rect 156064 303686 156092 304127
rect 156052 303680 156104 303686
rect 156052 303622 156104 303628
rect 156418 297936 156474 297945
rect 156418 297871 156474 297880
rect 154868 296686 155264 296714
rect 154868 294030 154896 296686
rect 156432 296002 156460 297871
rect 156420 295996 156472 296002
rect 156420 295938 156472 295944
rect 156328 295316 156380 295322
rect 156328 295258 156380 295264
rect 156340 294681 156368 295258
rect 156326 294672 156382 294681
rect 156326 294607 156382 294616
rect 154856 294024 154908 294030
rect 154856 293966 154908 293972
rect 154762 264752 154818 264761
rect 154762 264687 154818 264696
rect 154868 262041 154896 293966
rect 156234 288416 156290 288425
rect 156234 288351 156290 288360
rect 156248 287162 156276 288351
rect 156236 287156 156288 287162
rect 156236 287098 156288 287104
rect 156328 287088 156380 287094
rect 156328 287030 156380 287036
rect 156340 285161 156368 287030
rect 156326 285152 156382 285161
rect 156326 285087 156382 285096
rect 156512 274644 156564 274650
rect 156512 274586 156564 274592
rect 156524 273737 156552 274586
rect 156510 273728 156566 273737
rect 156510 273663 156566 273672
rect 155866 264208 155922 264217
rect 155866 264143 155922 264152
rect 154854 262032 154910 262041
rect 154854 261967 154910 261976
rect 68190 258768 68246 258777
rect 68190 258703 68246 258712
rect 68204 258058 68232 258703
rect 68192 258052 68244 258058
rect 68192 257994 68244 258000
rect 67914 250336 67970 250345
rect 67914 250271 67970 250280
rect 67928 248334 67956 250271
rect 67916 248328 67968 248334
rect 67916 248270 67968 248276
rect 154856 245676 154908 245682
rect 154856 245618 154908 245624
rect 73896 242072 73948 242078
rect 70306 242040 70362 242049
rect 150072 242072 150124 242078
rect 135994 242040 136050 242049
rect 73896 242014 73948 242020
rect 70306 241975 70362 241984
rect 70320 241942 70348 241975
rect 70308 241936 70360 241942
rect 69662 241904 69718 241913
rect 70308 241878 70360 241884
rect 69662 241839 69718 241848
rect 68816 241590 68968 241618
rect 69368 241590 69520 241618
rect 68940 240106 68968 241590
rect 69020 240168 69072 240174
rect 69020 240110 69072 240116
rect 68928 240100 68980 240106
rect 68928 240042 68980 240048
rect 67822 237144 67878 237153
rect 67822 237079 67878 237088
rect 67732 215280 67784 215286
rect 67732 215222 67784 215228
rect 69032 207670 69060 240110
rect 69492 238882 69520 241590
rect 69480 238876 69532 238882
rect 69480 238818 69532 238824
rect 69676 225865 69704 241839
rect 69768 241590 70104 241618
rect 70412 241590 70840 241618
rect 71576 241590 71728 241618
rect 72312 241590 72648 241618
rect 73048 241590 73108 241618
rect 69768 240174 69796 241590
rect 69756 240168 69808 240174
rect 69756 240110 69808 240116
rect 69662 225856 69718 225865
rect 69662 225791 69718 225800
rect 70412 224942 70440 241590
rect 71412 240100 71464 240106
rect 71412 240042 71464 240048
rect 71424 238649 71452 240042
rect 71700 239698 71728 241590
rect 72422 239864 72478 239873
rect 72422 239799 72478 239808
rect 71688 239692 71740 239698
rect 71688 239634 71740 239640
rect 71410 238640 71466 238649
rect 71410 238575 71466 238584
rect 70490 228440 70546 228449
rect 70490 228375 70546 228384
rect 70400 224936 70452 224942
rect 70400 224878 70452 224884
rect 69020 207664 69072 207670
rect 69020 207606 69072 207612
rect 67638 205592 67694 205601
rect 67638 205527 67694 205536
rect 70504 176730 70532 228375
rect 72436 192506 72464 239799
rect 72620 239465 72648 241590
rect 72606 239456 72662 239465
rect 72606 239391 72662 239400
rect 72516 237584 72568 237590
rect 72516 237526 72568 237532
rect 72528 222154 72556 237526
rect 72516 222148 72568 222154
rect 72516 222090 72568 222096
rect 73080 197985 73108 241590
rect 73172 241590 73784 241618
rect 73066 197976 73122 197985
rect 73066 197911 73122 197920
rect 72424 192500 72476 192506
rect 72424 192442 72476 192448
rect 73172 191826 73200 241590
rect 73804 239692 73856 239698
rect 73804 239634 73856 239640
rect 73816 204241 73844 239634
rect 73908 215218 73936 242014
rect 135364 241998 135994 242026
rect 76380 241936 76432 241942
rect 76380 241878 76432 241884
rect 74520 241590 74856 241618
rect 75072 241590 75408 241618
rect 74724 240780 74776 240786
rect 74724 240722 74776 240728
rect 74736 236609 74764 240722
rect 74828 240038 74856 241590
rect 75182 240136 75238 240145
rect 75182 240071 75238 240080
rect 74816 240032 74868 240038
rect 74816 239974 74868 239980
rect 74722 236600 74778 236609
rect 74722 236535 74778 236544
rect 73896 215212 73948 215218
rect 73896 215154 73948 215160
rect 73802 204232 73858 204241
rect 73802 204167 73858 204176
rect 75196 200025 75224 240071
rect 75380 239698 75408 241590
rect 75472 241590 75808 241618
rect 75472 240145 75500 241590
rect 76392 241346 76420 241878
rect 76544 241590 77064 241618
rect 77280 241590 77340 241618
rect 76392 241318 76696 241346
rect 75458 240136 75514 240145
rect 75458 240071 75514 240080
rect 76564 240100 76616 240106
rect 76564 240042 76616 240048
rect 75368 239692 75420 239698
rect 75368 239634 75420 239640
rect 75828 239692 75880 239698
rect 75828 239634 75880 239640
rect 75276 238876 75328 238882
rect 75276 238818 75328 238824
rect 75288 209710 75316 238818
rect 75840 228993 75868 239634
rect 76576 238513 76604 240042
rect 76562 238504 76618 238513
rect 76562 238439 76618 238448
rect 75826 228984 75882 228993
rect 75826 228919 75882 228928
rect 75276 209704 75328 209710
rect 75276 209646 75328 209652
rect 76576 201414 76604 238439
rect 76668 211138 76696 241318
rect 77036 238754 77064 241590
rect 77312 240106 77340 241590
rect 77404 241590 78016 241618
rect 78752 241590 79088 241618
rect 79488 241590 79916 241618
rect 80224 241590 80560 241618
rect 80776 241590 81388 241618
rect 81512 241590 81848 241618
rect 82248 241590 82584 241618
rect 77300 240100 77352 240106
rect 77300 240042 77352 240048
rect 77036 238726 77248 238754
rect 77220 223553 77248 238726
rect 77206 223544 77262 223553
rect 77206 223479 77262 223488
rect 77404 212430 77432 241590
rect 79060 239562 79088 241590
rect 79048 239556 79100 239562
rect 79048 239498 79100 239504
rect 77392 212424 77444 212430
rect 77392 212366 77444 212372
rect 76656 211132 76708 211138
rect 76656 211074 76708 211080
rect 76564 201408 76616 201414
rect 76564 201350 76616 201356
rect 75182 200016 75238 200025
rect 75182 199951 75238 199960
rect 79888 195974 79916 241590
rect 79968 239556 80020 239562
rect 79968 239498 80020 239504
rect 79876 195968 79928 195974
rect 79876 195910 79928 195916
rect 79980 192545 80008 239498
rect 80532 239290 80560 241590
rect 80520 239284 80572 239290
rect 80520 239226 80572 239232
rect 81256 239284 81308 239290
rect 81256 239226 81308 239232
rect 81268 218822 81296 239226
rect 81256 218816 81308 218822
rect 81256 218758 81308 218764
rect 81360 193866 81388 241590
rect 81820 239426 81848 241590
rect 82556 240786 82584 241590
rect 82970 241369 82998 241604
rect 83108 241590 83720 241618
rect 84456 241590 84792 241618
rect 85192 241590 85528 241618
rect 85928 241590 86080 241618
rect 82956 241360 83012 241369
rect 82956 241295 83012 241304
rect 82544 240780 82596 240786
rect 82544 240722 82596 240728
rect 81808 239420 81860 239426
rect 81808 239362 81860 239368
rect 82728 239420 82780 239426
rect 82728 239362 82780 239368
rect 82740 223582 82768 239362
rect 82728 223576 82780 223582
rect 82728 223518 82780 223524
rect 83108 202162 83136 241590
rect 84106 241224 84162 241233
rect 84106 241159 84162 241168
rect 83464 240032 83516 240038
rect 83464 239974 83516 239980
rect 83476 204950 83504 239974
rect 84120 224913 84148 241159
rect 84764 239426 84792 241590
rect 84842 239456 84898 239465
rect 84752 239420 84804 239426
rect 84842 239391 84898 239400
rect 84752 239362 84804 239368
rect 84856 226001 84884 239391
rect 84842 225992 84898 226001
rect 84842 225927 84898 225936
rect 84106 224904 84162 224913
rect 84106 224839 84162 224848
rect 85500 209137 85528 241590
rect 86052 240106 86080 241590
rect 86144 241590 86480 241618
rect 86972 241590 87216 241618
rect 87952 241590 88288 241618
rect 88688 241590 89024 241618
rect 89424 241590 89576 241618
rect 90160 241590 90496 241618
rect 90896 241590 91048 241618
rect 91632 241590 91968 241618
rect 92184 241590 92336 241618
rect 92920 241604 93164 241618
rect 86040 240100 86092 240106
rect 86040 240042 86092 240048
rect 86144 238754 86172 241590
rect 86868 240100 86920 240106
rect 86868 240042 86920 240048
rect 85592 238726 86172 238754
rect 85592 229770 85620 238726
rect 85580 229764 85632 229770
rect 85580 229706 85632 229712
rect 85486 209128 85542 209137
rect 85486 209063 85542 209072
rect 83464 204944 83516 204950
rect 83464 204886 83516 204892
rect 83096 202156 83148 202162
rect 83096 202098 83148 202104
rect 86880 200802 86908 240042
rect 86972 217841 87000 241590
rect 86958 217832 87014 217841
rect 86958 217767 87014 217776
rect 86868 200796 86920 200802
rect 86868 200738 86920 200744
rect 88260 196625 88288 241590
rect 88996 239834 89024 241590
rect 88984 239828 89036 239834
rect 88984 239770 89036 239776
rect 88246 196616 88302 196625
rect 88246 196551 88302 196560
rect 81348 193860 81400 193866
rect 81348 193802 81400 193808
rect 79966 192536 80022 192545
rect 79966 192471 80022 192480
rect 73160 191820 73212 191826
rect 73160 191762 73212 191768
rect 89548 189786 89576 241590
rect 90468 240106 90496 241590
rect 90456 240100 90508 240106
rect 90456 240042 90508 240048
rect 90916 240100 90968 240106
rect 90916 240042 90968 240048
rect 89628 239828 89680 239834
rect 89628 239770 89680 239776
rect 89536 189780 89588 189786
rect 89536 189722 89588 189728
rect 89640 189038 89668 239770
rect 90928 220153 90956 240042
rect 90914 220144 90970 220153
rect 90914 220079 90970 220088
rect 89628 189032 89680 189038
rect 89628 188974 89680 188980
rect 91020 185609 91048 241590
rect 91940 240106 91968 241590
rect 91928 240100 91980 240106
rect 91928 240042 91980 240048
rect 92308 215937 92336 241590
rect 92906 241590 93164 241604
rect 93656 241590 93716 241618
rect 92906 241466 92934 241590
rect 92894 241460 92946 241466
rect 92894 241402 92946 241408
rect 92388 240100 92440 240106
rect 92388 240042 92440 240048
rect 92294 215928 92350 215937
rect 92294 215863 92350 215872
rect 92400 209681 92428 240042
rect 92386 209672 92442 209681
rect 92386 209607 92442 209616
rect 93136 200122 93164 241590
rect 93688 218657 93716 241590
rect 94378 241369 94406 241604
rect 95128 241590 95188 241618
rect 93858 241360 93914 241369
rect 93858 241295 93914 241304
rect 94364 241360 94420 241369
rect 94364 241295 94420 241304
rect 93872 222194 93900 241295
rect 93780 222166 93900 222194
rect 93780 220862 93808 222166
rect 93768 220856 93820 220862
rect 93768 220798 93820 220804
rect 93674 218648 93730 218657
rect 93674 218583 93730 218592
rect 93124 200116 93176 200122
rect 93124 200058 93176 200064
rect 93780 191729 93808 220798
rect 93766 191720 93822 191729
rect 93766 191655 93822 191664
rect 95160 189689 95188 241590
rect 95252 241590 95864 241618
rect 96600 241590 96660 241618
rect 97336 241590 97764 241618
rect 97888 241590 97948 241618
rect 98624 241590 99052 241618
rect 99360 241590 99420 241618
rect 95252 205630 95280 241590
rect 96632 238746 96660 241590
rect 97736 238754 97764 241590
rect 96620 238740 96672 238746
rect 97736 238726 97856 238754
rect 96620 238682 96672 238688
rect 95240 205624 95292 205630
rect 95240 205566 95292 205572
rect 97828 198626 97856 238726
rect 97816 198620 97868 198626
rect 97816 198562 97868 198568
rect 95146 189680 95202 189689
rect 95146 189615 95202 189624
rect 91006 185600 91062 185609
rect 91006 185535 91062 185544
rect 97920 183025 97948 241590
rect 99024 238754 99052 241590
rect 99392 240106 99420 241590
rect 99484 241590 100096 241618
rect 100832 241590 101168 241618
rect 101568 241590 101996 241618
rect 99380 240100 99432 240106
rect 99380 240042 99432 240048
rect 99024 238726 99328 238754
rect 99300 188329 99328 238726
rect 99484 206922 99512 241590
rect 100668 240100 100720 240106
rect 100668 240042 100720 240048
rect 100680 207641 100708 240042
rect 101140 239698 101168 241590
rect 101128 239692 101180 239698
rect 101128 239634 101180 239640
rect 101968 221513 101996 241590
rect 102152 241590 102304 241618
rect 103040 241590 103468 241618
rect 102048 239692 102100 239698
rect 102048 239634 102100 239640
rect 101954 221504 102010 221513
rect 101954 221439 102010 221448
rect 102060 212401 102088 239634
rect 102152 231878 102180 241590
rect 102140 231872 102192 231878
rect 102140 231814 102192 231820
rect 102152 231713 102180 231814
rect 102138 231704 102194 231713
rect 102138 231639 102194 231648
rect 102046 212392 102102 212401
rect 102046 212327 102102 212336
rect 100666 207632 100722 207641
rect 100666 207567 100722 207576
rect 99472 206916 99524 206922
rect 99472 206858 99524 206864
rect 103440 191049 103468 241590
rect 103532 241590 103592 241618
rect 104328 241590 104848 241618
rect 103532 233209 103560 241590
rect 103518 233200 103574 233209
rect 103518 233135 103574 233144
rect 104164 231872 104216 231878
rect 104164 231814 104216 231820
rect 104176 193225 104204 231814
rect 104820 217326 104848 241590
rect 104912 241590 105064 241618
rect 105800 241590 106136 241618
rect 106536 241590 106872 241618
rect 107272 241590 107516 241618
rect 104808 217320 104860 217326
rect 104808 217262 104860 217268
rect 104912 211070 104940 241590
rect 106108 240854 106136 241590
rect 106096 240848 106148 240854
rect 106096 240790 106148 240796
rect 106844 239970 106872 241590
rect 106832 239964 106884 239970
rect 106832 239906 106884 239912
rect 106740 232552 106792 232558
rect 106740 232494 106792 232500
rect 106752 231713 106780 232494
rect 106738 231704 106794 231713
rect 106738 231639 106794 231648
rect 106924 228404 106976 228410
rect 106924 228346 106976 228352
rect 104900 211064 104952 211070
rect 104900 211006 104952 211012
rect 106936 195906 106964 228346
rect 107488 220726 107516 241590
rect 107672 241590 108008 241618
rect 108744 241590 108988 241618
rect 109296 241590 109632 241618
rect 110032 241590 110276 241618
rect 110768 241590 111104 241618
rect 111504 241590 111748 241618
rect 107568 239964 107620 239970
rect 107568 239906 107620 239912
rect 107476 220720 107528 220726
rect 107476 220662 107528 220668
rect 106924 195900 106976 195906
rect 106924 195842 106976 195848
rect 107580 193905 107608 239906
rect 107672 238678 107700 241590
rect 107660 238672 107712 238678
rect 107660 238614 107712 238620
rect 108304 238060 108356 238066
rect 108304 238002 108356 238008
rect 108316 233170 108344 238002
rect 108304 233164 108356 233170
rect 108304 233106 108356 233112
rect 108960 227225 108988 241590
rect 109604 239290 109632 241590
rect 109592 239284 109644 239290
rect 109592 239226 109644 239232
rect 108946 227216 109002 227225
rect 108946 227151 109002 227160
rect 110248 224874 110276 241590
rect 111076 239970 111104 241590
rect 111064 239964 111116 239970
rect 111064 239906 111116 239912
rect 111616 239964 111668 239970
rect 111616 239906 111668 239912
rect 110328 239284 110380 239290
rect 110328 239226 110380 239232
rect 110236 224868 110288 224874
rect 110236 224810 110288 224816
rect 110340 217977 110368 239226
rect 110326 217968 110382 217977
rect 110326 217903 110382 217912
rect 111628 203561 111656 239906
rect 111614 203552 111670 203561
rect 111614 203487 111670 203496
rect 111720 200705 111748 241590
rect 111812 241590 112240 241618
rect 112976 241590 113128 241618
rect 113712 241590 114232 241618
rect 114448 241590 114508 241618
rect 115000 241590 115336 241618
rect 115736 241590 115796 241618
rect 111812 215966 111840 241590
rect 111800 215960 111852 215966
rect 111800 215902 111852 215908
rect 113100 208350 113128 241590
rect 114204 238754 114232 241590
rect 114204 238726 114416 238754
rect 114388 231742 114416 238726
rect 114376 231736 114428 231742
rect 114376 231678 114428 231684
rect 114480 219337 114508 241590
rect 115308 240106 115336 241590
rect 115296 240100 115348 240106
rect 115296 240042 115348 240048
rect 115202 232656 115258 232665
rect 115202 232591 115258 232600
rect 115216 222193 115244 232591
rect 115202 222184 115258 222193
rect 115202 222119 115258 222128
rect 114466 219328 114522 219337
rect 114466 219263 114522 219272
rect 113088 208344 113140 208350
rect 113088 208286 113140 208292
rect 115768 202745 115796 241590
rect 116044 241590 116472 241618
rect 116872 241590 117208 241618
rect 117944 241590 118464 241618
rect 115940 240168 115992 240174
rect 115940 240110 115992 240116
rect 115848 240100 115900 240106
rect 115848 240042 115900 240048
rect 115754 202736 115810 202745
rect 115754 202671 115810 202680
rect 111706 200696 111762 200705
rect 111706 200631 111762 200640
rect 107566 193896 107622 193905
rect 107566 193831 107622 193840
rect 104162 193216 104218 193225
rect 104162 193151 104218 193160
rect 103426 191040 103482 191049
rect 103426 190975 103482 190984
rect 113088 189100 113140 189106
rect 113088 189042 113140 189048
rect 99286 188320 99342 188329
rect 99286 188255 99342 188264
rect 106188 185020 106240 185026
rect 106188 184962 106240 184968
rect 100668 183660 100720 183666
rect 100668 183602 100720 183608
rect 97906 183016 97962 183025
rect 97906 182951 97962 182960
rect 98918 182200 98974 182209
rect 98918 182135 98974 182144
rect 98932 177585 98960 182135
rect 98918 177576 98974 177585
rect 98918 177511 98974 177520
rect 100680 176769 100708 183602
rect 102048 182232 102100 182238
rect 102048 182174 102100 182180
rect 100758 179480 100814 179489
rect 100758 179415 100814 179424
rect 100772 176905 100800 179415
rect 102060 177585 102088 182174
rect 106200 177585 106228 184962
rect 108948 183592 109000 183598
rect 108948 183534 109000 183540
rect 108960 177585 108988 183534
rect 113100 177585 113128 189042
rect 115860 187649 115888 240042
rect 115952 237386 115980 240110
rect 115940 237380 115992 237386
rect 115940 237322 115992 237328
rect 116044 235657 116072 241590
rect 116584 240780 116636 240786
rect 116584 240722 116636 240728
rect 116030 235648 116086 235657
rect 116030 235583 116086 235592
rect 116596 226302 116624 240722
rect 116872 240174 116900 241590
rect 116860 240168 116912 240174
rect 116860 240110 116912 240116
rect 118436 238754 118464 241590
rect 118666 241369 118694 241604
rect 118896 241590 119416 241618
rect 120152 241590 120488 241618
rect 120704 241590 121040 241618
rect 121440 241590 121776 241618
rect 122176 241590 122696 241618
rect 118652 241360 118708 241369
rect 118652 241295 118708 241304
rect 118436 238726 118648 238754
rect 116584 226296 116636 226302
rect 116584 226238 116636 226244
rect 118620 199442 118648 238726
rect 118896 235890 118924 241590
rect 120460 240106 120488 241590
rect 120724 240168 120776 240174
rect 120724 240110 120776 240116
rect 120448 240100 120500 240106
rect 120448 240042 120500 240048
rect 120736 237318 120764 240110
rect 121012 239970 121040 241590
rect 121748 240106 121776 241590
rect 121368 240100 121420 240106
rect 121368 240042 121420 240048
rect 121736 240100 121788 240106
rect 121736 240042 121788 240048
rect 121000 239964 121052 239970
rect 121000 239906 121052 239912
rect 120724 237312 120776 237318
rect 120724 237254 120776 237260
rect 118884 235884 118936 235890
rect 118884 235826 118936 235832
rect 118896 234666 118924 235826
rect 118884 234660 118936 234666
rect 118884 234602 118936 234608
rect 119344 234660 119396 234666
rect 119344 234602 119396 234608
rect 119356 223417 119384 234602
rect 119342 223408 119398 223417
rect 119342 223343 119398 223352
rect 121380 202881 121408 240042
rect 122102 233880 122158 233889
rect 122102 233815 122158 233824
rect 122116 228857 122144 233815
rect 122102 228848 122158 228857
rect 122102 228783 122158 228792
rect 122668 215257 122696 241590
rect 122852 241590 122912 241618
rect 123036 241590 123648 241618
rect 124384 241590 124720 241618
rect 125120 241590 125548 241618
rect 125856 241590 126192 241618
rect 126408 241590 126928 241618
rect 127144 241590 127480 241618
rect 122748 240100 122800 240106
rect 122748 240042 122800 240048
rect 122654 215248 122710 215257
rect 122654 215183 122710 215192
rect 122760 204921 122788 240042
rect 122852 212498 122880 241590
rect 122932 239964 122984 239970
rect 122932 239906 122984 239912
rect 122944 238513 122972 239906
rect 122930 238504 122986 238513
rect 122930 238439 122986 238448
rect 123036 234530 123064 241590
rect 124692 240106 124720 241590
rect 124864 240848 124916 240854
rect 124864 240790 124916 240796
rect 124680 240100 124732 240106
rect 124680 240042 124732 240048
rect 124128 235272 124180 235278
rect 124128 235214 124180 235220
rect 123024 234524 123076 234530
rect 123024 234466 123076 234472
rect 122840 212492 122892 212498
rect 122840 212434 122892 212440
rect 124140 206961 124168 235214
rect 124876 231810 124904 240790
rect 125416 240100 125468 240106
rect 125416 240042 125468 240048
rect 125322 233336 125378 233345
rect 125322 233271 125378 233280
rect 124864 231804 124916 231810
rect 124864 231746 124916 231752
rect 125336 231674 125364 233271
rect 125324 231668 125376 231674
rect 125324 231610 125376 231616
rect 125428 228410 125456 240042
rect 125416 228404 125468 228410
rect 125416 228346 125468 228352
rect 124126 206952 124182 206961
rect 124126 206887 124182 206896
rect 122746 204912 122802 204921
rect 122746 204847 122802 204856
rect 121366 202872 121422 202881
rect 124140 202842 124168 206887
rect 125520 202842 125548 241590
rect 126164 239737 126192 241590
rect 126150 239728 126206 239737
rect 126150 239663 126206 239672
rect 126900 213761 126928 241590
rect 126980 240100 127032 240106
rect 126980 240042 127032 240048
rect 126992 233238 127020 240042
rect 127452 240038 127480 241590
rect 127544 241590 127880 241618
rect 128616 241590 128952 241618
rect 129352 241590 129596 241618
rect 130088 241590 130424 241618
rect 130824 241590 131068 241618
rect 131560 241590 131896 241618
rect 132112 241590 132356 241618
rect 132848 241590 133184 241618
rect 133584 241590 133736 241618
rect 134320 241590 134656 241618
rect 127544 240106 127572 241590
rect 127532 240100 127584 240106
rect 127532 240042 127584 240048
rect 127440 240032 127492 240038
rect 127440 239974 127492 239980
rect 128268 240032 128320 240038
rect 128268 239974 128320 239980
rect 126980 233232 127032 233238
rect 126980 233174 127032 233180
rect 126886 213752 126942 213761
rect 126886 213687 126942 213696
rect 121366 202807 121422 202816
rect 124128 202836 124180 202842
rect 124128 202778 124180 202784
rect 125508 202836 125560 202842
rect 125508 202778 125560 202784
rect 118608 199436 118660 199442
rect 118608 199378 118660 199384
rect 128280 195945 128308 239974
rect 128924 239290 128952 241590
rect 128912 239284 128964 239290
rect 128912 239226 128964 239232
rect 129568 230353 129596 241590
rect 130396 240106 130424 241590
rect 130384 240100 130436 240106
rect 130384 240042 130436 240048
rect 130936 240100 130988 240106
rect 130936 240042 130988 240048
rect 129648 239284 129700 239290
rect 129648 239226 129700 239232
rect 129554 230344 129610 230353
rect 129554 230279 129610 230288
rect 128360 218816 128412 218822
rect 128360 218758 128412 218764
rect 128372 211041 128400 218758
rect 128358 211032 128414 211041
rect 128358 210967 128414 210976
rect 129660 202201 129688 239226
rect 130948 219434 130976 240042
rect 130936 219428 130988 219434
rect 130936 219370 130988 219376
rect 131040 216646 131068 241590
rect 131868 240106 131896 241590
rect 131856 240100 131908 240106
rect 131856 240042 131908 240048
rect 131028 216640 131080 216646
rect 131028 216582 131080 216588
rect 132328 214577 132356 241590
rect 132408 240100 132460 240106
rect 132408 240042 132460 240048
rect 132314 214568 132370 214577
rect 132314 214503 132370 214512
rect 132420 209778 132448 240042
rect 133156 239970 133184 241590
rect 133144 239964 133196 239970
rect 133144 239906 133196 239912
rect 133512 231736 133564 231742
rect 133512 231678 133564 231684
rect 133602 231704 133658 231713
rect 133524 231441 133552 231678
rect 133602 231639 133658 231648
rect 133510 231432 133566 231441
rect 133510 231367 133566 231376
rect 133616 230518 133644 231639
rect 133604 230512 133656 230518
rect 133604 230454 133656 230460
rect 132408 209772 132460 209778
rect 132408 209714 132460 209720
rect 133708 207777 133736 241590
rect 134628 240106 134656 241590
rect 134720 241590 135056 241618
rect 134616 240100 134668 240106
rect 134616 240042 134668 240048
rect 133788 239964 133840 239970
rect 133788 239906 133840 239912
rect 133694 207768 133750 207777
rect 133694 207703 133750 207712
rect 129646 202192 129702 202201
rect 129646 202127 129702 202136
rect 133800 198121 133828 239906
rect 134720 238754 134748 241590
rect 135168 240100 135220 240106
rect 135168 240042 135220 240048
rect 133892 238726 134748 238754
rect 133892 221474 133920 238726
rect 135180 227361 135208 240042
rect 135364 235278 135392 241998
rect 135994 241975 136050 241984
rect 136914 242040 136970 242049
rect 138202 242040 138258 242049
rect 136970 241998 137264 242026
rect 136914 241975 136970 241984
rect 146758 242040 146814 242049
rect 138258 241998 138888 242026
rect 146464 241998 146758 242026
rect 138202 241975 138258 241984
rect 136528 241590 136588 241618
rect 136088 240168 136140 240174
rect 136088 240110 136140 240116
rect 136100 237318 136128 240110
rect 136088 237312 136140 237318
rect 136088 237254 136140 237260
rect 135352 235272 135404 235278
rect 135352 235214 135404 235220
rect 135166 227352 135222 227361
rect 135166 227287 135222 227296
rect 134524 227044 134576 227050
rect 134524 226986 134576 226992
rect 133880 221468 133932 221474
rect 133880 221410 133932 221416
rect 134536 213246 134564 226986
rect 136560 220697 136588 241590
rect 136928 238754 136956 241975
rect 137816 241590 137968 241618
rect 136744 238726 136956 238754
rect 136744 237289 136772 238726
rect 136730 237280 136786 237289
rect 136730 237215 136786 237224
rect 136744 236065 136772 237215
rect 136730 236056 136786 236065
rect 136730 235991 136786 236000
rect 137282 236056 137338 236065
rect 137282 235991 137338 236000
rect 137296 224641 137324 235991
rect 137282 224632 137338 224641
rect 137282 224567 137338 224576
rect 136546 220688 136602 220697
rect 136546 220623 136602 220632
rect 134524 213240 134576 213246
rect 134524 213182 134576 213188
rect 137940 204270 137968 241590
rect 138860 240786 138888 241998
rect 150072 242014 150124 242020
rect 146758 241975 146814 241984
rect 138952 241590 139288 241618
rect 140024 241590 140544 241618
rect 140760 241590 141096 241618
rect 141496 241590 141832 241618
rect 142232 241590 142292 241618
rect 138848 240780 138900 240786
rect 138848 240722 138900 240728
rect 138952 240106 138980 241590
rect 138020 240100 138072 240106
rect 138020 240042 138072 240048
rect 138940 240100 138992 240106
rect 138940 240042 138992 240048
rect 138032 235890 138060 240042
rect 140516 238754 140544 241590
rect 141068 239562 141096 241590
rect 141804 239873 141832 241590
rect 142264 239970 142292 241590
rect 142356 241590 142968 241618
rect 143704 241590 144040 241618
rect 142252 239964 142304 239970
rect 142252 239906 142304 239912
rect 141790 239864 141846 239873
rect 141790 239799 141846 239808
rect 141056 239556 141108 239562
rect 141056 239498 141108 239504
rect 142068 239556 142120 239562
rect 142068 239498 142120 239504
rect 140516 238726 140728 238754
rect 138020 235884 138072 235890
rect 138020 235826 138072 235832
rect 138662 233064 138718 233073
rect 138662 232999 138718 233008
rect 137928 204264 137980 204270
rect 137928 204206 137980 204212
rect 138676 202745 138704 232999
rect 140042 229800 140098 229809
rect 140042 229735 140098 229744
rect 138662 202736 138718 202745
rect 138662 202671 138718 202680
rect 133786 198112 133842 198121
rect 133786 198047 133842 198056
rect 138676 197305 138704 202671
rect 140056 201385 140084 229735
rect 140700 209001 140728 238726
rect 140778 233336 140834 233345
rect 140778 233271 140834 233280
rect 140792 231577 140820 233271
rect 140778 231568 140834 231577
rect 140778 231503 140834 231512
rect 142080 230450 142108 239498
rect 142356 234433 142384 241590
rect 144012 240106 144040 241590
rect 144242 241466 144270 241604
rect 144932 241590 144992 241618
rect 145728 241590 146248 241618
rect 147200 241590 147628 241618
rect 147936 241590 148272 241618
rect 148672 241590 148916 241618
rect 149408 241590 149560 241618
rect 144230 241460 144282 241466
rect 144230 241402 144282 241408
rect 144000 240100 144052 240106
rect 144000 240042 144052 240048
rect 144828 240100 144880 240106
rect 144828 240042 144880 240048
rect 143448 239964 143500 239970
rect 143448 239906 143500 239912
rect 142342 234424 142398 234433
rect 142342 234359 142398 234368
rect 142068 230444 142120 230450
rect 142068 230386 142120 230392
rect 142804 216708 142856 216714
rect 142804 216650 142856 216656
rect 142816 209710 142844 216650
rect 142804 209704 142856 209710
rect 142804 209646 142856 209652
rect 140686 208992 140742 209001
rect 140686 208927 140742 208936
rect 140042 201376 140098 201385
rect 140042 201311 140098 201320
rect 138662 197296 138718 197305
rect 143460 197266 143488 239906
rect 144840 230382 144868 240042
rect 144932 233073 144960 241590
rect 144918 233064 144974 233073
rect 144918 232999 144974 233008
rect 146116 230512 146168 230518
rect 146116 230454 146168 230460
rect 144828 230376 144880 230382
rect 144828 230318 144880 230324
rect 144184 229764 144236 229770
rect 144184 229706 144236 229712
rect 144196 209098 144224 229706
rect 146128 229090 146156 230454
rect 146116 229084 146168 229090
rect 146116 229026 146168 229032
rect 144184 209092 144236 209098
rect 144184 209034 144236 209040
rect 146220 203590 146248 241590
rect 147600 231742 147628 241590
rect 147680 240780 147732 240786
rect 147680 240722 147732 240728
rect 147692 240106 147720 240722
rect 147680 240100 147732 240106
rect 147680 240042 147732 240048
rect 148244 239834 148272 241590
rect 148232 239828 148284 239834
rect 148232 239770 148284 239776
rect 147588 231736 147640 231742
rect 147588 231678 147640 231684
rect 148324 230376 148376 230382
rect 148324 230318 148376 230324
rect 148336 220794 148364 230318
rect 148888 229770 148916 241590
rect 149532 240786 149560 241590
rect 149624 241590 149960 241618
rect 149520 240780 149572 240786
rect 149520 240722 149572 240728
rect 148968 239828 149020 239834
rect 148968 239770 149020 239776
rect 148876 229764 148928 229770
rect 148876 229706 148928 229712
rect 148324 220788 148376 220794
rect 148324 220730 148376 220736
rect 147678 214024 147734 214033
rect 147678 213959 147734 213968
rect 147692 212430 147720 213959
rect 147680 212424 147732 212430
rect 147680 212366 147732 212372
rect 148980 211818 149008 239770
rect 149624 239630 149652 241590
rect 149060 239624 149112 239630
rect 149060 239566 149112 239572
rect 149612 239624 149664 239630
rect 149612 239566 149664 239572
rect 149072 237289 149100 239566
rect 150084 238754 150112 242014
rect 154026 241768 154082 241777
rect 154026 241703 154082 241712
rect 149716 238726 150112 238754
rect 150544 241590 150696 241618
rect 151432 241590 151768 241618
rect 149716 237318 149744 238726
rect 149704 237312 149756 237318
rect 149058 237280 149114 237289
rect 149704 237254 149756 237260
rect 149058 237215 149114 237224
rect 150544 235793 150572 241590
rect 150530 235784 150586 235793
rect 150530 235719 150586 235728
rect 151174 233880 151230 233889
rect 151174 233815 151230 233824
rect 151082 232520 151138 232529
rect 151082 232455 151138 232464
rect 151096 227730 151124 232455
rect 151188 228857 151216 233815
rect 151174 228848 151230 228857
rect 151174 228783 151230 228792
rect 151084 227724 151136 227730
rect 151084 227666 151136 227672
rect 151084 225616 151136 225622
rect 151084 225558 151136 225564
rect 151096 215218 151124 225558
rect 151084 215212 151136 215218
rect 151084 215154 151136 215160
rect 148968 211812 149020 211818
rect 148968 211754 149020 211760
rect 146208 203584 146260 203590
rect 146208 203526 146260 203532
rect 138662 197231 138718 197240
rect 143448 197260 143500 197266
rect 143448 197202 143500 197208
rect 128266 195936 128322 195945
rect 128266 195871 128322 195880
rect 151740 195265 151768 241590
rect 151924 241590 152168 241618
rect 152904 241590 153148 241618
rect 153640 241590 153976 241618
rect 151924 237318 151952 241590
rect 152464 240848 152516 240854
rect 152464 240790 152516 240796
rect 151912 237312 151964 237318
rect 151912 237254 151964 237260
rect 152476 226001 152504 240790
rect 152462 225992 152518 226001
rect 152462 225927 152518 225936
rect 153120 210905 153148 241590
rect 153948 239290 153976 241590
rect 153936 239284 153988 239290
rect 153936 239226 153988 239232
rect 154040 238754 154068 241703
rect 154376 241590 154436 241618
rect 153856 238726 154068 238754
rect 153856 234598 153884 238726
rect 153844 234592 153896 234598
rect 153844 234534 153896 234540
rect 153106 210896 153162 210905
rect 153106 210831 153162 210840
rect 154408 205057 154436 241590
rect 154868 241505 154896 245618
rect 155316 244384 155368 244390
rect 155316 244326 155368 244332
rect 155222 242992 155278 243001
rect 155222 242927 155278 242936
rect 154854 241496 154910 241505
rect 154854 241431 154910 241440
rect 154488 239284 154540 239290
rect 154488 239226 154540 239232
rect 154394 205048 154450 205057
rect 154394 204983 154450 204992
rect 154500 202337 154528 239226
rect 155236 222902 155264 242927
rect 155328 227662 155356 244326
rect 155880 243438 155908 264143
rect 156418 259040 156474 259049
rect 156418 258975 156474 258984
rect 156432 258126 156460 258975
rect 156420 258120 156472 258126
rect 156420 258062 156472 258068
rect 156420 253632 156472 253638
rect 156418 253600 156420 253609
rect 156472 253600 156474 253609
rect 156418 253535 156474 253544
rect 156418 249520 156474 249529
rect 156418 249455 156474 249464
rect 156432 248470 156460 249455
rect 156420 248464 156472 248470
rect 156420 248406 156472 248412
rect 156050 244080 156106 244089
rect 156050 244015 156106 244024
rect 155408 243432 155460 243438
rect 155408 243374 155460 243380
rect 155868 243432 155920 243438
rect 155868 243374 155920 243380
rect 155420 235890 155448 243374
rect 155880 243030 155908 243374
rect 155868 243024 155920 243030
rect 155868 242966 155920 242972
rect 156064 242962 156092 244015
rect 156052 242956 156104 242962
rect 156052 242898 156104 242904
rect 155408 235884 155460 235890
rect 155408 235826 155460 235832
rect 155684 235816 155736 235822
rect 155684 235758 155736 235764
rect 155696 235657 155724 235758
rect 155682 235648 155738 235657
rect 155682 235583 155738 235592
rect 155316 227656 155368 227662
rect 155316 227598 155368 227604
rect 156616 227497 156644 318543
rect 156708 303657 156736 353903
rect 157246 319968 157302 319977
rect 157246 319903 157302 319912
rect 157260 319530 157288 319903
rect 157248 319524 157300 319530
rect 157248 319466 157300 319472
rect 157246 318880 157302 318889
rect 157246 318815 157248 318824
rect 157300 318815 157302 318824
rect 157248 318786 157300 318792
rect 157246 316976 157302 316985
rect 157352 316962 157380 364919
rect 157302 316934 157380 316962
rect 157246 316911 157302 316920
rect 157260 316810 157288 316911
rect 157248 316804 157300 316810
rect 157248 316746 157300 316752
rect 157246 315888 157302 315897
rect 157302 315846 157380 315874
rect 157246 315823 157302 315832
rect 157246 312624 157302 312633
rect 157352 312594 157380 315846
rect 157246 312559 157302 312568
rect 157340 312588 157392 312594
rect 157260 311914 157288 312559
rect 157340 312530 157392 312536
rect 157248 311908 157300 311914
rect 157248 311850 157300 311856
rect 157246 311536 157302 311545
rect 157246 311471 157302 311480
rect 157260 310554 157288 311471
rect 157248 310548 157300 310554
rect 157248 310490 157300 310496
rect 157246 310448 157302 310457
rect 157246 310383 157302 310392
rect 157154 309632 157210 309641
rect 157154 309567 157210 309576
rect 157168 308417 157196 309567
rect 157260 309233 157288 310383
rect 157246 309224 157302 309233
rect 157246 309159 157302 309168
rect 157154 308408 157210 308417
rect 157154 308343 157210 308352
rect 157246 306368 157302 306377
rect 157246 306303 157248 306312
rect 157300 306303 157302 306312
rect 157248 306274 157300 306280
rect 157246 305280 157302 305289
rect 157246 305215 157248 305224
rect 157300 305215 157302 305224
rect 157248 305186 157300 305192
rect 156694 303648 156750 303657
rect 156694 303583 156750 303592
rect 156708 296857 156736 303583
rect 157246 303104 157302 303113
rect 157246 303039 157302 303048
rect 157260 302258 157288 303039
rect 157248 302252 157300 302258
rect 157248 302194 157300 302200
rect 156786 302016 156842 302025
rect 156786 301951 156842 301960
rect 156800 300898 156828 301951
rect 156788 300892 156840 300898
rect 156788 300834 156840 300840
rect 157154 300112 157210 300121
rect 157154 300047 157210 300056
rect 157168 299538 157196 300047
rect 157156 299532 157208 299538
rect 157156 299474 157208 299480
rect 157248 299464 157300 299470
rect 157248 299406 157300 299412
rect 157260 299033 157288 299406
rect 157246 299024 157302 299033
rect 157246 298959 157302 298968
rect 156694 296848 156750 296857
rect 156694 296783 156750 296792
rect 157246 292768 157302 292777
rect 157522 292768 157578 292777
rect 157246 292703 157302 292712
rect 157352 292726 157522 292754
rect 157260 292602 157288 292703
rect 157248 292596 157300 292602
rect 157248 292538 157300 292544
rect 157352 292482 157380 292726
rect 157522 292703 157578 292712
rect 157260 292454 157380 292482
rect 156786 291680 156842 291689
rect 156786 291615 156842 291624
rect 156800 291242 156828 291615
rect 156788 291236 156840 291242
rect 156788 291178 156840 291184
rect 156694 291136 156750 291145
rect 156694 291071 156750 291080
rect 156708 290193 156736 291071
rect 157260 290601 157288 292454
rect 157246 290592 157302 290601
rect 157246 290527 157302 290536
rect 156694 290184 156750 290193
rect 156694 290119 156750 290128
rect 156708 288266 156736 290119
rect 156786 289504 156842 289513
rect 156786 289439 156842 289448
rect 156800 288454 156828 289439
rect 156788 288448 156840 288454
rect 156788 288390 156840 288396
rect 156708 288238 156828 288266
rect 156694 287328 156750 287337
rect 156694 287263 156750 287272
rect 156708 275233 156736 287263
rect 156694 275224 156750 275233
rect 156694 275159 156750 275168
rect 156694 259856 156750 259865
rect 156694 259791 156750 259800
rect 156602 227488 156658 227497
rect 156602 227423 156658 227432
rect 155224 222896 155276 222902
rect 155224 222838 155276 222844
rect 156616 218754 156644 227423
rect 156604 218748 156656 218754
rect 156604 218690 156656 218696
rect 154486 202328 154542 202337
rect 154486 202263 154542 202272
rect 156708 199345 156736 259791
rect 156800 247353 156828 288238
rect 157246 286240 157302 286249
rect 157246 286175 157302 286184
rect 157260 285734 157288 286175
rect 157248 285728 157300 285734
rect 157248 285670 157300 285676
rect 157248 284368 157300 284374
rect 157246 284336 157248 284345
rect 157300 284336 157302 284345
rect 157246 284271 157302 284280
rect 157246 283248 157302 283257
rect 157246 283183 157302 283192
rect 157260 282946 157288 283183
rect 157248 282940 157300 282946
rect 157248 282882 157300 282888
rect 157156 282872 157208 282878
rect 157156 282814 157208 282820
rect 157168 282169 157196 282814
rect 157154 282160 157210 282169
rect 157154 282095 157210 282104
rect 157248 281512 157300 281518
rect 157248 281454 157300 281460
rect 157260 281081 157288 281454
rect 157246 281072 157302 281081
rect 157246 281007 157302 281016
rect 157064 280832 157116 280838
rect 157064 280774 157116 280780
rect 156970 279984 157026 279993
rect 156970 279919 157026 279928
rect 156984 278866 157012 279919
rect 156972 278860 157024 278866
rect 156972 278802 157024 278808
rect 156878 276720 156934 276729
rect 156878 276655 156934 276664
rect 156892 276078 156920 276655
rect 156880 276072 156932 276078
rect 156880 276014 156932 276020
rect 157076 275913 157104 280774
rect 157248 279064 157300 279070
rect 157248 279006 157300 279012
rect 157260 278905 157288 279006
rect 157246 278896 157302 278905
rect 157246 278831 157302 278840
rect 157246 277808 157302 277817
rect 157246 277743 157302 277752
rect 157260 277438 157288 277743
rect 157248 277432 157300 277438
rect 157248 277374 157300 277380
rect 157062 275904 157118 275913
rect 157062 275839 157118 275848
rect 156878 274816 156934 274825
rect 156878 274751 156934 274760
rect 156892 264246 156920 274751
rect 157154 272640 157210 272649
rect 157154 272575 157210 272584
rect 157168 271182 157196 272575
rect 157246 271552 157302 271561
rect 157246 271487 157302 271496
rect 157156 271176 157208 271182
rect 157156 271118 157208 271124
rect 157260 270570 157288 271487
rect 157248 270564 157300 270570
rect 157248 270506 157300 270512
rect 157246 270464 157302 270473
rect 157246 270399 157302 270408
rect 157260 269142 157288 270399
rect 157248 269136 157300 269142
rect 157248 269078 157300 269084
rect 157248 268388 157300 268394
rect 157248 268330 157300 268336
rect 157260 268297 157288 268330
rect 157246 268288 157302 268297
rect 157246 268223 157302 268232
rect 157248 267708 157300 267714
rect 157248 267650 157300 267656
rect 157260 267481 157288 267650
rect 157246 267472 157302 267481
rect 157246 267407 157302 267416
rect 157248 266348 157300 266354
rect 157248 266290 157300 266296
rect 157260 265305 157288 266290
rect 157246 265296 157302 265305
rect 157246 265231 157302 265240
rect 156880 264240 156932 264246
rect 156880 264182 156932 264188
rect 157246 263120 157302 263129
rect 157246 263055 157302 263064
rect 157260 262274 157288 263055
rect 157248 262268 157300 262274
rect 157248 262210 157300 262216
rect 156880 257984 156932 257990
rect 156878 257952 156880 257961
rect 156932 257952 156934 257961
rect 156878 257887 156934 257896
rect 157246 256864 157302 256873
rect 157246 256799 157248 256808
rect 157300 256799 157302 256808
rect 157248 256770 157300 256776
rect 157246 255776 157302 255785
rect 157246 255711 157302 255720
rect 157260 255338 157288 255711
rect 157248 255332 157300 255338
rect 157248 255274 157300 255280
rect 157246 254688 157302 254697
rect 157246 254623 157302 254632
rect 157260 253978 157288 254623
rect 157248 253972 157300 253978
rect 157248 253914 157300 253920
rect 156880 251388 156932 251394
rect 156880 251330 156932 251336
rect 156786 247344 156842 247353
rect 156786 247279 156842 247288
rect 156788 245744 156840 245750
rect 156788 245686 156840 245692
rect 156800 233170 156828 245686
rect 156892 242185 156920 251330
rect 157246 250608 157302 250617
rect 157246 250543 157302 250552
rect 157260 249830 157288 250543
rect 157248 249824 157300 249830
rect 157248 249766 157300 249772
rect 157156 249756 157208 249762
rect 157156 249698 157208 249704
rect 157168 248441 157196 249698
rect 157154 248432 157210 248441
rect 157154 248367 157210 248376
rect 156970 245168 157026 245177
rect 156970 245103 157026 245112
rect 156984 244322 157012 245103
rect 156972 244316 157024 244322
rect 156972 244258 157024 244264
rect 156878 242176 156934 242185
rect 156878 242111 156934 242120
rect 156878 240816 156934 240825
rect 156878 240751 156934 240760
rect 156788 233164 156840 233170
rect 156788 233106 156840 233112
rect 156892 229090 156920 240751
rect 157996 235249 158024 438126
rect 158076 400920 158128 400926
rect 158076 400862 158128 400868
rect 158088 307873 158116 400862
rect 158720 380180 158772 380186
rect 158720 380122 158772 380128
rect 158168 327208 158220 327214
rect 158168 327150 158220 327156
rect 158180 318102 158208 327150
rect 158168 318096 158220 318102
rect 158168 318038 158220 318044
rect 158074 307864 158130 307873
rect 158074 307799 158130 307808
rect 157982 235240 158038 235249
rect 157982 235175 158038 235184
rect 156880 229084 156932 229090
rect 156880 229026 156932 229032
rect 158088 220726 158116 307799
rect 158732 306338 158760 380122
rect 159364 356040 159416 356046
rect 159364 355982 159416 355988
rect 158812 332716 158864 332722
rect 158812 332658 158864 332664
rect 158824 327758 158852 332658
rect 159376 331226 159404 355982
rect 159546 335472 159602 335481
rect 159546 335407 159602 335416
rect 159364 331220 159416 331226
rect 159364 331162 159416 331168
rect 159456 329928 159508 329934
rect 159456 329870 159508 329876
rect 159362 327856 159418 327865
rect 159362 327791 159418 327800
rect 158812 327752 158864 327758
rect 158812 327694 158864 327700
rect 158720 306332 158772 306338
rect 158720 306274 158772 306280
rect 158732 302938 158760 306274
rect 158720 302932 158772 302938
rect 158720 302874 158772 302880
rect 158626 295352 158682 295361
rect 158626 295287 158682 295296
rect 158168 253224 158220 253230
rect 158168 253166 158220 253172
rect 158180 227225 158208 253166
rect 158640 247722 158668 295287
rect 159376 273329 159404 327791
rect 159468 291145 159496 329870
rect 159560 322153 159588 335407
rect 159546 322144 159602 322153
rect 159546 322079 159602 322088
rect 160112 319530 160140 449958
rect 160744 370524 160796 370530
rect 160744 370466 160796 370472
rect 160190 342544 160246 342553
rect 160190 342479 160246 342488
rect 160204 336025 160232 342479
rect 160190 336016 160246 336025
rect 160190 335951 160246 335960
rect 160100 319524 160152 319530
rect 160100 319466 160152 319472
rect 160008 295384 160060 295390
rect 160008 295326 160060 295332
rect 159640 291236 159692 291242
rect 159640 291178 159692 291184
rect 159454 291136 159510 291145
rect 159454 291071 159510 291080
rect 159546 282160 159602 282169
rect 159546 282095 159602 282104
rect 159456 273964 159508 273970
rect 159456 273906 159508 273912
rect 159362 273320 159418 273329
rect 159362 273255 159418 273264
rect 158720 256760 158772 256766
rect 158720 256702 158772 256708
rect 158732 253638 158760 256702
rect 158720 253632 158772 253638
rect 158720 253574 158772 253580
rect 159364 251932 159416 251938
rect 159364 251874 159416 251880
rect 158628 247716 158680 247722
rect 158628 247658 158680 247664
rect 158718 235240 158774 235249
rect 158718 235175 158774 235184
rect 158166 227216 158222 227225
rect 158166 227151 158222 227160
rect 158076 220720 158128 220726
rect 158076 220662 158128 220668
rect 156694 199336 156750 199345
rect 156694 199271 156750 199280
rect 158732 198626 158760 235175
rect 159376 222154 159404 251874
rect 159468 231742 159496 273906
rect 159560 257990 159588 282095
rect 159652 267034 159680 291178
rect 159640 267028 159692 267034
rect 159640 266970 159692 266976
rect 159548 257984 159600 257990
rect 159548 257926 159600 257932
rect 159548 254584 159600 254590
rect 159548 254526 159600 254532
rect 159560 235822 159588 254526
rect 159548 235816 159600 235822
rect 159548 235758 159600 235764
rect 159456 231736 159508 231742
rect 159456 231678 159508 231684
rect 160020 230353 160048 295326
rect 160100 278860 160152 278866
rect 160100 278802 160152 278808
rect 160112 276690 160140 278802
rect 160100 276684 160152 276690
rect 160100 276626 160152 276632
rect 160006 230344 160062 230353
rect 160006 230279 160062 230288
rect 160756 226370 160784 370466
rect 160928 341012 160980 341018
rect 160928 340954 160980 340960
rect 160836 334076 160888 334082
rect 160836 334018 160888 334024
rect 160848 260166 160876 334018
rect 160940 329118 160968 340954
rect 160928 329112 160980 329118
rect 160928 329054 160980 329060
rect 161020 328500 161072 328506
rect 161020 328442 161072 328448
rect 161032 325038 161060 328442
rect 161020 325032 161072 325038
rect 161020 324974 161072 324980
rect 160926 315072 160982 315081
rect 160926 315007 160982 315016
rect 160940 289105 160968 315007
rect 160926 289096 160982 289105
rect 160926 289031 160982 289040
rect 161492 280154 161520 454038
rect 166264 443692 166316 443698
rect 166264 443634 166316 443640
rect 162860 409896 162912 409902
rect 162860 409838 162912 409844
rect 162768 403640 162820 403646
rect 162768 403582 162820 403588
rect 162780 403034 162808 403582
rect 161572 403028 161624 403034
rect 161572 402970 161624 402976
rect 162768 403028 162820 403034
rect 162768 402970 162820 402976
rect 161584 295390 161612 402970
rect 162124 346520 162176 346526
rect 162124 346462 162176 346468
rect 161756 331220 161808 331226
rect 161756 331162 161808 331168
rect 161768 326398 161796 331162
rect 162136 330546 162164 346462
rect 162306 335744 162362 335753
rect 162306 335679 162362 335688
rect 162124 330540 162176 330546
rect 162124 330482 162176 330488
rect 162216 326936 162268 326942
rect 162216 326878 162268 326884
rect 161756 326392 161808 326398
rect 161756 326334 161808 326340
rect 162124 318844 162176 318850
rect 162124 318786 162176 318792
rect 162136 305658 162164 318786
rect 162124 305652 162176 305658
rect 162124 305594 162176 305600
rect 162122 295488 162178 295497
rect 162122 295423 162178 295432
rect 161572 295384 161624 295390
rect 161572 295326 161624 295332
rect 161400 280126 161520 280154
rect 161400 279070 161428 280126
rect 161388 279064 161440 279070
rect 161388 279006 161440 279012
rect 160928 261588 160980 261594
rect 160928 261530 160980 261536
rect 160836 260160 160888 260166
rect 160836 260102 160888 260108
rect 160836 244316 160888 244322
rect 160836 244258 160888 244264
rect 160744 226364 160796 226370
rect 160744 226306 160796 226312
rect 159364 222148 159416 222154
rect 159364 222090 159416 222096
rect 158720 198620 158772 198626
rect 158720 198562 158772 198568
rect 160756 195945 160784 226306
rect 160742 195936 160798 195945
rect 160742 195871 160798 195880
rect 151726 195256 151782 195265
rect 151726 195191 151782 195200
rect 133788 190528 133840 190534
rect 133788 190470 133840 190476
rect 131028 187740 131080 187746
rect 131028 187682 131080 187688
rect 115846 187640 115902 187649
rect 115846 187575 115902 187584
rect 128268 186380 128320 186386
rect 128268 186322 128320 186328
rect 121368 184952 121420 184958
rect 121368 184894 121420 184900
rect 118514 180840 118570 180849
rect 118514 180775 118570 180784
rect 113362 179616 113418 179625
rect 113362 179551 113418 179560
rect 102046 177576 102102 177585
rect 102046 177511 102102 177520
rect 106186 177576 106242 177585
rect 106186 177511 106242 177520
rect 108946 177576 109002 177585
rect 108946 177511 109002 177520
rect 113086 177576 113142 177585
rect 113086 177511 113142 177520
rect 113376 177041 113404 179551
rect 115848 178084 115900 178090
rect 115848 178026 115900 178032
rect 115860 177041 115888 178026
rect 118528 177449 118556 180775
rect 121380 177585 121408 184894
rect 124954 180976 125010 180985
rect 124954 180911 125010 180920
rect 125968 180940 126020 180946
rect 121920 179444 121972 179450
rect 121920 179386 121972 179392
rect 121366 177576 121422 177585
rect 121366 177511 121422 177520
rect 118514 177440 118570 177449
rect 118514 177375 118570 177384
rect 113362 177032 113418 177041
rect 113362 176967 113418 176976
rect 115846 177032 115902 177041
rect 115846 176967 115902 176976
rect 117962 177032 118018 177041
rect 117962 176967 118018 176976
rect 100758 176896 100814 176905
rect 100758 176831 100814 176840
rect 117976 176769 118004 176967
rect 121932 176769 121960 179386
rect 123300 178152 123352 178158
rect 123300 178094 123352 178100
rect 123312 176769 123340 178094
rect 124968 177585 124996 180911
rect 125968 180882 126020 180888
rect 125980 177585 126008 180882
rect 128280 177585 128308 186322
rect 129464 179512 129516 179518
rect 129464 179454 129516 179460
rect 124954 177576 125010 177585
rect 124954 177511 125010 177520
rect 125966 177576 126022 177585
rect 125966 177511 126022 177520
rect 128266 177576 128322 177585
rect 128266 177511 128322 177520
rect 128176 176860 128228 176866
rect 128176 176802 128228 176808
rect 128188 176769 128216 176802
rect 129476 176769 129504 179454
rect 131040 177313 131068 187682
rect 132408 182300 132460 182306
rect 132408 182242 132460 182248
rect 132420 177585 132448 182242
rect 133800 177585 133828 190470
rect 160848 181393 160876 244258
rect 160940 202881 160968 261530
rect 161400 224777 161428 279006
rect 162136 237153 162164 295423
rect 162228 291854 162256 326878
rect 162320 323610 162348 335679
rect 162308 323604 162360 323610
rect 162308 323546 162360 323552
rect 162584 323468 162636 323474
rect 162584 323410 162636 323416
rect 162596 319462 162624 323410
rect 162584 319456 162636 319462
rect 162584 319398 162636 319404
rect 162308 305244 162360 305250
rect 162308 305186 162360 305192
rect 162216 291848 162268 291854
rect 162216 291790 162268 291796
rect 162320 279478 162348 305186
rect 162308 279472 162360 279478
rect 162308 279414 162360 279420
rect 162216 274712 162268 274718
rect 162216 274654 162268 274660
rect 162228 251394 162256 274654
rect 162306 273864 162362 273873
rect 162306 273799 162362 273808
rect 162216 251388 162268 251394
rect 162216 251330 162268 251336
rect 162214 245712 162270 245721
rect 162214 245647 162270 245656
rect 162122 237144 162178 237153
rect 162122 237079 162178 237088
rect 161386 224768 161442 224777
rect 161386 224703 161442 224712
rect 162228 211857 162256 245647
rect 162320 240854 162348 273799
rect 162398 243536 162454 243545
rect 162398 243471 162454 243480
rect 162308 240848 162360 240854
rect 162308 240790 162360 240796
rect 162412 225622 162440 243471
rect 162400 225616 162452 225622
rect 162400 225558 162452 225564
rect 162214 211848 162270 211857
rect 162214 211783 162270 211792
rect 162872 210905 162900 409838
rect 164240 373312 164292 373318
rect 164240 373254 164292 373260
rect 163596 336864 163648 336870
rect 163596 336806 163648 336812
rect 163504 321972 163556 321978
rect 163504 321914 163556 321920
rect 163516 300257 163544 321914
rect 163608 320890 163636 336806
rect 163686 328944 163742 328953
rect 163686 328879 163742 328888
rect 163596 320884 163648 320890
rect 163596 320826 163648 320832
rect 163700 315314 163728 328879
rect 164252 324290 164280 373254
rect 164884 370592 164936 370598
rect 164884 370534 164936 370540
rect 164240 324284 164292 324290
rect 164240 324226 164292 324232
rect 163688 315308 163740 315314
rect 163688 315250 163740 315256
rect 163502 300248 163558 300257
rect 163502 300183 163558 300192
rect 163504 296744 163556 296750
rect 163504 296686 163556 296692
rect 162858 210896 162914 210905
rect 162858 210831 162914 210840
rect 160926 202872 160982 202881
rect 160926 202807 160982 202816
rect 163516 197266 163544 296686
rect 163594 280120 163650 280129
rect 163594 280055 163650 280064
rect 163608 234433 163636 280055
rect 164148 263628 164200 263634
rect 164148 263570 164200 263576
rect 164160 249898 164188 263570
rect 164148 249892 164200 249898
rect 164148 249834 164200 249840
rect 164160 249762 164188 249834
rect 164148 249756 164200 249762
rect 164148 249698 164200 249704
rect 163594 234424 163650 234433
rect 163594 234359 163650 234368
rect 163504 197260 163556 197266
rect 163504 197202 163556 197208
rect 160834 181384 160890 181393
rect 160834 181319 160890 181328
rect 148232 180872 148284 180878
rect 148232 180814 148284 180820
rect 148244 177585 148272 180814
rect 132406 177576 132462 177585
rect 132406 177511 132462 177520
rect 133786 177576 133842 177585
rect 133786 177511 133842 177520
rect 148230 177576 148286 177585
rect 148230 177511 148286 177520
rect 131026 177304 131082 177313
rect 131026 177239 131082 177248
rect 158996 176792 159048 176798
rect 100666 176760 100722 176769
rect 67548 176724 67600 176730
rect 67548 176666 67600 176672
rect 70492 176724 70544 176730
rect 100666 176695 100722 176704
rect 117962 176760 118018 176769
rect 117962 176695 118018 176704
rect 121918 176760 121974 176769
rect 121918 176695 121974 176704
rect 123298 176760 123354 176769
rect 123298 176695 123354 176704
rect 128174 176760 128230 176769
rect 128174 176695 128230 176704
rect 129462 176760 129518 176769
rect 129462 176695 129518 176704
rect 136086 176760 136142 176769
rect 136086 176695 136088 176704
rect 70492 176666 70544 176672
rect 136140 176695 136142 176704
rect 158994 176760 158996 176769
rect 159048 176760 159050 176769
rect 158994 176695 159050 176704
rect 136088 176666 136140 176672
rect 66166 129296 66222 129305
rect 66166 129231 66222 129240
rect 65522 128072 65578 128081
rect 65522 128007 65578 128016
rect 65536 127022 65564 128007
rect 65524 127016 65576 127022
rect 65524 126958 65576 126964
rect 65982 125216 66038 125225
rect 65982 125151 66038 125160
rect 65996 93158 66024 125151
rect 66074 122632 66130 122641
rect 66074 122567 66130 122576
rect 65984 93152 66036 93158
rect 65984 93094 66036 93100
rect 66088 82793 66116 122567
rect 66180 87650 66208 129231
rect 67454 123584 67510 123593
rect 67454 123519 67510 123528
rect 67362 102368 67418 102377
rect 67362 102303 67418 102312
rect 67270 100736 67326 100745
rect 67270 100671 67326 100680
rect 67284 89010 67312 100671
rect 67376 94518 67404 102303
rect 67364 94512 67416 94518
rect 67364 94454 67416 94460
rect 67272 89004 67324 89010
rect 67272 88946 67324 88952
rect 66168 87644 66220 87650
rect 66168 87586 66220 87592
rect 66074 82784 66130 82793
rect 66074 82719 66130 82728
rect 67468 78441 67496 123519
rect 67560 93226 67588 176666
rect 163516 176633 163544 197202
rect 163502 176624 163558 176633
rect 163502 176559 163558 176568
rect 164896 176254 164924 370534
rect 165066 338328 165122 338337
rect 165066 338263 165122 338272
rect 164976 331356 165028 331362
rect 164976 331298 165028 331304
rect 164988 272610 165016 331298
rect 165080 309806 165108 338263
rect 165068 309800 165120 309806
rect 165068 309742 165120 309748
rect 165158 282704 165214 282713
rect 165158 282639 165214 282648
rect 164976 272604 165028 272610
rect 164976 272546 165028 272552
rect 165068 272536 165120 272542
rect 165068 272478 165120 272484
rect 164974 269784 165030 269793
rect 164974 269719 165030 269728
rect 164988 203697 165016 269719
rect 165080 240106 165108 272478
rect 165172 253230 165200 282639
rect 165160 253224 165212 253230
rect 165160 253166 165212 253172
rect 165068 240100 165120 240106
rect 165068 240042 165120 240048
rect 166276 236745 166304 443634
rect 166356 392012 166408 392018
rect 166356 391954 166408 391960
rect 166368 300966 166396 391954
rect 168380 389224 168432 389230
rect 168380 389166 168432 389172
rect 167000 367804 167052 367810
rect 167000 367746 167052 367752
rect 166448 360324 166500 360330
rect 166448 360266 166500 360272
rect 166460 312662 166488 360266
rect 166538 335608 166594 335617
rect 166538 335543 166594 335552
rect 166552 316742 166580 335543
rect 166540 316736 166592 316742
rect 166540 316678 166592 316684
rect 166448 312656 166500 312662
rect 166448 312598 166500 312604
rect 166540 311908 166592 311914
rect 166540 311850 166592 311856
rect 166448 310548 166500 310554
rect 166448 310490 166500 310496
rect 166356 300960 166408 300966
rect 166356 300902 166408 300908
rect 166368 295322 166396 300902
rect 166356 295316 166408 295322
rect 166356 295258 166408 295264
rect 166356 285728 166408 285734
rect 166356 285670 166408 285676
rect 166262 236736 166318 236745
rect 166262 236671 166318 236680
rect 166276 227361 166304 236671
rect 166262 227352 166318 227361
rect 166262 227287 166318 227296
rect 166368 220726 166396 285670
rect 166460 275330 166488 310490
rect 166552 294642 166580 311850
rect 167012 299470 167040 367746
rect 167642 352064 167698 352073
rect 167642 351999 167698 352008
rect 167656 315353 167684 351999
rect 167642 315344 167698 315353
rect 167642 315279 167698 315288
rect 167736 309188 167788 309194
rect 167736 309130 167788 309136
rect 167000 299464 167052 299470
rect 167000 299406 167052 299412
rect 167012 298790 167040 299406
rect 167000 298784 167052 298790
rect 167000 298726 167052 298732
rect 166540 294636 166592 294642
rect 166540 294578 166592 294584
rect 167642 284336 167698 284345
rect 167642 284271 167698 284280
rect 166540 277432 166592 277438
rect 166540 277374 166592 277380
rect 166448 275324 166500 275330
rect 166448 275266 166500 275272
rect 166552 253230 166580 277374
rect 166540 253224 166592 253230
rect 166540 253166 166592 253172
rect 167656 235958 167684 284271
rect 167748 274650 167776 309130
rect 167828 291236 167880 291242
rect 167828 291178 167880 291184
rect 167840 280838 167868 291178
rect 167828 280832 167880 280838
rect 167828 280774 167880 280780
rect 167828 276072 167880 276078
rect 167828 276014 167880 276020
rect 167736 274644 167788 274650
rect 167736 274586 167788 274592
rect 167736 261520 167788 261526
rect 167736 261462 167788 261468
rect 167644 235952 167696 235958
rect 167644 235894 167696 235900
rect 167748 230382 167776 261462
rect 167840 260137 167868 276014
rect 168392 260953 168420 389166
rect 169036 286385 169064 458215
rect 179420 452668 179472 452674
rect 179420 452610 179472 452616
rect 178040 449948 178092 449954
rect 178040 449890 178092 449896
rect 173808 449200 173860 449206
rect 173808 449142 173860 449148
rect 173820 448594 173848 449142
rect 173808 448588 173860 448594
rect 173808 448530 173860 448536
rect 170404 447160 170456 447166
rect 170404 447102 170456 447108
rect 169760 438932 169812 438938
rect 169760 438874 169812 438880
rect 169116 384328 169168 384334
rect 169116 384270 169168 384276
rect 169022 286376 169078 286385
rect 169022 286311 169078 286320
rect 169036 275369 169064 286311
rect 169022 275360 169078 275369
rect 169022 275295 169078 275304
rect 168378 260944 168434 260953
rect 168378 260879 168434 260888
rect 167826 260128 167882 260137
rect 167826 260063 167882 260072
rect 168380 255332 168432 255338
rect 168380 255274 168432 255280
rect 168392 251870 168420 255274
rect 168380 251864 168432 251870
rect 168380 251806 168432 251812
rect 169128 249937 169156 384270
rect 169208 332648 169260 332654
rect 169208 332590 169260 332596
rect 169220 298858 169248 332590
rect 169208 298852 169260 298858
rect 169208 298794 169260 298800
rect 169300 285728 169352 285734
rect 169300 285670 169352 285676
rect 169206 274816 169262 274825
rect 169206 274751 169262 274760
rect 169114 249928 169170 249937
rect 169024 249892 169076 249898
rect 169114 249863 169170 249872
rect 169024 249834 169076 249840
rect 167828 249756 167880 249762
rect 167828 249698 167880 249704
rect 166908 230376 166960 230382
rect 166908 230318 166960 230324
rect 167736 230376 167788 230382
rect 167736 230318 167788 230324
rect 166920 229770 166948 230318
rect 166908 229764 166960 229770
rect 166908 229706 166960 229712
rect 166356 220720 166408 220726
rect 166356 220662 166408 220668
rect 164974 203688 165030 203697
rect 164974 203623 165030 203632
rect 166816 202156 166868 202162
rect 166816 202098 166868 202104
rect 166828 198626 166856 202098
rect 166816 198620 166868 198626
rect 166816 198562 166868 198568
rect 166262 198112 166318 198121
rect 166262 198047 166318 198056
rect 165436 179512 165488 179518
rect 165436 179454 165488 179460
rect 164976 178152 165028 178158
rect 164976 178094 165028 178100
rect 164884 176248 164936 176254
rect 164884 176190 164936 176196
rect 119436 175976 119488 175982
rect 119436 175918 119488 175924
rect 119448 175001 119476 175918
rect 135260 175228 135312 175234
rect 135260 175170 135312 175176
rect 119434 174992 119490 175001
rect 119434 174927 119490 174936
rect 135272 174865 135300 175170
rect 135258 174856 135314 174865
rect 135258 174791 135314 174800
rect 164988 169726 165016 178094
rect 165068 175976 165120 175982
rect 165068 175918 165120 175924
rect 164976 169720 165028 169726
rect 164976 169662 165028 169668
rect 165080 167006 165108 175918
rect 165448 172514 165476 179454
rect 165436 172508 165488 172514
rect 165436 172450 165488 172456
rect 165068 167000 165120 167006
rect 165068 166942 165120 166948
rect 166276 134638 166304 198047
rect 166920 192574 166948 229706
rect 167840 220697 167868 249698
rect 167826 220688 167882 220697
rect 167826 220623 167882 220632
rect 167840 219434 167868 220623
rect 167656 219406 167868 219434
rect 167000 204944 167052 204950
rect 167000 204886 167052 204892
rect 167012 202774 167040 204886
rect 167000 202768 167052 202774
rect 167000 202710 167052 202716
rect 166908 192568 166960 192574
rect 166908 192510 166960 192516
rect 167656 181490 167684 219406
rect 167736 182232 167788 182238
rect 167736 182174 167788 182180
rect 167644 181484 167696 181490
rect 167644 181426 167696 181432
rect 166448 180940 166500 180946
rect 166448 180882 166500 180888
rect 166354 179480 166410 179489
rect 166354 179415 166410 179424
rect 166368 157350 166396 179415
rect 166460 171086 166488 180882
rect 167000 176248 167052 176254
rect 167000 176190 167052 176196
rect 167012 175953 167040 176190
rect 166998 175944 167054 175953
rect 166998 175879 167054 175888
rect 166538 175536 166594 175545
rect 166538 175471 166594 175480
rect 166448 171080 166500 171086
rect 166448 171022 166500 171028
rect 166552 165578 166580 175471
rect 167642 171592 167698 171601
rect 167642 171527 167698 171536
rect 166540 165572 166592 165578
rect 166540 165514 166592 165520
rect 166356 157344 166408 157350
rect 166356 157286 166408 157292
rect 167656 152522 167684 171527
rect 167748 158710 167776 182174
rect 167826 180976 167882 180985
rect 167826 180911 167882 180920
rect 167840 169658 167868 180911
rect 169036 180130 169064 249834
rect 169128 233209 169156 249863
rect 169220 249762 169248 274751
rect 169312 274718 169340 285670
rect 169300 274712 169352 274718
rect 169300 274654 169352 274660
rect 169300 262880 169352 262886
rect 169300 262822 169352 262828
rect 169208 249756 169260 249762
rect 169208 249698 169260 249704
rect 169312 240825 169340 262822
rect 169772 261594 169800 438874
rect 170416 306374 170444 447102
rect 173256 366376 173308 366382
rect 173256 366318 173308 366324
rect 173162 343904 173218 343913
rect 173162 343839 173218 343848
rect 171874 338464 171930 338473
rect 171874 338399 171930 338408
rect 171784 334008 171836 334014
rect 171784 333950 171836 333956
rect 170586 306504 170642 306513
rect 170586 306439 170642 306448
rect 170600 306374 170628 306439
rect 170416 306346 170628 306374
rect 170402 291408 170458 291417
rect 170402 291343 170458 291352
rect 169760 261588 169812 261594
rect 169760 261530 169812 261536
rect 169772 261225 169800 261530
rect 169758 261216 169814 261225
rect 169758 261151 169814 261160
rect 170416 251938 170444 291343
rect 170496 258120 170548 258126
rect 170496 258062 170548 258068
rect 170404 251932 170456 251938
rect 170404 251874 170456 251880
rect 169760 249076 169812 249082
rect 169760 249018 169812 249024
rect 169772 242214 169800 249018
rect 170402 246256 170458 246265
rect 170402 246191 170458 246200
rect 169760 242208 169812 242214
rect 169760 242150 169812 242156
rect 169298 240816 169354 240825
rect 169298 240751 169354 240760
rect 169758 236736 169814 236745
rect 169758 236671 169760 236680
rect 169812 236671 169814 236680
rect 169760 236642 169812 236648
rect 169114 233200 169170 233209
rect 169114 233135 169170 233144
rect 169114 202328 169170 202337
rect 169114 202263 169170 202272
rect 169024 180124 169076 180130
rect 169024 180066 169076 180072
rect 169022 177032 169078 177041
rect 169022 176967 169078 176976
rect 167828 169652 167880 169658
rect 167828 169594 167880 169600
rect 169036 161430 169064 176967
rect 169024 161424 169076 161430
rect 169024 161366 169076 161372
rect 167736 158704 167788 158710
rect 167736 158646 167788 158652
rect 167644 152516 167696 152522
rect 167644 152458 167696 152464
rect 166356 147688 166408 147694
rect 166356 147630 166408 147636
rect 166264 134632 166316 134638
rect 166264 134574 166316 134580
rect 164884 129804 164936 129810
rect 164884 129746 164936 129752
rect 67638 126304 67694 126313
rect 67638 126239 67694 126248
rect 67548 93220 67600 93226
rect 67548 93162 67600 93168
rect 67652 81394 67680 126239
rect 67730 120864 67786 120873
rect 67730 120799 67786 120808
rect 67744 86290 67772 120799
rect 100666 94752 100722 94761
rect 100666 94687 100722 94696
rect 100680 93906 100708 94687
rect 124864 94512 124916 94518
rect 135812 94512 135864 94518
rect 124864 94454 124916 94460
rect 133878 94480 133934 94489
rect 100668 93900 100720 93906
rect 100668 93842 100720 93848
rect 117134 93528 117190 93537
rect 117134 93463 117190 93472
rect 121734 93528 121790 93537
rect 121734 93463 121790 93472
rect 110142 93256 110198 93265
rect 97264 93220 97316 93226
rect 110142 93191 110198 93200
rect 113822 93256 113878 93265
rect 117148 93226 117176 93463
rect 113822 93191 113878 93200
rect 117136 93220 117188 93226
rect 97264 93162 97316 93168
rect 84382 92440 84438 92449
rect 84382 92375 84438 92384
rect 89074 92440 89130 92449
rect 89074 92375 89130 92384
rect 84396 91254 84424 92375
rect 88984 91792 89036 91798
rect 88984 91734 89036 91740
rect 84384 91248 84436 91254
rect 75366 91216 75422 91225
rect 84384 91190 84436 91196
rect 86222 91216 86278 91225
rect 75366 91151 75422 91160
rect 86222 91151 86278 91160
rect 86866 91216 86922 91225
rect 86866 91151 86922 91160
rect 88246 91216 88302 91225
rect 88246 91151 88302 91160
rect 75380 88233 75408 91151
rect 75366 88224 75422 88233
rect 75366 88159 75422 88168
rect 67732 86284 67784 86290
rect 67732 86226 67784 86232
rect 86236 85513 86264 91151
rect 86222 85504 86278 85513
rect 86222 85439 86278 85448
rect 83464 84856 83516 84862
rect 83464 84798 83516 84804
rect 67640 81388 67692 81394
rect 67640 81330 67692 81336
rect 67454 78432 67510 78441
rect 67454 78367 67510 78376
rect 74446 77888 74502 77897
rect 74446 77823 74502 77832
rect 70214 76664 70270 76673
rect 70214 76599 70270 76608
rect 64418 69728 64474 69737
rect 64418 69663 64474 69672
rect 66166 61432 66222 61441
rect 66166 61367 66222 61376
rect 63408 25560 63460 25566
rect 63408 25502 63460 25508
rect 66180 3534 66208 61367
rect 68926 53136 68982 53145
rect 68926 53071 68982 53080
rect 66720 7676 66772 7682
rect 66720 7618 66772 7624
rect 63224 3528 63276 3534
rect 63224 3470 63276 3476
rect 65524 3528 65576 3534
rect 65524 3470 65576 3476
rect 66168 3528 66220 3534
rect 66168 3470 66220 3476
rect 63236 480 63264 3470
rect 64326 3360 64382 3369
rect 64326 3295 64382 3304
rect 64340 480 64368 3295
rect 65536 480 65564 3470
rect 66732 480 66760 7618
rect 68940 3534 68968 53071
rect 70228 16574 70256 76599
rect 73066 73944 73122 73953
rect 73066 73879 73122 73888
rect 71044 33856 71096 33862
rect 71044 33798 71096 33804
rect 70228 16546 70348 16574
rect 69112 4888 69164 4894
rect 69112 4830 69164 4836
rect 67916 3528 67968 3534
rect 67916 3470 67968 3476
rect 68928 3528 68980 3534
rect 68928 3470 68980 3476
rect 67928 480 67956 3470
rect 69124 480 69152 4830
rect 70320 480 70348 16546
rect 71056 3602 71084 33798
rect 71504 11824 71556 11830
rect 71504 11766 71556 11772
rect 71044 3596 71096 3602
rect 71044 3538 71096 3544
rect 71516 480 71544 11766
rect 73080 3534 73108 73879
rect 74460 3534 74488 77823
rect 75826 64288 75882 64297
rect 75826 64223 75882 64232
rect 75840 3534 75868 64223
rect 77208 60036 77260 60042
rect 77208 59978 77260 59984
rect 77220 3534 77248 59978
rect 79968 58676 80020 58682
rect 79968 58618 80020 58624
rect 77392 9036 77444 9042
rect 77392 8978 77444 8984
rect 72608 3528 72660 3534
rect 72608 3470 72660 3476
rect 73068 3528 73120 3534
rect 73068 3470 73120 3476
rect 73804 3528 73856 3534
rect 73804 3470 73856 3476
rect 74448 3528 74500 3534
rect 74448 3470 74500 3476
rect 75000 3528 75052 3534
rect 75000 3470 75052 3476
rect 75828 3528 75880 3534
rect 75828 3470 75880 3476
rect 76196 3528 76248 3534
rect 76196 3470 76248 3476
rect 77208 3528 77260 3534
rect 77208 3470 77260 3476
rect 72620 480 72648 3470
rect 73816 480 73844 3470
rect 75012 480 75040 3470
rect 76208 480 76236 3470
rect 77404 480 77432 8978
rect 79980 6914 80008 58618
rect 81346 40624 81402 40633
rect 81346 40559 81402 40568
rect 79704 6886 80008 6914
rect 78588 3460 78640 3466
rect 78588 3402 78640 3408
rect 78600 480 78628 3402
rect 79704 480 79732 6886
rect 81360 3534 81388 40559
rect 83476 31142 83504 84798
rect 86880 83502 86908 91151
rect 86868 83496 86920 83502
rect 86868 83438 86920 83444
rect 88260 82822 88288 91151
rect 88248 82816 88300 82822
rect 88248 82758 88300 82764
rect 88996 73137 89024 91734
rect 89088 91186 89116 92375
rect 96342 91896 96398 91905
rect 96342 91831 96398 91840
rect 93214 91760 93270 91769
rect 93214 91695 93270 91704
rect 91006 91216 91062 91225
rect 89076 91180 89128 91186
rect 91006 91151 91062 91160
rect 91926 91216 91982 91225
rect 91926 91151 91982 91160
rect 89076 91122 89128 91128
rect 91020 74526 91048 91151
rect 91940 88097 91968 91151
rect 93228 89729 93256 91695
rect 95146 91216 95202 91225
rect 95146 91151 95202 91160
rect 93214 89720 93270 89729
rect 93214 89655 93270 89664
rect 91926 88088 91982 88097
rect 91926 88023 91982 88032
rect 95160 81326 95188 91151
rect 96356 85377 96384 91831
rect 96342 85368 96398 85377
rect 96342 85303 96398 85312
rect 95148 81320 95200 81326
rect 95148 81262 95200 81268
rect 95146 75304 95202 75313
rect 95146 75239 95202 75248
rect 91008 74520 91060 74526
rect 91008 74462 91060 74468
rect 88982 73128 89038 73137
rect 88982 73063 89038 73072
rect 87602 62928 87658 62937
rect 87602 62863 87658 62872
rect 86866 61568 86922 61577
rect 86866 61503 86922 61512
rect 86776 44872 86828 44878
rect 86776 44814 86828 44820
rect 83464 31136 83516 31142
rect 83464 31078 83516 31084
rect 83464 26988 83516 26994
rect 83464 26930 83516 26936
rect 82728 24132 82780 24138
rect 82728 24074 82780 24080
rect 82740 3534 82768 24074
rect 80888 3528 80940 3534
rect 80888 3470 80940 3476
rect 81348 3528 81400 3534
rect 81348 3470 81400 3476
rect 82084 3528 82136 3534
rect 82084 3470 82136 3476
rect 82728 3528 82780 3534
rect 82728 3470 82780 3476
rect 83280 3528 83332 3534
rect 83280 3470 83332 3476
rect 80900 480 80928 3470
rect 82096 480 82124 3470
rect 83292 480 83320 3470
rect 83476 3398 83504 26930
rect 84108 22772 84160 22778
rect 84108 22714 84160 22720
rect 84120 3534 84148 22714
rect 86788 16574 86816 44814
rect 86696 16546 86816 16574
rect 85488 14544 85540 14550
rect 85488 14486 85540 14492
rect 85500 3534 85528 14486
rect 85672 3596 85724 3602
rect 85672 3538 85724 3544
rect 84108 3528 84160 3534
rect 84108 3470 84160 3476
rect 84476 3528 84528 3534
rect 84476 3470 84528 3476
rect 85488 3528 85540 3534
rect 85488 3470 85540 3476
rect 83464 3392 83516 3398
rect 83464 3334 83516 3340
rect 84488 480 84516 3470
rect 85684 480 85712 3538
rect 86696 3482 86724 16546
rect 86880 6914 86908 61503
rect 86788 6886 86908 6914
rect 86788 3602 86816 6886
rect 86776 3596 86828 3602
rect 86776 3538 86828 3544
rect 86696 3454 86908 3482
rect 87616 3466 87644 62863
rect 89626 58576 89682 58585
rect 89626 58511 89682 58520
rect 88248 43444 88300 43450
rect 88248 43386 88300 43392
rect 88260 6914 88288 43386
rect 87984 6886 88288 6914
rect 86880 480 86908 3454
rect 87604 3460 87656 3466
rect 87604 3402 87656 3408
rect 87984 480 88012 6886
rect 89640 3330 89668 58511
rect 93768 57248 93820 57254
rect 93768 57190 93820 57196
rect 91008 55888 91060 55894
rect 91008 55830 91060 55836
rect 91020 3534 91048 55830
rect 90364 3528 90416 3534
rect 90364 3470 90416 3476
rect 91008 3528 91060 3534
rect 91008 3470 91060 3476
rect 91560 3528 91612 3534
rect 91560 3470 91612 3476
rect 89168 3324 89220 3330
rect 89168 3266 89220 3272
rect 89628 3324 89680 3330
rect 89628 3266 89680 3272
rect 89180 480 89208 3266
rect 90376 480 90404 3470
rect 91572 480 91600 3470
rect 93780 3466 93808 57190
rect 95056 26920 95108 26926
rect 95056 26862 95108 26868
rect 95068 3466 95096 26862
rect 92756 3460 92808 3466
rect 92756 3402 92808 3408
rect 93768 3460 93820 3466
rect 93768 3402 93820 3408
rect 93952 3460 94004 3466
rect 93952 3402 94004 3408
rect 95056 3460 95108 3466
rect 95056 3402 95108 3408
rect 92768 480 92796 3402
rect 93964 480 93992 3402
rect 95160 480 95188 75239
rect 97276 46306 97304 93162
rect 106924 93152 106976 93158
rect 106924 93094 106976 93100
rect 106832 92608 106884 92614
rect 106832 92550 106884 92556
rect 99104 92540 99156 92546
rect 99104 92482 99156 92488
rect 99116 92449 99144 92482
rect 106844 92449 106872 92550
rect 99102 92440 99158 92449
rect 99102 92375 99158 92384
rect 106830 92440 106886 92449
rect 106830 92375 106886 92384
rect 99286 91760 99342 91769
rect 99286 91695 99342 91704
rect 97906 91352 97962 91361
rect 97906 91287 97962 91296
rect 97814 91216 97870 91225
rect 97814 91151 97870 91160
rect 97828 84182 97856 91151
rect 97816 84176 97868 84182
rect 97816 84118 97868 84124
rect 97920 80034 97948 91287
rect 99194 91216 99250 91225
rect 99194 91151 99250 91160
rect 97908 80028 97960 80034
rect 97908 79970 97960 79976
rect 99208 71738 99236 91151
rect 99300 89593 99328 91695
rect 102046 91352 102102 91361
rect 102046 91287 102102 91296
rect 100022 91216 100078 91225
rect 100022 91151 100078 91160
rect 101218 91216 101274 91225
rect 101218 91151 101274 91160
rect 101954 91216 102010 91225
rect 101954 91151 102010 91160
rect 99286 89584 99342 89593
rect 99286 89519 99342 89528
rect 100036 86737 100064 91151
rect 101232 86873 101260 91151
rect 101218 86864 101274 86873
rect 101218 86799 101274 86808
rect 100022 86728 100078 86737
rect 100022 86663 100078 86672
rect 99286 82104 99342 82113
rect 99286 82039 99342 82048
rect 99196 71732 99248 71738
rect 99196 71674 99248 71680
rect 97908 54528 97960 54534
rect 97908 54470 97960 54476
rect 97264 46300 97316 46306
rect 97264 46242 97316 46248
rect 96528 18692 96580 18698
rect 96528 18634 96580 18640
rect 96540 6914 96568 18634
rect 96264 6886 96568 6914
rect 96264 480 96292 6886
rect 97920 3466 97948 54470
rect 99300 3466 99328 82039
rect 101968 78577 101996 91151
rect 101954 78568 102010 78577
rect 101954 78503 102010 78512
rect 102060 70378 102088 91287
rect 103426 91216 103482 91225
rect 104438 91216 104494 91225
rect 103426 91151 103482 91160
rect 104256 91180 104308 91186
rect 102048 70372 102100 70378
rect 102048 70314 102100 70320
rect 103440 69018 103468 91151
rect 104438 91151 104494 91160
rect 105542 91216 105598 91225
rect 105542 91151 105598 91160
rect 106094 91216 106150 91225
rect 106094 91151 106150 91160
rect 104256 91122 104308 91128
rect 104162 71224 104218 71233
rect 104162 71159 104218 71168
rect 103428 69012 103480 69018
rect 103428 68954 103480 68960
rect 101404 68332 101456 68338
rect 101404 68274 101456 68280
rect 101416 53106 101444 68274
rect 101404 53100 101456 53106
rect 101404 53042 101456 53048
rect 102048 53100 102100 53106
rect 102048 53042 102100 53048
rect 100668 20052 100720 20058
rect 100668 19994 100720 20000
rect 100680 3466 100708 19994
rect 102060 3466 102088 53042
rect 103428 50380 103480 50386
rect 103428 50322 103480 50328
rect 103440 6914 103468 50322
rect 104176 8974 104204 71159
rect 104268 64870 104296 91122
rect 104452 85542 104480 91151
rect 105556 88330 105584 91151
rect 105544 88324 105596 88330
rect 105544 88266 105596 88272
rect 104440 85536 104492 85542
rect 104440 85478 104492 85484
rect 106108 66162 106136 91151
rect 106936 80073 106964 93094
rect 109682 92440 109738 92449
rect 109682 92375 109738 92384
rect 107566 91216 107622 91225
rect 107566 91151 107622 91160
rect 108486 91216 108542 91225
rect 108486 91151 108542 91160
rect 107016 87644 107068 87650
rect 107016 87586 107068 87592
rect 106922 80064 106978 80073
rect 106922 79999 106978 80008
rect 106188 76560 106240 76566
rect 106188 76502 106240 76508
rect 106096 66156 106148 66162
rect 106096 66098 106148 66104
rect 104256 64864 104308 64870
rect 104256 64806 104308 64812
rect 104532 10328 104584 10334
rect 104532 10270 104584 10276
rect 104164 8968 104216 8974
rect 104164 8910 104216 8916
rect 103348 6886 103468 6914
rect 97448 3460 97500 3466
rect 97448 3402 97500 3408
rect 97908 3460 97960 3466
rect 97908 3402 97960 3408
rect 98644 3460 98696 3466
rect 98644 3402 98696 3408
rect 99288 3460 99340 3466
rect 99288 3402 99340 3408
rect 99840 3460 99892 3466
rect 99840 3402 99892 3408
rect 100668 3460 100720 3466
rect 100668 3402 100720 3408
rect 101036 3460 101088 3466
rect 101036 3402 101088 3408
rect 102048 3460 102100 3466
rect 102048 3402 102100 3408
rect 97460 480 97488 3402
rect 98656 480 98684 3402
rect 99852 480 99880 3402
rect 101048 480 101076 3402
rect 102232 2100 102284 2106
rect 102232 2042 102284 2048
rect 102244 480 102272 2042
rect 103348 480 103376 6886
rect 104544 480 104572 10270
rect 106200 3466 106228 76502
rect 107028 75886 107056 87586
rect 107016 75880 107068 75886
rect 107016 75822 107068 75828
rect 107580 67590 107608 91151
rect 108304 89004 108356 89010
rect 108304 88946 108356 88952
rect 107568 67584 107620 67590
rect 107568 67526 107620 67532
rect 108316 66230 108344 88946
rect 108500 87961 108528 91151
rect 109696 91118 109724 92375
rect 109684 91112 109736 91118
rect 109684 91054 109736 91060
rect 108486 87952 108542 87961
rect 108486 87887 108542 87896
rect 108304 66224 108356 66230
rect 108304 66166 108356 66172
rect 110156 56574 110184 93191
rect 112444 92540 112496 92546
rect 112444 92482 112496 92488
rect 110696 92472 110748 92478
rect 110694 92440 110696 92449
rect 110748 92440 110750 92449
rect 110694 92375 110750 92384
rect 111522 92440 111578 92449
rect 111522 92375 111578 92384
rect 111064 91248 111116 91254
rect 110234 91216 110290 91225
rect 111064 91190 111116 91196
rect 110234 91151 110290 91160
rect 110248 84153 110276 91151
rect 110234 84144 110290 84153
rect 110234 84079 110290 84088
rect 111076 82754 111104 91190
rect 111536 91050 111564 92375
rect 111524 91044 111576 91050
rect 111524 90986 111576 90992
rect 111064 82748 111116 82754
rect 111064 82690 111116 82696
rect 111708 75200 111760 75206
rect 111708 75142 111760 75148
rect 110144 56568 110196 56574
rect 110144 56510 110196 56516
rect 108948 51740 109000 51746
rect 108948 51682 109000 51688
rect 106922 42120 106978 42129
rect 106922 42055 106978 42064
rect 106936 6914 106964 42055
rect 107016 8968 107068 8974
rect 107016 8910 107068 8916
rect 106844 6886 106964 6914
rect 105728 3460 105780 3466
rect 105728 3402 105780 3408
rect 106188 3460 106240 3466
rect 106188 3402 106240 3408
rect 105740 480 105768 3402
rect 106844 2174 106872 6886
rect 107028 3482 107056 8910
rect 106936 3454 107056 3482
rect 108960 3466 108988 51682
rect 111616 35284 111668 35290
rect 111616 35226 111668 35232
rect 110328 32496 110380 32502
rect 110328 32438 110380 32444
rect 110340 3466 110368 32438
rect 108120 3460 108172 3466
rect 106832 2168 106884 2174
rect 106832 2110 106884 2116
rect 106936 480 106964 3454
rect 108120 3402 108172 3408
rect 108948 3460 109000 3466
rect 108948 3402 109000 3408
rect 109316 3460 109368 3466
rect 109316 3402 109368 3408
rect 110328 3460 110380 3466
rect 110328 3402 110380 3408
rect 110512 3460 110564 3466
rect 110512 3402 110564 3408
rect 108132 480 108160 3402
rect 109328 480 109356 3402
rect 110524 480 110552 3402
rect 111628 480 111656 35226
rect 111720 3466 111748 75142
rect 112456 57934 112484 92482
rect 112718 91216 112774 91225
rect 112718 91151 112774 91160
rect 112732 86970 112760 91151
rect 113836 89457 113864 93191
rect 117136 93162 117188 93168
rect 121748 93158 121776 93463
rect 121736 93152 121788 93158
rect 121736 93094 121788 93100
rect 116584 92608 116636 92614
rect 116584 92550 116636 92556
rect 114282 91352 114338 91361
rect 114282 91287 114338 91296
rect 115754 91352 115810 91361
rect 115754 91287 115810 91296
rect 113822 89448 113878 89457
rect 113822 89383 113878 89392
rect 112720 86964 112772 86970
rect 112720 86906 112772 86912
rect 112444 57928 112496 57934
rect 112444 57870 112496 57876
rect 114296 52426 114324 91287
rect 114374 91216 114430 91225
rect 114374 91151 114430 91160
rect 114388 60722 114416 91151
rect 115204 91112 115256 91118
rect 115204 91054 115256 91060
rect 114376 60716 114428 60722
rect 114376 60658 114428 60664
rect 115216 55214 115244 91054
rect 115768 85474 115796 91287
rect 115846 91216 115902 91225
rect 115846 91151 115902 91160
rect 115756 85468 115808 85474
rect 115756 85410 115808 85416
rect 115860 62014 115888 91151
rect 116596 67522 116624 92550
rect 124126 92440 124182 92449
rect 124126 92375 124182 92384
rect 119802 91760 119858 91769
rect 119802 91695 119858 91704
rect 118606 91352 118662 91361
rect 118606 91287 118662 91296
rect 118514 91216 118570 91225
rect 118514 91151 118570 91160
rect 117228 73840 117280 73846
rect 117228 73782 117280 73788
rect 116584 67516 116636 67522
rect 116584 67458 116636 67464
rect 115848 62008 115900 62014
rect 115848 61950 115900 61956
rect 115204 55208 115256 55214
rect 115204 55150 115256 55156
rect 114284 52420 114336 52426
rect 114284 52362 114336 52368
rect 115848 49088 115900 49094
rect 115848 49030 115900 49036
rect 112444 39432 112496 39438
rect 112444 39374 112496 39380
rect 112456 13190 112484 39374
rect 112444 13184 112496 13190
rect 112444 13126 112496 13132
rect 112812 10396 112864 10402
rect 112812 10338 112864 10344
rect 111708 3460 111760 3466
rect 111708 3402 111760 3408
rect 112824 480 112852 10338
rect 115860 3466 115888 49030
rect 117240 3466 117268 73782
rect 118528 53786 118556 91151
rect 118516 53780 118568 53786
rect 118516 53722 118568 53728
rect 118620 48278 118648 91287
rect 119816 89690 119844 91695
rect 124034 91488 124090 91497
rect 124034 91423 124090 91432
rect 119894 91216 119950 91225
rect 119894 91151 119950 91160
rect 120446 91216 120502 91225
rect 120446 91151 120502 91160
rect 120722 91216 120778 91225
rect 120722 91151 120778 91160
rect 122746 91216 122802 91225
rect 122746 91151 122802 91160
rect 119804 89684 119856 89690
rect 119804 89626 119856 89632
rect 119908 51066 119936 91151
rect 120460 85241 120488 91151
rect 120736 88262 120764 91151
rect 120724 88256 120776 88262
rect 120724 88198 120776 88204
rect 120446 85232 120502 85241
rect 120446 85167 120502 85176
rect 122760 78674 122788 91151
rect 122748 78668 122800 78674
rect 122748 78610 122800 78616
rect 119988 71052 120040 71058
rect 119988 70994 120040 71000
rect 119896 51060 119948 51066
rect 119896 51002 119948 51008
rect 118608 48272 118660 48278
rect 118608 48214 118660 48220
rect 118608 13184 118660 13190
rect 118608 13126 118660 13132
rect 118620 3466 118648 13126
rect 119896 6248 119948 6254
rect 119896 6190 119948 6196
rect 115204 3460 115256 3466
rect 115204 3402 115256 3408
rect 115848 3460 115900 3466
rect 115848 3402 115900 3408
rect 116400 3460 116452 3466
rect 116400 3402 116452 3408
rect 117228 3460 117280 3466
rect 117228 3402 117280 3408
rect 117596 3460 117648 3466
rect 117596 3402 117648 3408
rect 118608 3460 118660 3466
rect 118608 3402 118660 3408
rect 118792 3460 118844 3466
rect 118792 3402 118844 3408
rect 114008 3392 114060 3398
rect 114008 3334 114060 3340
rect 114020 480 114048 3334
rect 115216 480 115244 3402
rect 116412 480 116440 3402
rect 117608 480 117636 3402
rect 118804 480 118832 3402
rect 119908 480 119936 6190
rect 120000 3466 120028 70994
rect 122102 65648 122158 65657
rect 122102 65583 122158 65592
rect 119988 3460 120040 3466
rect 119988 3402 120040 3408
rect 122116 3369 122144 65583
rect 124048 64802 124076 91423
rect 124140 90982 124168 92375
rect 124128 90976 124180 90982
rect 124128 90918 124180 90924
rect 124126 83464 124182 83473
rect 124126 83399 124182 83408
rect 124036 64796 124088 64802
rect 124036 64738 124088 64744
rect 122748 28280 122800 28286
rect 122748 28222 122800 28228
rect 122102 3360 122158 3369
rect 122760 3330 122788 28222
rect 124140 3534 124168 83399
rect 124876 63442 124904 94454
rect 135812 94454 135864 94460
rect 133878 94415 133934 94424
rect 133892 92478 133920 94415
rect 135824 93673 135852 94454
rect 135810 93664 135866 93673
rect 135810 93599 135866 93608
rect 135994 93664 136050 93673
rect 135994 93599 136050 93608
rect 136008 93401 136036 93599
rect 135994 93392 136050 93401
rect 135994 93327 136050 93336
rect 133880 92472 133932 92478
rect 136088 92472 136140 92478
rect 133880 92414 133932 92420
rect 136086 92440 136088 92449
rect 136140 92440 136142 92449
rect 136086 92375 136142 92384
rect 151450 92440 151506 92449
rect 151450 92375 151506 92384
rect 125414 91352 125470 91361
rect 125414 91287 125470 91296
rect 126886 91352 126942 91361
rect 126886 91287 126942 91296
rect 125428 70310 125456 91287
rect 125506 91216 125562 91225
rect 125506 91151 125562 91160
rect 126794 91216 126850 91225
rect 126794 91151 126850 91160
rect 125416 70304 125468 70310
rect 125416 70246 125468 70252
rect 125520 63510 125548 91151
rect 126808 84114 126836 91151
rect 126796 84108 126848 84114
rect 126796 84050 126848 84056
rect 126244 83496 126296 83502
rect 126244 83438 126296 83444
rect 126256 73098 126284 83438
rect 126900 79966 126928 91287
rect 128266 91216 128322 91225
rect 128266 91151 128322 91160
rect 129646 91216 129702 91225
rect 129646 91151 129702 91160
rect 132406 91216 132462 91225
rect 132406 91151 132462 91160
rect 126888 79960 126940 79966
rect 126888 79902 126940 79908
rect 128280 77246 128308 91151
rect 128268 77240 128320 77246
rect 128268 77182 128320 77188
rect 126244 73092 126296 73098
rect 126244 73034 126296 73040
rect 125508 63504 125560 63510
rect 125508 63446 125560 63452
rect 124864 63436 124916 63442
rect 124864 63378 124916 63384
rect 129660 59362 129688 91151
rect 130382 68504 130438 68513
rect 130382 68439 130438 68448
rect 129648 59356 129700 59362
rect 129648 59298 129700 59304
rect 125508 44940 125560 44946
rect 125508 44882 125560 44888
rect 125520 3534 125548 44882
rect 126244 21480 126296 21486
rect 126244 21422 126296 21428
rect 126256 3602 126284 21422
rect 126244 3596 126296 3602
rect 126244 3538 126296 3544
rect 130396 3534 130424 68439
rect 132420 62082 132448 91151
rect 151464 91118 151492 92375
rect 159364 91860 159416 91866
rect 159364 91802 159416 91808
rect 151542 91352 151598 91361
rect 151542 91287 151598 91296
rect 151452 91112 151504 91118
rect 151452 91054 151504 91060
rect 150440 86284 150492 86290
rect 150440 86226 150492 86232
rect 150452 81433 150480 86226
rect 150438 81424 150494 81433
rect 150438 81359 150494 81368
rect 142802 80880 142858 80889
rect 142802 80815 142858 80824
rect 132408 62076 132460 62082
rect 132408 62018 132460 62024
rect 136454 11656 136510 11665
rect 136454 11591 136510 11600
rect 132958 8936 133014 8945
rect 132958 8871 133014 8880
rect 123484 3528 123536 3534
rect 123484 3470 123536 3476
rect 124128 3528 124180 3534
rect 124128 3470 124180 3476
rect 124680 3528 124732 3534
rect 124680 3470 124732 3476
rect 125508 3528 125560 3534
rect 125508 3470 125560 3476
rect 129372 3528 129424 3534
rect 129372 3470 129424 3476
rect 130384 3528 130436 3534
rect 130384 3470 130436 3476
rect 122102 3295 122158 3304
rect 122288 3324 122340 3330
rect 122288 3266 122340 3272
rect 122748 3324 122800 3330
rect 122748 3266 122800 3272
rect 121092 2168 121144 2174
rect 121092 2110 121144 2116
rect 121104 480 121132 2110
rect 122300 480 122328 3266
rect 123496 480 123524 3470
rect 124692 480 124720 3470
rect 125874 3360 125930 3369
rect 125874 3295 125930 3304
rect 125888 480 125916 3295
rect 129384 480 129412 3470
rect 132972 480 133000 8871
rect 136468 480 136496 11591
rect 142816 8974 142844 80815
rect 151556 73166 151584 91287
rect 151634 91216 151690 91225
rect 151634 91151 151690 91160
rect 152462 91216 152518 91225
rect 152462 91151 152518 91160
rect 151648 78606 151676 91151
rect 152476 86902 152504 91151
rect 157340 91112 157392 91118
rect 157340 91054 157392 91060
rect 157352 89622 157380 91054
rect 157340 89616 157392 89622
rect 157340 89558 157392 89564
rect 152464 86896 152516 86902
rect 152464 86838 152516 86844
rect 159376 79966 159404 91802
rect 159364 79960 159416 79966
rect 159364 79902 159416 79908
rect 151636 78600 151688 78606
rect 151636 78542 151688 78548
rect 151544 73160 151596 73166
rect 151544 73102 151596 73108
rect 164896 69018 164924 129746
rect 166264 122868 166316 122874
rect 166264 122810 166316 122816
rect 165068 107704 165120 107710
rect 165068 107646 165120 107652
rect 164976 95940 165028 95946
rect 164976 95882 165028 95888
rect 164988 73098 165016 95882
rect 165080 90817 165108 107646
rect 165066 90808 165122 90817
rect 165066 90743 165122 90752
rect 166276 88262 166304 122810
rect 166368 92478 166396 147630
rect 169024 144968 169076 144974
rect 169024 144910 169076 144916
rect 167828 129056 167880 129062
rect 167828 128998 167880 129004
rect 167736 113824 167788 113830
rect 167736 113766 167788 113772
rect 166446 112024 166502 112033
rect 166446 111959 166502 111968
rect 166460 93906 166488 111959
rect 167644 110492 167696 110498
rect 167644 110434 167696 110440
rect 166540 105596 166592 105602
rect 166540 105538 166592 105544
rect 166448 93900 166500 93906
rect 166448 93842 166500 93848
rect 166356 92472 166408 92478
rect 166356 92414 166408 92420
rect 166552 89690 166580 105538
rect 166540 89684 166592 89690
rect 166540 89626 166592 89632
rect 166264 88256 166316 88262
rect 166264 88198 166316 88204
rect 167656 86737 167684 110434
rect 167748 94518 167776 113766
rect 167840 111761 167868 128998
rect 168288 115252 168340 115258
rect 168288 115194 168340 115200
rect 167826 111752 167882 111761
rect 167826 111687 167882 111696
rect 168300 110129 168328 115194
rect 168286 110120 168342 110129
rect 168286 110055 168342 110064
rect 168012 108996 168064 109002
rect 168012 108938 168064 108944
rect 168024 108769 168052 108938
rect 168010 108760 168066 108769
rect 168010 108695 168066 108704
rect 167918 105496 167974 105505
rect 167918 105431 167974 105440
rect 167828 98048 167880 98054
rect 167828 97990 167880 97996
rect 167736 94512 167788 94518
rect 167736 94454 167788 94460
rect 167642 86728 167698 86737
rect 167642 86663 167698 86672
rect 167840 85513 167868 97990
rect 167932 93537 167960 105431
rect 167918 93528 167974 93537
rect 167918 93463 167974 93472
rect 169036 92177 169064 144910
rect 169128 141438 169156 202263
rect 169758 189816 169814 189825
rect 169758 189751 169814 189760
rect 169772 189106 169800 189751
rect 169760 189100 169812 189106
rect 169760 189042 169812 189048
rect 169206 179616 169262 179625
rect 169206 179551 169262 179560
rect 169220 164218 169248 179551
rect 169208 164212 169260 164218
rect 169208 164154 169260 164160
rect 169206 151056 169262 151065
rect 169206 150991 169262 151000
rect 169116 141432 169168 141438
rect 169116 141374 169168 141380
rect 169116 122120 169168 122126
rect 169116 122062 169168 122068
rect 169022 92168 169078 92177
rect 169022 92103 169078 92112
rect 169128 90982 169156 122062
rect 169220 109002 169248 150991
rect 170416 135930 170444 246191
rect 170508 182889 170536 258062
rect 170600 237318 170628 306346
rect 171796 247790 171824 333950
rect 171888 281450 171916 338399
rect 172060 324284 172112 324290
rect 172060 324226 172112 324232
rect 172072 315382 172100 324226
rect 171968 315376 172020 315382
rect 171968 315318 172020 315324
rect 172060 315376 172112 315382
rect 172060 315318 172112 315324
rect 171876 281444 171928 281450
rect 171876 281386 171928 281392
rect 171980 269074 172008 315318
rect 171968 269068 172020 269074
rect 171968 269010 172020 269016
rect 171968 260160 172020 260166
rect 171968 260102 172020 260108
rect 171876 258732 171928 258738
rect 171876 258674 171928 258680
rect 171784 247784 171836 247790
rect 171784 247726 171836 247732
rect 170588 237312 170640 237318
rect 170588 237254 170640 237260
rect 171784 211812 171836 211818
rect 171784 211754 171836 211760
rect 170588 189168 170640 189174
rect 170588 189110 170640 189116
rect 170494 182880 170550 182889
rect 170494 182815 170550 182824
rect 170494 180840 170550 180849
rect 170494 180775 170550 180784
rect 170508 166938 170536 180775
rect 170496 166932 170548 166938
rect 170496 166874 170548 166880
rect 170600 164150 170628 189110
rect 170588 164144 170640 164150
rect 170588 164086 170640 164092
rect 171796 142866 171824 211754
rect 171888 191729 171916 258674
rect 171980 219366 172008 260102
rect 171968 219360 172020 219366
rect 171968 219302 172020 219308
rect 172796 217320 172848 217326
rect 172796 217262 172848 217268
rect 172808 212401 172836 217262
rect 172426 212392 172482 212401
rect 172426 212327 172482 212336
rect 172794 212392 172850 212401
rect 172794 212327 172850 212336
rect 172440 211206 172468 212327
rect 172428 211200 172480 211206
rect 172428 211142 172480 211148
rect 171968 192500 172020 192506
rect 171968 192442 172020 192448
rect 171874 191720 171930 191729
rect 171874 191655 171930 191664
rect 171980 178770 172008 192442
rect 172060 182300 172112 182306
rect 172060 182242 172112 182248
rect 171968 178764 172020 178770
rect 171968 178706 172020 178712
rect 171876 178084 171928 178090
rect 171876 178026 171928 178032
rect 171888 165510 171916 178026
rect 172072 173874 172100 182242
rect 172060 173868 172112 173874
rect 172060 173810 172112 173816
rect 171876 165504 171928 165510
rect 171876 165446 171928 165452
rect 173176 144226 173204 343839
rect 173268 298217 173296 366318
rect 173254 298208 173310 298217
rect 173254 298143 173310 298152
rect 173268 285734 173296 298143
rect 173440 291848 173492 291854
rect 173440 291790 173492 291796
rect 173256 285728 173308 285734
rect 173256 285670 173308 285676
rect 173452 235278 173480 291790
rect 173820 242214 173848 448530
rect 177396 396092 177448 396098
rect 177396 396034 177448 396040
rect 174728 358896 174780 358902
rect 174728 358838 174780 358844
rect 174634 347984 174690 347993
rect 174634 347919 174690 347928
rect 174542 330168 174598 330177
rect 174542 330103 174598 330112
rect 173808 242208 173860 242214
rect 173808 242150 173860 242156
rect 173820 239873 173848 242150
rect 173806 239864 173862 239873
rect 173806 239799 173862 239808
rect 173440 235272 173492 235278
rect 173440 235214 173492 235220
rect 173254 232792 173310 232801
rect 173254 232727 173310 232736
rect 173268 197334 173296 232727
rect 173256 197328 173308 197334
rect 173256 197270 173308 197276
rect 173254 178392 173310 178401
rect 173254 178327 173310 178336
rect 173268 162858 173296 178327
rect 173256 162852 173308 162858
rect 173256 162794 173308 162800
rect 173164 144220 173216 144226
rect 173164 144162 173216 144168
rect 171784 142860 171836 142866
rect 171784 142802 171836 142808
rect 171784 136672 171836 136678
rect 171784 136614 171836 136620
rect 170404 135924 170456 135930
rect 170404 135866 170456 135872
rect 170404 117360 170456 117366
rect 170404 117302 170456 117308
rect 169208 108996 169260 109002
rect 169208 108938 169260 108944
rect 169208 102808 169260 102814
rect 169208 102750 169260 102756
rect 169116 90976 169168 90982
rect 169116 90918 169168 90924
rect 169024 90364 169076 90370
rect 169024 90306 169076 90312
rect 167826 85504 167882 85513
rect 167826 85439 167882 85448
rect 164976 73092 165028 73098
rect 164976 73034 165028 73040
rect 164884 69012 164936 69018
rect 164884 68954 164936 68960
rect 160742 68368 160798 68377
rect 160742 68303 160798 68312
rect 146944 47592 146996 47598
rect 146944 47534 146996 47540
rect 142804 8968 142856 8974
rect 142804 8910 142856 8916
rect 146956 6186 146984 47534
rect 160756 10305 160784 68303
rect 169036 63442 169064 90306
rect 169220 78606 169248 102750
rect 169300 100768 169352 100774
rect 169300 100710 169352 100716
rect 169312 82754 169340 100710
rect 170416 91050 170444 117302
rect 170586 106856 170642 106865
rect 170586 106791 170642 106800
rect 170496 103556 170548 103562
rect 170496 103498 170548 103504
rect 170404 91044 170456 91050
rect 170404 90986 170456 90992
rect 169300 82748 169352 82754
rect 169300 82690 169352 82696
rect 170508 80073 170536 103498
rect 170600 85241 170628 106791
rect 170680 99408 170732 99414
rect 170680 99350 170732 99356
rect 170586 85232 170642 85241
rect 170586 85167 170642 85176
rect 170692 82822 170720 99350
rect 170680 82816 170732 82822
rect 170680 82758 170732 82764
rect 170494 80064 170550 80073
rect 170494 79999 170550 80008
rect 169208 78600 169260 78606
rect 169208 78542 169260 78548
rect 169024 63436 169076 63442
rect 169024 63378 169076 63384
rect 171796 62014 171824 136614
rect 173164 132524 173216 132530
rect 173164 132466 173216 132472
rect 171876 124908 171928 124914
rect 171876 124850 171928 124856
rect 171888 86902 171916 124850
rect 171968 109064 172020 109070
rect 171968 109006 172020 109012
rect 171876 86896 171928 86902
rect 171876 86838 171928 86844
rect 171874 84960 171930 84969
rect 171874 84895 171930 84904
rect 171888 73137 171916 84895
rect 171980 84182 172008 109006
rect 173176 87961 173204 132466
rect 173256 126268 173308 126274
rect 173256 126210 173308 126216
rect 173268 94489 173296 126210
rect 173348 109132 173400 109138
rect 173348 109074 173400 109080
rect 173254 94480 173310 94489
rect 173254 94415 173310 94424
rect 173162 87952 173218 87961
rect 173162 87887 173218 87896
rect 173256 87644 173308 87650
rect 173256 87586 173308 87592
rect 171968 84176 172020 84182
rect 171968 84118 172020 84124
rect 171874 73128 171930 73137
rect 171874 73063 171930 73072
rect 173268 67522 173296 87586
rect 173360 85377 173388 109074
rect 173440 101448 173492 101454
rect 173440 101390 173492 101396
rect 173346 85368 173402 85377
rect 173346 85303 173402 85312
rect 173452 77246 173480 101390
rect 173440 77240 173492 77246
rect 173440 77182 173492 77188
rect 173256 67516 173308 67522
rect 173256 67458 173308 67464
rect 171784 62008 171836 62014
rect 171784 61950 171836 61956
rect 174556 43518 174584 330103
rect 174648 253881 174676 347919
rect 174740 311166 174768 358838
rect 176108 356176 176160 356182
rect 176108 356118 176160 356124
rect 176014 342408 176070 342417
rect 176014 342343 176070 342352
rect 174728 311160 174780 311166
rect 174728 311102 174780 311108
rect 175924 270564 175976 270570
rect 175924 270506 175976 270512
rect 174728 264240 174780 264246
rect 174728 264182 174780 264188
rect 174634 253872 174690 253881
rect 174634 253807 174690 253816
rect 174636 243024 174688 243030
rect 174636 242966 174688 242972
rect 174648 196654 174676 242966
rect 174740 222154 174768 264182
rect 174728 222148 174780 222154
rect 174728 222090 174780 222096
rect 174636 196648 174688 196654
rect 174636 196590 174688 196596
rect 174636 186380 174688 186386
rect 174636 186322 174688 186328
rect 174648 171018 174676 186322
rect 174728 176792 174780 176798
rect 174728 176734 174780 176740
rect 174636 171012 174688 171018
rect 174636 170954 174688 170960
rect 174740 167686 174768 176734
rect 174728 167680 174780 167686
rect 174728 167622 174780 167628
rect 174636 127628 174688 127634
rect 174636 127570 174688 127576
rect 174648 78674 174676 127570
rect 174818 126304 174874 126313
rect 174818 126239 174874 126248
rect 174832 89593 174860 126239
rect 174818 89584 174874 89593
rect 174818 89519 174874 89528
rect 174728 88868 174780 88874
rect 174728 88810 174780 88816
rect 174636 78668 174688 78674
rect 174636 78610 174688 78616
rect 174740 52426 174768 88810
rect 175936 77994 175964 270506
rect 176028 236065 176056 342343
rect 176120 271862 176148 356118
rect 177304 326392 177356 326398
rect 177304 326334 177356 326340
rect 177316 283626 177344 326334
rect 177304 283620 177356 283626
rect 177304 283562 177356 283568
rect 177304 281444 177356 281450
rect 177304 281386 177356 281392
rect 176108 271856 176160 271862
rect 176108 271798 176160 271804
rect 176106 265160 176162 265169
rect 176106 265095 176162 265104
rect 176014 236056 176070 236065
rect 176014 235991 176070 236000
rect 176120 235929 176148 265095
rect 176106 235920 176162 235929
rect 176106 235855 176162 235864
rect 176120 219434 176148 235855
rect 176028 219406 176148 219434
rect 176028 198257 176056 219406
rect 176014 198248 176070 198257
rect 176014 198183 176070 198192
rect 176016 193860 176068 193866
rect 176016 193802 176068 193808
rect 176028 116521 176056 193802
rect 177316 138718 177344 281386
rect 177408 267889 177436 396034
rect 177488 339584 177540 339590
rect 177488 339526 177540 339532
rect 177500 276554 177528 339526
rect 177488 276548 177540 276554
rect 177488 276490 177540 276496
rect 177488 272604 177540 272610
rect 177488 272546 177540 272552
rect 177394 267880 177450 267889
rect 177394 267815 177450 267824
rect 177408 233073 177436 267815
rect 177500 253298 177528 272546
rect 177948 256828 178000 256834
rect 177948 256770 178000 256776
rect 177488 253292 177540 253298
rect 177488 253234 177540 253240
rect 177856 248464 177908 248470
rect 177856 248406 177908 248412
rect 177868 244934 177896 248406
rect 177856 244928 177908 244934
rect 177856 244870 177908 244876
rect 177394 233064 177450 233073
rect 177394 232999 177450 233008
rect 177960 180033 177988 256770
rect 178052 255270 178080 449890
rect 178776 350600 178828 350606
rect 178776 350542 178828 350548
rect 178682 341184 178738 341193
rect 178682 341119 178738 341128
rect 178696 330449 178724 341119
rect 178682 330440 178738 330449
rect 178682 330375 178738 330384
rect 178682 320784 178738 320793
rect 178682 320719 178738 320728
rect 178040 255264 178092 255270
rect 178040 255206 178092 255212
rect 178052 254590 178080 255206
rect 178040 254584 178092 254590
rect 178040 254526 178092 254532
rect 177946 180024 178002 180033
rect 177946 179959 178002 179968
rect 177394 178256 177450 178265
rect 177394 178191 177450 178200
rect 177408 162790 177436 178191
rect 177396 162784 177448 162790
rect 177396 162726 177448 162732
rect 177304 138712 177356 138718
rect 177304 138654 177356 138660
rect 177580 120148 177632 120154
rect 177580 120090 177632 120096
rect 176108 118720 176160 118726
rect 176108 118662 176160 118668
rect 176014 116512 176070 116521
rect 176014 116447 176070 116456
rect 176016 104916 176068 104922
rect 176016 104858 176068 104864
rect 175924 77988 175976 77994
rect 175924 77930 175976 77936
rect 176028 74526 176056 104858
rect 176120 89457 176148 118662
rect 177304 116000 177356 116006
rect 177304 115942 177356 115948
rect 176106 89448 176162 89457
rect 176106 89383 176162 89392
rect 176016 74520 176068 74526
rect 176016 74462 176068 74468
rect 177316 55214 177344 115942
rect 177488 110560 177540 110566
rect 177488 110502 177540 110508
rect 177396 97300 177448 97306
rect 177396 97242 177448 97248
rect 177304 55208 177356 55214
rect 177304 55150 177356 55156
rect 174728 52420 174780 52426
rect 174728 52362 174780 52368
rect 177408 48278 177436 97242
rect 177500 71738 177528 110502
rect 177592 93226 177620 120090
rect 177580 93220 177632 93226
rect 177580 93162 177632 93168
rect 177488 71732 177540 71738
rect 177488 71674 177540 71680
rect 177396 48272 177448 48278
rect 177396 48214 177448 48220
rect 174544 43512 174596 43518
rect 174544 43454 174596 43460
rect 160742 10296 160798 10305
rect 160742 10231 160798 10240
rect 146944 6180 146996 6186
rect 146944 6122 146996 6128
rect 178696 4865 178724 320719
rect 178788 314022 178816 350542
rect 178958 332888 179014 332897
rect 178958 332823 179014 332832
rect 178776 314016 178828 314022
rect 178776 313958 178828 313964
rect 178776 262268 178828 262274
rect 178776 262210 178828 262216
rect 178788 6186 178816 262210
rect 178868 249348 178920 249354
rect 178868 249290 178920 249296
rect 178880 224874 178908 249290
rect 178972 249121 179000 332823
rect 179432 253994 179460 452610
rect 201500 445800 201552 445806
rect 201500 445742 201552 445748
rect 193864 374060 193916 374066
rect 193864 374002 193916 374008
rect 180800 371272 180852 371278
rect 180800 371214 180852 371220
rect 180064 349172 180116 349178
rect 180064 349114 180116 349120
rect 179512 282940 179564 282946
rect 179512 282882 179564 282888
rect 179524 282198 179552 282882
rect 179512 282192 179564 282198
rect 179512 282134 179564 282140
rect 179340 253978 179460 253994
rect 179328 253972 179460 253978
rect 179380 253966 179460 253972
rect 179328 253914 179380 253920
rect 178958 249112 179014 249121
rect 178958 249047 179014 249056
rect 179340 235929 179368 253914
rect 179880 252612 179932 252618
rect 179880 252554 179932 252560
rect 179892 249354 179920 252554
rect 179880 249348 179932 249354
rect 179880 249290 179932 249296
rect 179326 235920 179382 235929
rect 179326 235855 179382 235864
rect 180076 233170 180104 349114
rect 180156 327140 180208 327146
rect 180156 327082 180208 327088
rect 180168 284306 180196 327082
rect 180156 284300 180208 284306
rect 180156 284242 180208 284248
rect 180708 282192 180760 282198
rect 180708 282134 180760 282140
rect 180340 253224 180392 253230
rect 180340 253166 180392 253172
rect 180154 236056 180210 236065
rect 180154 235991 180210 236000
rect 180064 233164 180116 233170
rect 180064 233106 180116 233112
rect 178868 224868 178920 224874
rect 178868 224810 178920 224816
rect 178880 182850 178908 224810
rect 180062 211848 180118 211857
rect 180062 211783 180118 211792
rect 178868 182844 178920 182850
rect 178868 182786 178920 182792
rect 178958 182200 179014 182209
rect 178958 182135 179014 182144
rect 178972 155922 179000 182135
rect 178960 155916 179012 155922
rect 178960 155858 179012 155864
rect 178868 134564 178920 134570
rect 178868 134506 178920 134512
rect 178880 88874 178908 134506
rect 178960 89004 179012 89010
rect 178960 88946 179012 88952
rect 178868 88868 178920 88874
rect 178868 88810 178920 88816
rect 178972 75886 179000 88946
rect 178960 75880 179012 75886
rect 178960 75822 179012 75828
rect 180076 47666 180104 211783
rect 180168 140078 180196 235991
rect 180246 231296 180302 231305
rect 180246 231231 180302 231240
rect 180260 198694 180288 231231
rect 180352 229090 180380 253166
rect 180340 229084 180392 229090
rect 180340 229026 180392 229032
rect 180248 198688 180300 198694
rect 180248 198630 180300 198636
rect 180720 186998 180748 282134
rect 180812 270473 180840 371214
rect 185582 367296 185638 367305
rect 185582 367231 185638 367240
rect 184296 354748 184348 354754
rect 184296 354690 184348 354696
rect 182822 346624 182878 346633
rect 182822 346559 182878 346568
rect 181444 278044 181496 278050
rect 181444 277986 181496 277992
rect 180798 270464 180854 270473
rect 180798 270399 180854 270408
rect 181258 270464 181314 270473
rect 181258 270399 181314 270408
rect 181272 269793 181300 270399
rect 181258 269784 181314 269793
rect 181258 269719 181314 269728
rect 181456 256834 181484 277986
rect 181536 276548 181588 276554
rect 181536 276490 181588 276496
rect 181444 256828 181496 256834
rect 181444 256770 181496 256776
rect 181442 253872 181498 253881
rect 181442 253807 181498 253816
rect 180708 186992 180760 186998
rect 180708 186934 180760 186940
rect 180248 183660 180300 183666
rect 180248 183602 180300 183608
rect 180260 157282 180288 183602
rect 180248 157276 180300 157282
rect 180248 157218 180300 157224
rect 180340 142180 180392 142186
rect 180340 142122 180392 142128
rect 180248 140820 180300 140826
rect 180248 140762 180300 140768
rect 180156 140072 180208 140078
rect 180156 140014 180208 140020
rect 180156 91792 180208 91798
rect 180156 91734 180208 91740
rect 180064 47660 180116 47666
rect 180064 47602 180116 47608
rect 178776 6180 178828 6186
rect 178776 6122 178828 6128
rect 180168 4894 180196 91734
rect 180260 70310 180288 140762
rect 180352 94081 180380 142122
rect 181456 136649 181484 253807
rect 181548 229770 181576 276490
rect 181628 269204 181680 269210
rect 181628 269146 181680 269152
rect 181640 234530 181668 269146
rect 182732 247716 182784 247722
rect 182732 247658 182784 247664
rect 182744 240009 182772 247658
rect 182730 240000 182786 240009
rect 182730 239935 182786 239944
rect 181628 234524 181680 234530
rect 181628 234466 181680 234472
rect 181536 229764 181588 229770
rect 181536 229706 181588 229712
rect 181640 191185 181668 234466
rect 181626 191176 181682 191185
rect 181626 191111 181682 191120
rect 181534 176896 181590 176905
rect 181534 176831 181590 176840
rect 181548 158642 181576 176831
rect 181536 158636 181588 158642
rect 181536 158578 181588 158584
rect 181536 137284 181588 137290
rect 181536 137226 181588 137232
rect 181442 136640 181498 136649
rect 181442 136575 181498 136584
rect 181444 131776 181496 131782
rect 181444 131718 181496 131724
rect 180338 94072 180394 94081
rect 180338 94007 180394 94016
rect 181456 91866 181484 131718
rect 181548 105505 181576 137226
rect 181628 106344 181680 106350
rect 181628 106286 181680 106292
rect 181534 105496 181590 105505
rect 181534 105431 181590 105440
rect 181536 103624 181588 103630
rect 181536 103566 181588 103572
rect 181444 91860 181496 91866
rect 181444 91802 181496 91808
rect 181442 84824 181498 84833
rect 181442 84759 181498 84768
rect 180248 70304 180300 70310
rect 180248 70246 180300 70252
rect 181456 14550 181484 84759
rect 181548 81394 181576 103566
rect 181640 88097 181668 106286
rect 181626 88088 181682 88097
rect 181626 88023 181682 88032
rect 181536 81388 181588 81394
rect 181536 81330 181588 81336
rect 182836 33833 182864 346559
rect 183006 291272 183062 291281
rect 183006 291207 183062 291216
rect 182916 290488 182968 290494
rect 182916 290430 182968 290436
rect 182928 282878 182956 290430
rect 182916 282872 182968 282878
rect 182916 282814 182968 282820
rect 182916 271856 182968 271862
rect 182916 271798 182968 271804
rect 182928 196761 182956 271798
rect 183020 230489 183048 291207
rect 184202 266384 184258 266393
rect 184202 266319 184258 266328
rect 183006 230480 183062 230489
rect 183006 230415 183062 230424
rect 182914 196752 182970 196761
rect 182914 196687 182970 196696
rect 182916 185020 182968 185026
rect 182916 184962 182968 184968
rect 182928 160070 182956 184962
rect 182916 160064 182968 160070
rect 182916 160006 182968 160012
rect 183008 150476 183060 150482
rect 183008 150418 183060 150424
rect 183020 115258 183048 150418
rect 183008 115252 183060 115258
rect 183008 115194 183060 115200
rect 182914 115152 182970 115161
rect 182914 115087 182970 115096
rect 182928 66162 182956 115087
rect 183100 114572 183152 114578
rect 183100 114514 183152 114520
rect 183112 88330 183140 114514
rect 183100 88324 183152 88330
rect 183100 88266 183152 88272
rect 182916 66156 182968 66162
rect 182916 66098 182968 66104
rect 182822 33824 182878 33833
rect 182822 33759 182878 33768
rect 181444 14544 181496 14550
rect 181444 14486 181496 14492
rect 184216 10305 184244 266319
rect 184308 259418 184336 354690
rect 184388 351960 184440 351966
rect 184388 351902 184440 351908
rect 184400 266529 184428 351902
rect 184478 285968 184534 285977
rect 184478 285903 184534 285912
rect 184386 266520 184442 266529
rect 184386 266455 184442 266464
rect 184296 259412 184348 259418
rect 184296 259354 184348 259360
rect 184492 219434 184520 285903
rect 184570 279576 184626 279585
rect 184570 279511 184626 279520
rect 184584 220833 184612 279511
rect 184848 256760 184900 256766
rect 184848 256702 184900 256708
rect 184570 220824 184626 220833
rect 184570 220759 184626 220768
rect 184308 219406 184520 219434
rect 184308 217841 184336 219406
rect 184294 217832 184350 217841
rect 184294 217767 184350 217776
rect 184308 178702 184336 217767
rect 184860 184210 184888 256702
rect 184848 184204 184900 184210
rect 184848 184146 184900 184152
rect 185596 178945 185624 367231
rect 186964 361616 187016 361622
rect 186964 361558 187016 361564
rect 185676 327752 185728 327758
rect 185676 327694 185728 327700
rect 185688 297401 185716 327694
rect 186976 318170 187004 361558
rect 192576 357536 192628 357542
rect 192576 357478 192628 357484
rect 191102 345264 191158 345273
rect 191102 345199 191158 345208
rect 187054 339824 187110 339833
rect 187054 339759 187110 339768
rect 187068 327758 187096 339759
rect 189722 334384 189778 334393
rect 189722 334319 189778 334328
rect 187056 327752 187108 327758
rect 187056 327694 187108 327700
rect 186964 318164 187016 318170
rect 186964 318106 187016 318112
rect 188436 316804 188488 316810
rect 188436 316746 188488 316752
rect 188344 300892 188396 300898
rect 188344 300834 188396 300840
rect 186964 298852 187016 298858
rect 186964 298794 187016 298800
rect 185674 297392 185730 297401
rect 185674 297327 185730 297336
rect 185674 294128 185730 294137
rect 185674 294063 185730 294072
rect 185688 262886 185716 294063
rect 185768 283620 185820 283626
rect 185768 283562 185820 283568
rect 185780 276758 185808 283562
rect 186976 277438 187004 298794
rect 187148 288516 187200 288522
rect 187148 288458 187200 288464
rect 186964 277432 187016 277438
rect 186964 277374 187016 277380
rect 185768 276752 185820 276758
rect 185768 276694 185820 276700
rect 186964 275392 187016 275398
rect 186964 275334 187016 275340
rect 186228 270564 186280 270570
rect 186228 270506 186280 270512
rect 185676 262880 185728 262886
rect 185676 262822 185728 262828
rect 185768 262268 185820 262274
rect 185768 262210 185820 262216
rect 185676 249892 185728 249898
rect 185676 249834 185728 249840
rect 185688 226302 185716 249834
rect 185780 245750 185808 262210
rect 185768 245744 185820 245750
rect 185768 245686 185820 245692
rect 185676 226296 185728 226302
rect 185676 226238 185728 226244
rect 185582 178936 185638 178945
rect 185582 178871 185638 178880
rect 184296 178696 184348 178702
rect 184296 178638 184348 178644
rect 185688 177313 185716 226238
rect 185780 202337 185808 245686
rect 186240 231577 186268 270506
rect 186320 253292 186372 253298
rect 186320 253234 186372 253240
rect 186332 252686 186360 253234
rect 186320 252680 186372 252686
rect 186320 252622 186372 252628
rect 185950 231568 186006 231577
rect 185950 231503 186006 231512
rect 186226 231568 186282 231577
rect 186226 231503 186282 231512
rect 185964 231169 185992 231503
rect 185950 231160 186006 231169
rect 185950 231095 186006 231104
rect 186976 219434 187004 275334
rect 187160 273970 187188 288458
rect 187148 273964 187200 273970
rect 187148 273906 187200 273912
rect 187056 273284 187108 273290
rect 187056 273226 187108 273232
rect 187068 245682 187096 273226
rect 187608 252680 187660 252686
rect 187608 252622 187660 252628
rect 187514 249112 187570 249121
rect 187514 249047 187570 249056
rect 187528 248577 187556 249047
rect 187514 248568 187570 248577
rect 187514 248503 187570 248512
rect 187056 245676 187108 245682
rect 187056 245618 187108 245624
rect 186964 219428 187016 219434
rect 186964 219370 187016 219376
rect 186976 218074 187004 219370
rect 186964 218068 187016 218074
rect 186964 218010 187016 218016
rect 186964 213240 187016 213246
rect 186964 213182 187016 213188
rect 186976 204105 187004 213182
rect 186962 204096 187018 204105
rect 186962 204031 187018 204040
rect 185766 202328 185822 202337
rect 185766 202263 185822 202272
rect 187068 194041 187096 245618
rect 187148 218068 187200 218074
rect 187148 218010 187200 218016
rect 187054 194032 187110 194041
rect 187054 193967 187110 193976
rect 186962 189680 187018 189689
rect 186962 189615 187018 189624
rect 185766 178120 185822 178129
rect 185766 178055 185822 178064
rect 185674 177304 185730 177313
rect 185674 177239 185730 177248
rect 185780 155854 185808 178055
rect 185768 155848 185820 155854
rect 185768 155790 185820 155796
rect 185676 153264 185728 153270
rect 185676 153206 185728 153212
rect 184388 146328 184440 146334
rect 184388 146270 184440 146276
rect 184296 144220 184348 144226
rect 184296 144162 184348 144168
rect 184308 28354 184336 144162
rect 184400 113830 184428 146270
rect 185584 134632 185636 134638
rect 185584 134574 185636 134580
rect 184388 113824 184440 113830
rect 184388 113766 184440 113772
rect 184480 113212 184532 113218
rect 184480 113154 184532 113160
rect 184492 85542 184520 113154
rect 184480 85536 184532 85542
rect 184480 85478 184532 85484
rect 184296 28348 184348 28354
rect 184296 28290 184348 28296
rect 185596 21321 185624 134574
rect 185688 89622 185716 153206
rect 185768 93220 185820 93226
rect 185768 93162 185820 93168
rect 185676 89616 185728 89622
rect 185676 89558 185728 89564
rect 185780 84114 185808 93162
rect 185768 84108 185820 84114
rect 185768 84050 185820 84056
rect 185582 21312 185638 21321
rect 185582 21247 185638 21256
rect 184202 10296 184258 10305
rect 184202 10231 184258 10240
rect 186976 8974 187004 189615
rect 187160 175273 187188 218010
rect 187528 217326 187556 248503
rect 187516 217320 187568 217326
rect 187516 217262 187568 217268
rect 187620 198121 187648 252622
rect 187698 228304 187754 228313
rect 187698 228239 187754 228248
rect 187712 220833 187740 228239
rect 187698 220824 187754 220833
rect 187698 220759 187754 220768
rect 187606 198112 187662 198121
rect 187606 198047 187662 198056
rect 187146 175264 187202 175273
rect 187146 175199 187202 175208
rect 187056 135312 187108 135318
rect 187056 135254 187108 135260
rect 187068 93945 187096 135254
rect 187148 122936 187200 122942
rect 187148 122878 187200 122884
rect 187054 93936 187110 93945
rect 187054 93871 187110 93880
rect 187160 93158 187188 122878
rect 187148 93152 187200 93158
rect 187148 93094 187200 93100
rect 188356 13025 188384 300834
rect 188448 256698 188476 316746
rect 188620 275324 188672 275330
rect 188620 275266 188672 275272
rect 188528 259480 188580 259486
rect 188528 259422 188580 259428
rect 188436 256692 188488 256698
rect 188436 256634 188488 256640
rect 188436 242956 188488 242962
rect 188436 242898 188488 242904
rect 188448 234598 188476 242898
rect 188436 234592 188488 234598
rect 188436 234534 188488 234540
rect 188540 211070 188568 259422
rect 188632 226302 188660 275266
rect 189736 244905 189764 334319
rect 189908 318096 189960 318102
rect 189908 318038 189960 318044
rect 189814 283520 189870 283529
rect 189814 283455 189870 283464
rect 189722 244896 189778 244905
rect 189722 244831 189778 244840
rect 188620 226296 188672 226302
rect 188620 226238 188672 226244
rect 189828 223417 189856 283455
rect 189920 264246 189948 318038
rect 191116 266286 191144 345199
rect 191196 338224 191248 338230
rect 191196 338166 191248 338172
rect 191208 317393 191236 338166
rect 191194 317384 191250 317393
rect 191194 317319 191250 317328
rect 192484 315376 192536 315382
rect 192484 315318 192536 315324
rect 191196 302932 191248 302938
rect 191196 302874 191248 302880
rect 191208 281450 191236 302874
rect 191654 288824 191710 288833
rect 191654 288759 191710 288768
rect 191196 281444 191248 281450
rect 191196 281386 191248 281392
rect 191196 271176 191248 271182
rect 191196 271118 191248 271124
rect 191104 266280 191156 266286
rect 191104 266222 191156 266228
rect 189908 264240 189960 264246
rect 189908 264182 189960 264188
rect 189908 261588 189960 261594
rect 189908 261530 189960 261536
rect 189920 231810 189948 261530
rect 191104 251252 191156 251258
rect 191104 251194 191156 251200
rect 190368 245472 190420 245478
rect 190368 245414 190420 245420
rect 190000 244928 190052 244934
rect 190000 244870 190052 244876
rect 190012 231810 190040 244870
rect 189908 231804 189960 231810
rect 189908 231746 189960 231752
rect 190000 231804 190052 231810
rect 190000 231746 190052 231752
rect 189814 223408 189870 223417
rect 189814 223343 189870 223352
rect 189920 219434 189948 231746
rect 189736 219406 189948 219434
rect 189736 216073 189764 219406
rect 189722 216064 189778 216073
rect 189722 215999 189778 216008
rect 188528 211064 188580 211070
rect 188528 211006 188580 211012
rect 188434 204912 188490 204921
rect 188434 204847 188490 204856
rect 188448 86358 188476 204847
rect 188540 185706 188568 211006
rect 189724 200796 189776 200802
rect 189724 200738 189776 200744
rect 188620 187740 188672 187746
rect 188620 187682 188672 187688
rect 188528 185700 188580 185706
rect 188528 185642 188580 185648
rect 188632 173806 188660 187682
rect 188620 173800 188672 173806
rect 188620 173742 188672 173748
rect 189736 145625 189764 200738
rect 190380 189825 190408 245414
rect 191116 244497 191144 251194
rect 191208 249762 191236 271118
rect 191196 249756 191248 249762
rect 191196 249698 191248 249704
rect 191196 247104 191248 247110
rect 191196 247046 191248 247052
rect 191102 244488 191158 244497
rect 191102 244423 191158 244432
rect 190828 228404 190880 228410
rect 190828 228346 190880 228352
rect 190840 226137 190868 228346
rect 190826 226128 190882 226137
rect 190826 226063 190882 226072
rect 190366 189816 190422 189825
rect 190366 189751 190422 189760
rect 189722 145616 189778 145625
rect 189722 145551 189778 145560
rect 189816 143608 189868 143614
rect 189816 143550 189868 143556
rect 188526 136640 188582 136649
rect 188526 136575 188582 136584
rect 188436 86352 188488 86358
rect 188436 86294 188488 86300
rect 188540 24206 188568 136575
rect 189722 113792 189778 113801
rect 189722 113727 189778 113736
rect 189736 60722 189764 113727
rect 189828 101454 189856 143550
rect 191116 133113 191144 244423
rect 191208 216646 191236 247046
rect 191668 228449 191696 288759
rect 191748 279472 191800 279478
rect 191748 279414 191800 279420
rect 191654 228440 191710 228449
rect 191654 228375 191710 228384
rect 191196 216640 191248 216646
rect 191196 216582 191248 216588
rect 191208 203726 191236 216582
rect 191656 215960 191708 215966
rect 191656 215902 191708 215908
rect 191668 213858 191696 215902
rect 191656 213852 191708 213858
rect 191656 213794 191708 213800
rect 191196 203720 191248 203726
rect 191196 203662 191248 203668
rect 191288 203584 191340 203590
rect 191288 203526 191340 203532
rect 191300 198694 191328 203526
rect 191288 198688 191340 198694
rect 191288 198630 191340 198636
rect 191196 189780 191248 189786
rect 191196 189722 191248 189728
rect 191102 133104 191158 133113
rect 191102 133039 191158 133048
rect 191104 124228 191156 124234
rect 191104 124170 191156 124176
rect 189906 118824 189962 118833
rect 189906 118759 189962 118768
rect 189816 101448 189868 101454
rect 189816 101390 189868 101396
rect 189920 86970 189948 118759
rect 189908 86964 189960 86970
rect 189908 86906 189960 86912
rect 191116 64802 191144 124170
rect 191208 89049 191236 189722
rect 191760 188358 191788 279414
rect 191840 277840 191892 277846
rect 191840 277782 191892 277788
rect 191852 277438 191880 277782
rect 191840 277432 191892 277438
rect 191840 277374 191892 277380
rect 191852 245478 191880 277374
rect 191840 245472 191892 245478
rect 191840 245414 191892 245420
rect 192496 233209 192524 315318
rect 192588 302297 192616 357478
rect 192574 302288 192630 302297
rect 192574 302223 192630 302232
rect 193126 302288 193182 302297
rect 193126 302223 193182 302232
rect 192576 284980 192628 284986
rect 192576 284922 192628 284928
rect 192588 268394 192616 284922
rect 193140 277953 193168 302223
rect 193126 277944 193182 277953
rect 193126 277879 193182 277888
rect 193876 272377 193904 374002
rect 196624 362976 196676 362982
rect 196624 362918 196676 362924
rect 195334 360224 195390 360233
rect 195334 360159 195390 360168
rect 195244 345092 195296 345098
rect 195244 345034 195296 345040
rect 195152 320204 195204 320210
rect 195152 320146 195204 320152
rect 195164 319433 195192 320146
rect 195150 319424 195206 319433
rect 195150 319359 195206 319368
rect 193956 299600 194008 299606
rect 193956 299542 194008 299548
rect 193968 290494 193996 299542
rect 193956 290488 194008 290494
rect 193956 290430 194008 290436
rect 194048 285728 194100 285734
rect 194048 285670 194100 285676
rect 193862 272368 193918 272377
rect 193862 272303 193918 272312
rect 192576 268388 192628 268394
rect 192576 268330 192628 268336
rect 192588 256426 192616 268330
rect 193956 267028 194008 267034
rect 193956 266970 194008 266976
rect 192758 260944 192814 260953
rect 192758 260879 192814 260888
rect 192576 256420 192628 256426
rect 192576 256362 192628 256368
rect 192668 253972 192720 253978
rect 192668 253914 192720 253920
rect 192576 244316 192628 244322
rect 192576 244258 192628 244264
rect 192482 233200 192538 233209
rect 192482 233135 192538 233144
rect 191840 221468 191892 221474
rect 191840 221410 191892 221416
rect 191852 216646 191880 221410
rect 191930 220960 191986 220969
rect 191930 220895 191986 220904
rect 191840 216640 191892 216646
rect 191840 216582 191892 216588
rect 191944 213926 191972 220895
rect 191932 213920 191984 213926
rect 191932 213862 191984 213868
rect 192484 211200 192536 211206
rect 192484 211142 192536 211148
rect 191748 188352 191800 188358
rect 191748 188294 191800 188300
rect 192496 179926 192524 211142
rect 192588 191146 192616 244258
rect 192680 225865 192708 253914
rect 192772 244322 192800 260879
rect 193864 256420 193916 256426
rect 193864 256362 193916 256368
rect 192760 244316 192812 244322
rect 192760 244258 192812 244264
rect 192760 241528 192812 241534
rect 192760 241470 192812 241476
rect 192772 228857 192800 241470
rect 192758 228848 192814 228857
rect 192758 228783 192814 228792
rect 192666 225856 192722 225865
rect 192666 225791 192722 225800
rect 192576 191140 192628 191146
rect 192576 191082 192628 191088
rect 192668 190528 192720 190534
rect 192668 190470 192720 190476
rect 192484 179920 192536 179926
rect 192484 179862 192536 179868
rect 192576 179444 192628 179450
rect 192576 179386 192628 179392
rect 192588 168366 192616 179386
rect 192680 175166 192708 190470
rect 193876 177342 193904 256362
rect 193968 240825 193996 266970
rect 194060 264217 194088 285670
rect 194508 276684 194560 276690
rect 194508 276626 194560 276632
rect 194046 264208 194102 264217
rect 194046 264143 194102 264152
rect 194416 247784 194468 247790
rect 194416 247726 194468 247732
rect 194428 245206 194456 247726
rect 194520 246090 194548 276626
rect 194874 270464 194930 270473
rect 194874 270399 194930 270408
rect 194888 269890 194916 270399
rect 194876 269884 194928 269890
rect 194876 269826 194928 269832
rect 195256 247042 195284 345034
rect 195348 307834 195376 360159
rect 195428 329860 195480 329866
rect 195428 329802 195480 329808
rect 195440 318102 195468 329802
rect 195428 318096 195480 318102
rect 195428 318038 195480 318044
rect 195336 307828 195388 307834
rect 195336 307770 195388 307776
rect 195336 298240 195388 298246
rect 195336 298182 195388 298188
rect 195348 267714 195376 298182
rect 195426 291544 195482 291553
rect 195426 291479 195482 291488
rect 195440 280129 195468 291479
rect 195426 280120 195482 280129
rect 195426 280055 195482 280064
rect 195520 270632 195572 270638
rect 195520 270574 195572 270580
rect 195428 269136 195480 269142
rect 195428 269078 195480 269084
rect 195336 267708 195388 267714
rect 195336 267650 195388 267656
rect 195440 257446 195468 269078
rect 195532 261526 195560 270574
rect 195888 266416 195940 266422
rect 195888 266358 195940 266364
rect 195520 261520 195572 261526
rect 195520 261462 195572 261468
rect 195428 257440 195480 257446
rect 195428 257382 195480 257388
rect 195796 251864 195848 251870
rect 195796 251806 195848 251812
rect 195704 249756 195756 249762
rect 195704 249698 195756 249704
rect 195244 247036 195296 247042
rect 195244 246978 195296 246984
rect 194508 246084 194560 246090
rect 194508 246026 194560 246032
rect 195336 246084 195388 246090
rect 195336 246026 195388 246032
rect 194416 245200 194468 245206
rect 194416 245142 194468 245148
rect 194428 245018 194456 245142
rect 194428 244990 194548 245018
rect 194414 244896 194470 244905
rect 194414 244831 194470 244840
rect 193954 240816 194010 240825
rect 193954 240751 194010 240760
rect 193954 215928 194010 215937
rect 193954 215863 194010 215872
rect 193968 204921 193996 215863
rect 194428 214577 194456 244831
rect 194414 214568 194470 214577
rect 194414 214503 194470 214512
rect 193954 204912 194010 204921
rect 193954 204847 194010 204856
rect 194520 189786 194548 244990
rect 195244 222896 195296 222902
rect 195244 222838 195296 222844
rect 195256 212430 195284 222838
rect 195244 212424 195296 212430
rect 195244 212366 195296 212372
rect 195242 205048 195298 205057
rect 195348 205018 195376 246026
rect 195716 240514 195744 249698
rect 195704 240508 195756 240514
rect 195704 240450 195756 240456
rect 195612 229764 195664 229770
rect 195612 229706 195664 229712
rect 195624 224874 195652 229706
rect 195808 228410 195836 251806
rect 195900 229129 195928 266358
rect 195980 255264 196032 255270
rect 195978 255232 195980 255241
rect 196032 255232 196034 255241
rect 195978 255167 196034 255176
rect 196348 249824 196400 249830
rect 196348 249766 196400 249772
rect 196360 245070 196388 249766
rect 196348 245064 196400 245070
rect 196348 245006 196400 245012
rect 196636 235657 196664 362918
rect 198002 349480 198058 349489
rect 198002 349415 198058 349424
rect 196714 347848 196770 347857
rect 196714 347783 196770 347792
rect 196728 330614 196756 347783
rect 196716 330608 196768 330614
rect 196716 330550 196768 330556
rect 196716 329180 196768 329186
rect 196716 329122 196768 329128
rect 196728 264489 196756 329122
rect 198016 309262 198044 349415
rect 200762 342272 200818 342281
rect 200762 342207 200818 342216
rect 198094 329896 198150 329905
rect 198094 329831 198150 329840
rect 198108 313954 198136 329831
rect 199474 322144 199530 322153
rect 199474 322079 199530 322088
rect 199384 319524 199436 319530
rect 199384 319466 199436 319472
rect 198096 313948 198148 313954
rect 198096 313890 198148 313896
rect 198096 309800 198148 309806
rect 198096 309742 198148 309748
rect 198004 309256 198056 309262
rect 198004 309198 198056 309204
rect 198108 305046 198136 309742
rect 198648 309256 198700 309262
rect 198648 309198 198700 309204
rect 198096 305040 198148 305046
rect 198096 304982 198148 304988
rect 198556 305040 198608 305046
rect 198556 304982 198608 304988
rect 196808 295384 196860 295390
rect 196808 295326 196860 295332
rect 196820 281518 196848 295326
rect 198094 292904 198150 292913
rect 198094 292839 198150 292848
rect 197358 291408 197414 291417
rect 197358 291343 197414 291352
rect 197372 290494 197400 291343
rect 197360 290488 197412 290494
rect 197360 290430 197412 290436
rect 198002 287464 198058 287473
rect 198002 287399 198058 287408
rect 197360 284300 197412 284306
rect 197360 284242 197412 284248
rect 197372 283801 197400 284242
rect 197358 283792 197414 283801
rect 197358 283727 197414 283736
rect 197358 282432 197414 282441
rect 197358 282367 197414 282376
rect 197372 282198 197400 282367
rect 197360 282192 197412 282198
rect 197360 282134 197412 282140
rect 196808 281512 196860 281518
rect 196808 281454 196860 281460
rect 197360 281444 197412 281450
rect 197360 281386 197412 281392
rect 197372 280809 197400 281386
rect 197358 280800 197414 280809
rect 197358 280735 197414 280744
rect 197358 280256 197414 280265
rect 197358 280191 197414 280200
rect 197372 278050 197400 280191
rect 197452 279472 197504 279478
rect 197450 279440 197452 279449
rect 197504 279440 197506 279449
rect 197450 279375 197506 279384
rect 197450 278624 197506 278633
rect 197450 278559 197506 278568
rect 197360 278044 197412 278050
rect 197360 277986 197412 277992
rect 197358 277944 197414 277953
rect 197358 277879 197414 277888
rect 197372 277273 197400 277879
rect 197464 277846 197492 278559
rect 197452 277840 197504 277846
rect 197452 277782 197504 277788
rect 197358 277264 197414 277273
rect 197358 277199 197414 277208
rect 197544 276752 197596 276758
rect 197358 276720 197414 276729
rect 197544 276694 197596 276700
rect 197358 276655 197360 276664
rect 197412 276655 197414 276664
rect 197360 276626 197412 276632
rect 197450 275904 197506 275913
rect 197450 275839 197506 275848
rect 197358 273728 197414 273737
rect 197358 273663 197414 273672
rect 197372 273290 197400 273663
rect 197360 273284 197412 273290
rect 197360 273226 197412 273232
rect 197358 272912 197414 272921
rect 197358 272847 197414 272856
rect 197372 271930 197400 272847
rect 197464 272542 197492 275839
rect 197556 274553 197584 276694
rect 197542 274544 197598 274553
rect 197542 274479 197598 274488
rect 197452 272536 197504 272542
rect 197452 272478 197504 272484
rect 197360 271924 197412 271930
rect 197360 271866 197412 271872
rect 197818 271552 197874 271561
rect 197818 271487 197874 271496
rect 197358 271008 197414 271017
rect 197358 270943 197414 270952
rect 197372 270570 197400 270943
rect 197832 270638 197860 271487
rect 197820 270632 197872 270638
rect 197820 270574 197872 270580
rect 197360 270564 197412 270570
rect 197360 270506 197412 270512
rect 197358 270192 197414 270201
rect 197358 270127 197414 270136
rect 197372 269210 197400 270127
rect 197452 269884 197504 269890
rect 197452 269826 197504 269832
rect 197464 269385 197492 269826
rect 197450 269376 197506 269385
rect 197450 269311 197506 269320
rect 197360 269204 197412 269210
rect 197360 269146 197412 269152
rect 197360 269068 197412 269074
rect 197360 269010 197412 269016
rect 197372 268841 197400 269010
rect 197358 268832 197414 268841
rect 197358 268767 197414 268776
rect 198016 267734 198044 287399
rect 197924 267706 198044 267734
rect 197360 266280 197412 266286
rect 197360 266222 197412 266228
rect 197372 265849 197400 266222
rect 197358 265840 197414 265849
rect 197358 265775 197414 265784
rect 196714 264480 196770 264489
rect 196714 264415 196770 264424
rect 197358 263664 197414 263673
rect 197358 263599 197360 263608
rect 197412 263599 197414 263608
rect 197360 263570 197412 263576
rect 197358 263120 197414 263129
rect 197358 263055 197414 263064
rect 197372 262274 197400 263055
rect 197360 262268 197412 262274
rect 197360 262210 197412 262216
rect 197450 260128 197506 260137
rect 197450 260063 197506 260072
rect 197464 259486 197492 260063
rect 197452 259480 197504 259486
rect 197452 259422 197504 259428
rect 197360 259412 197412 259418
rect 197360 259354 197412 259360
rect 197372 258777 197400 259354
rect 197358 258768 197414 258777
rect 197924 258738 197952 267706
rect 198002 267200 198058 267209
rect 198002 267135 198058 267144
rect 198016 266422 198044 267135
rect 198004 266416 198056 266422
rect 198004 266358 198056 266364
rect 198108 266354 198136 292839
rect 198568 282985 198596 304982
rect 198554 282976 198610 282985
rect 198554 282911 198610 282920
rect 198660 278089 198688 309198
rect 199396 294545 199424 319466
rect 199488 302190 199516 322079
rect 199476 302184 199528 302190
rect 199476 302126 199528 302132
rect 200776 301345 200804 342207
rect 201408 302184 201460 302190
rect 201408 302126 201460 302132
rect 200118 301336 200174 301345
rect 200118 301271 200174 301280
rect 200762 301336 200818 301345
rect 200762 301271 200818 301280
rect 199382 294536 199438 294545
rect 199382 294471 199438 294480
rect 198738 287328 198794 287337
rect 198738 287263 198794 287272
rect 198752 283529 198780 287263
rect 199474 287192 199530 287201
rect 199474 287127 199530 287136
rect 199384 285796 199436 285802
rect 199384 285738 199436 285744
rect 198738 283520 198794 283529
rect 198738 283455 198794 283464
rect 198646 278080 198702 278089
rect 198646 278015 198702 278024
rect 198646 274544 198702 274553
rect 198646 274479 198702 274488
rect 198096 266348 198148 266354
rect 198096 266290 198148 266296
rect 198094 262304 198150 262313
rect 198094 262239 198150 262248
rect 197358 258703 197414 258712
rect 197912 258732 197964 258738
rect 197912 258674 197964 258680
rect 197358 257952 197414 257961
rect 197358 257887 197414 257896
rect 197372 256834 197400 257887
rect 197360 256828 197412 256834
rect 197360 256770 197412 256776
rect 197360 256692 197412 256698
rect 197360 256634 197412 256640
rect 197372 255785 197400 256634
rect 197358 255776 197414 255785
rect 197358 255711 197414 255720
rect 197358 254416 197414 254425
rect 197358 254351 197414 254360
rect 197372 253978 197400 254351
rect 197360 253972 197412 253978
rect 197360 253914 197412 253920
rect 197450 253600 197506 253609
rect 197450 253535 197506 253544
rect 197358 253056 197414 253065
rect 197358 252991 197414 253000
rect 197372 252618 197400 252991
rect 197464 252686 197492 253535
rect 197452 252680 197504 252686
rect 197452 252622 197504 252628
rect 197360 252612 197412 252618
rect 197360 252554 197412 252560
rect 197358 252240 197414 252249
rect 197358 252175 197414 252184
rect 197372 251258 197400 252175
rect 197452 251864 197504 251870
rect 197452 251806 197504 251812
rect 197464 251705 197492 251806
rect 197450 251696 197506 251705
rect 197450 251631 197506 251640
rect 197360 251252 197412 251258
rect 197360 251194 197412 251200
rect 197358 250880 197414 250889
rect 197358 250815 197414 250824
rect 197372 249898 197400 250815
rect 197360 249892 197412 249898
rect 197360 249834 197412 249840
rect 197360 249756 197412 249762
rect 197360 249698 197412 249704
rect 197372 249529 197400 249698
rect 197358 249520 197414 249529
rect 197358 249455 197414 249464
rect 197450 247888 197506 247897
rect 197450 247823 197506 247832
rect 197464 247110 197492 247823
rect 197452 247104 197504 247110
rect 197452 247046 197504 247052
rect 197360 247036 197412 247042
rect 197360 246978 197412 246984
rect 197372 245993 197400 246978
rect 197358 245984 197414 245993
rect 197358 245919 197414 245928
rect 197360 245200 197412 245206
rect 197358 245168 197360 245177
rect 197412 245168 197414 245177
rect 197358 245103 197414 245112
rect 196714 243808 196770 243817
rect 196714 243743 196770 243752
rect 196622 235648 196678 235657
rect 196622 235583 196678 235592
rect 195886 229120 195942 229129
rect 195886 229055 195942 229064
rect 195796 228404 195848 228410
rect 195796 228346 195848 228352
rect 195612 224868 195664 224874
rect 195612 224810 195664 224816
rect 196728 224641 196756 243743
rect 197360 242208 197412 242214
rect 197266 242176 197322 242185
rect 197360 242150 197412 242156
rect 197266 242111 197322 242120
rect 196714 224632 196770 224641
rect 196714 224567 196770 224576
rect 196622 221504 196678 221513
rect 196622 221439 196678 221448
rect 196254 212528 196310 212537
rect 196254 212463 196310 212472
rect 196268 211857 196296 212463
rect 196254 211848 196310 211857
rect 196254 211783 196310 211792
rect 195242 204983 195298 204992
rect 195336 205012 195388 205018
rect 194508 189780 194560 189786
rect 194508 189722 194560 189728
rect 193864 177336 193916 177342
rect 193864 177278 193916 177284
rect 192668 175160 192720 175166
rect 192668 175102 192720 175108
rect 192576 168360 192628 168366
rect 192576 168302 192628 168308
rect 192576 153332 192628 153338
rect 192576 153274 192628 153280
rect 192484 138032 192536 138038
rect 192484 137974 192536 137980
rect 191288 94512 191340 94518
rect 191288 94454 191340 94460
rect 191194 89040 191250 89049
rect 191194 88975 191250 88984
rect 191104 64796 191156 64802
rect 191104 64738 191156 64744
rect 189724 60716 189776 60722
rect 189724 60658 189776 60664
rect 191300 53786 191328 94454
rect 191288 53780 191340 53786
rect 191288 53722 191340 53728
rect 192496 51066 192524 137974
rect 192588 73166 192616 153274
rect 194508 152516 194560 152522
rect 194508 152458 194560 152464
rect 194520 150414 194548 152458
rect 194508 150408 194560 150414
rect 194508 150350 194560 150356
rect 193864 142860 193916 142866
rect 193864 142802 193916 142808
rect 192668 108316 192720 108322
rect 192668 108258 192720 108264
rect 192680 87650 192708 108258
rect 192668 87644 192720 87650
rect 192668 87586 192720 87592
rect 192576 73160 192628 73166
rect 192576 73102 192628 73108
rect 192484 51060 192536 51066
rect 192484 51002 192536 51008
rect 188528 24200 188580 24206
rect 188528 24142 188580 24148
rect 193876 15881 193904 142802
rect 193956 120216 194008 120222
rect 193956 120158 194008 120164
rect 193968 85474 193996 120158
rect 193956 85468 194008 85474
rect 193956 85410 194008 85416
rect 195256 84862 195284 204983
rect 195336 204954 195388 204960
rect 195336 183592 195388 183598
rect 195336 183534 195388 183540
rect 195348 161362 195376 183534
rect 195336 161356 195388 161362
rect 195336 161298 195388 161304
rect 195336 127016 195388 127022
rect 195336 126958 195388 126964
rect 195244 84856 195296 84862
rect 195244 84798 195296 84804
rect 195244 82136 195296 82142
rect 195244 82078 195296 82084
rect 195256 15978 195284 82078
rect 195348 80034 195376 126958
rect 195336 80028 195388 80034
rect 195336 79970 195388 79976
rect 195244 15972 195296 15978
rect 195244 15914 195296 15920
rect 193862 15872 193918 15881
rect 193862 15807 193918 15816
rect 188342 13016 188398 13025
rect 188342 12951 188398 12960
rect 186964 8968 187016 8974
rect 186964 8910 187016 8916
rect 180156 4888 180208 4894
rect 178682 4856 178738 4865
rect 180156 4830 180208 4836
rect 178682 4791 178738 4800
rect 196636 3369 196664 221439
rect 197280 211857 197308 242111
rect 197372 241641 197400 242150
rect 198108 241777 198136 262239
rect 198660 257514 198688 274479
rect 199396 261594 199424 285738
rect 199384 261588 199436 261594
rect 199384 261530 199436 261536
rect 198648 257508 198700 257514
rect 198648 257450 198700 257456
rect 199384 257508 199436 257514
rect 199384 257450 199436 257456
rect 198646 256592 198702 256601
rect 198646 256527 198702 256536
rect 198094 241768 198150 241777
rect 198094 241703 198150 241712
rect 197358 241632 197414 241641
rect 197358 241567 197414 241576
rect 198004 217320 198056 217326
rect 198004 217262 198056 217268
rect 197358 214024 197414 214033
rect 197358 213959 197414 213968
rect 197372 213314 197400 213959
rect 197360 213308 197412 213314
rect 197360 213250 197412 213256
rect 197266 211848 197322 211857
rect 197266 211783 197322 211792
rect 196714 198248 196770 198257
rect 196714 198183 196770 198192
rect 196728 189689 196756 198183
rect 196714 189680 196770 189689
rect 196714 189615 196770 189624
rect 198016 181529 198044 217262
rect 198002 181520 198058 181529
rect 198002 181455 198058 181464
rect 198004 179920 198056 179926
rect 198004 179862 198056 179868
rect 197360 178764 197412 178770
rect 197360 178706 197412 178712
rect 197372 177993 197400 178706
rect 197358 177984 197414 177993
rect 197358 177919 197414 177928
rect 196808 128376 196860 128382
rect 196808 128318 196860 128324
rect 196820 86873 196848 128318
rect 196806 86864 196862 86873
rect 196806 86799 196862 86808
rect 196716 86284 196768 86290
rect 196716 86226 196768 86232
rect 196728 20058 196756 86226
rect 198016 39273 198044 179862
rect 198108 178673 198136 241703
rect 198660 241369 198688 256527
rect 198740 245064 198792 245070
rect 198740 245006 198792 245012
rect 198646 241360 198702 241369
rect 198646 241295 198702 241304
rect 198660 240174 198688 241295
rect 198648 240168 198700 240174
rect 198648 240110 198700 240116
rect 198752 239494 198780 245006
rect 198740 239488 198792 239494
rect 198740 239430 198792 239436
rect 198832 235272 198884 235278
rect 198832 235214 198884 235220
rect 198738 231976 198794 231985
rect 198738 231911 198794 231920
rect 198752 231130 198780 231911
rect 198740 231124 198792 231130
rect 198740 231066 198792 231072
rect 198844 230382 198872 235214
rect 198832 230376 198884 230382
rect 198832 230318 198884 230324
rect 198738 202464 198794 202473
rect 198738 202399 198794 202408
rect 198752 200122 198780 202399
rect 198740 200116 198792 200122
rect 198740 200058 198792 200064
rect 199396 193866 199424 257450
rect 199488 249801 199516 287127
rect 199566 285696 199622 285705
rect 199566 285631 199622 285640
rect 199580 273873 199608 285631
rect 200132 285326 200160 301271
rect 201420 300898 201448 302126
rect 201408 300892 201460 300898
rect 201408 300834 201460 300840
rect 201420 296714 201448 300834
rect 201328 296686 201448 296714
rect 200396 291168 200448 291174
rect 200396 291110 200448 291116
rect 200120 285320 200172 285326
rect 200120 285262 200172 285268
rect 200026 284608 200082 284617
rect 200026 284543 200082 284552
rect 199658 284472 199714 284481
rect 199658 284407 199714 284416
rect 199672 275398 199700 284407
rect 200040 282713 200068 284543
rect 200408 284172 200436 291110
rect 200488 285320 200540 285326
rect 200488 285262 200540 285268
rect 200500 284186 200528 285262
rect 200500 284158 200790 284186
rect 201328 284172 201356 296686
rect 201512 296041 201540 445742
rect 582392 432614 582420 484599
rect 582654 471472 582710 471481
rect 582654 471407 582710 471416
rect 582470 458144 582526 458153
rect 582470 458079 582526 458088
rect 582484 449206 582512 458079
rect 582472 449200 582524 449206
rect 582472 449142 582524 449148
rect 582380 432608 582432 432614
rect 582380 432550 582432 432556
rect 582378 431624 582434 431633
rect 582378 431559 582434 431568
rect 582392 403646 582420 431559
rect 582470 418296 582526 418305
rect 582470 418231 582526 418240
rect 582380 403640 582432 403646
rect 582380 403582 582432 403588
rect 242164 374128 242216 374134
rect 242164 374070 242216 374076
rect 215392 368620 215444 368626
rect 215392 368562 215444 368568
rect 209044 367124 209096 367130
rect 209044 367066 209096 367072
rect 204904 364472 204956 364478
rect 204904 364414 204956 364420
rect 204258 361856 204314 361865
rect 204258 361791 204314 361800
rect 202786 329080 202842 329089
rect 202786 329015 202842 329024
rect 201684 307828 201736 307834
rect 201684 307770 201736 307776
rect 201498 296032 201554 296041
rect 201498 295967 201554 295976
rect 201408 291848 201460 291854
rect 201408 291790 201460 291796
rect 201420 291553 201448 291790
rect 201406 291544 201462 291553
rect 201406 291479 201462 291488
rect 201696 284172 201724 307770
rect 202234 288552 202290 288561
rect 202234 288487 202290 288496
rect 202248 285705 202276 288487
rect 202234 285696 202290 285705
rect 202234 285631 202290 285640
rect 202248 284172 202276 285631
rect 202800 284172 202828 329015
rect 204272 291174 204300 361791
rect 204352 343664 204404 343670
rect 204352 343606 204404 343612
rect 204364 306374 204392 343606
rect 204916 320958 204944 364414
rect 208124 363656 208176 363662
rect 208124 363598 208176 363604
rect 206282 352200 206338 352209
rect 206282 352135 206338 352144
rect 204904 320952 204956 320958
rect 204904 320894 204956 320900
rect 204364 306346 204760 306374
rect 204260 291168 204312 291174
rect 204260 291110 204312 291116
rect 203154 288824 203210 288833
rect 203154 288759 203210 288768
rect 203168 284172 203196 288759
rect 203706 287192 203762 287201
rect 203706 287127 203762 287136
rect 203720 284172 203748 287127
rect 204628 285728 204680 285734
rect 204628 285670 204680 285676
rect 204258 284336 204314 284345
rect 204258 284271 204314 284280
rect 204272 284172 204300 284271
rect 204640 284172 204668 285670
rect 204732 283914 204760 306346
rect 206296 295361 206324 352135
rect 206376 335368 206428 335374
rect 206376 335310 206428 335316
rect 206282 295352 206338 295361
rect 206282 295287 206338 295296
rect 206098 287464 206154 287473
rect 206098 287399 206154 287408
rect 205548 285796 205600 285802
rect 205548 285738 205600 285744
rect 205560 284172 205588 285738
rect 206112 284172 206140 287399
rect 206388 285734 206416 335310
rect 207662 334248 207718 334257
rect 207662 334183 207718 334192
rect 207676 307902 207704 334183
rect 207664 307896 207716 307902
rect 207664 307838 207716 307844
rect 207676 296714 207704 307838
rect 207584 296686 207704 296714
rect 206650 295352 206706 295361
rect 206650 295287 206706 295296
rect 206376 285728 206428 285734
rect 206376 285670 206428 285676
rect 206664 284172 206692 295287
rect 207020 285728 207072 285734
rect 207020 285670 207072 285676
rect 205362 283928 205418 283937
rect 204732 283886 205362 283914
rect 207032 283914 207060 285670
rect 207584 284172 207612 296686
rect 208136 284172 208164 363598
rect 208490 332752 208546 332761
rect 208490 332687 208546 332696
rect 208400 300960 208452 300966
rect 208400 300902 208452 300908
rect 208412 285326 208440 300902
rect 208400 285320 208452 285326
rect 208400 285262 208452 285268
rect 207110 283928 207166 283937
rect 207032 283900 207110 283914
rect 207046 283886 207110 283900
rect 205362 283863 205418 283872
rect 208504 283914 208532 332687
rect 209056 287201 209084 367066
rect 214564 360256 214616 360262
rect 214564 360198 214616 360204
rect 213184 358828 213236 358834
rect 213184 358770 213236 358776
rect 211804 343732 211856 343738
rect 211804 343674 211856 343680
rect 209134 339688 209190 339697
rect 209134 339623 209190 339632
rect 209148 298353 209176 339623
rect 210424 319456 210476 319462
rect 210424 319398 210476 319404
rect 210436 318850 210464 319398
rect 210424 318844 210476 318850
rect 210424 318786 210476 318792
rect 210436 316034 210464 318786
rect 210436 316006 210556 316034
rect 209134 298344 209190 298353
rect 209134 298279 209190 298288
rect 209410 298344 209466 298353
rect 209410 298279 209466 298288
rect 209042 287192 209098 287201
rect 209042 287127 209098 287136
rect 208676 285320 208728 285326
rect 208676 285262 208728 285268
rect 208688 284186 208716 285262
rect 208688 284158 209070 284186
rect 209424 284172 209452 298279
rect 210422 296032 210478 296041
rect 210422 295967 210478 295976
rect 210436 289785 210464 295967
rect 210422 289776 210478 289785
rect 210422 289711 210478 289720
rect 210436 287054 210464 289711
rect 210344 287026 210464 287054
rect 210344 284186 210372 287026
rect 209990 284158 210372 284186
rect 210528 284172 210556 316006
rect 211816 306474 211844 343674
rect 213196 327826 213224 358770
rect 213184 327820 213236 327826
rect 213184 327762 213236 327768
rect 212906 327312 212962 327321
rect 212906 327247 212962 327256
rect 211894 315344 211950 315353
rect 211894 315279 211950 315288
rect 211804 306468 211856 306474
rect 211804 306410 211856 306416
rect 211816 296714 211844 306410
rect 211908 306374 211936 315279
rect 211908 306346 212120 306374
rect 211448 296686 211844 296714
rect 210882 285968 210938 285977
rect 210882 285903 210938 285912
rect 210896 284172 210924 285903
rect 211448 284172 211476 296686
rect 211986 287192 212042 287201
rect 211986 287127 212042 287136
rect 212000 284617 212028 287127
rect 211986 284608 212042 284617
rect 211986 284543 212042 284552
rect 212000 284172 212028 284543
rect 212092 284186 212120 306346
rect 212354 284336 212410 284345
rect 212354 284271 212410 284280
rect 212368 284186 212396 284271
rect 212092 284172 212396 284186
rect 212920 284172 212948 327247
rect 214576 311234 214604 360198
rect 214654 351112 214710 351121
rect 214654 351047 214710 351056
rect 214564 311228 214616 311234
rect 214564 311170 214616 311176
rect 214668 306374 214696 351047
rect 214668 306346 214788 306374
rect 214760 303686 214788 306346
rect 213184 303680 213236 303686
rect 213184 303622 213236 303628
rect 214748 303680 214800 303686
rect 214748 303622 214800 303628
rect 213196 293282 213224 303622
rect 213184 293276 213236 293282
rect 213184 293218 213236 293224
rect 213182 291816 213238 291825
rect 213182 291751 213238 291760
rect 213196 286385 213224 291751
rect 213182 286376 213238 286385
rect 213182 286311 213238 286320
rect 213196 284186 213224 286311
rect 213828 285796 213880 285802
rect 213828 285738 213880 285744
rect 212092 284158 212382 284172
rect 213196 284158 213486 284186
rect 213840 284172 213868 285738
rect 214564 285728 214616 285734
rect 214564 285670 214616 285676
rect 214576 284986 214604 285670
rect 214564 284980 214616 284986
rect 214564 284922 214616 284928
rect 214760 284172 214788 303622
rect 215298 298072 215354 298081
rect 215298 298007 215354 298016
rect 215312 296993 215340 298007
rect 215298 296984 215354 296993
rect 215298 296919 215354 296928
rect 215312 284172 215340 296919
rect 215404 285802 215432 368562
rect 218242 365936 218298 365945
rect 218242 365871 218298 365880
rect 216034 337104 216090 337113
rect 216034 337039 216090 337048
rect 215944 331288 215996 331294
rect 215944 331230 215996 331236
rect 215850 311944 215906 311953
rect 215850 311879 215906 311888
rect 215392 285796 215444 285802
rect 215392 285738 215444 285744
rect 215864 284172 215892 311879
rect 215956 298081 215984 331230
rect 216048 311953 216076 337039
rect 217322 331256 217378 331265
rect 217322 331191 217378 331200
rect 217336 314702 217364 331191
rect 217324 314696 217376 314702
rect 217324 314638 217376 314644
rect 217968 314696 218020 314702
rect 217968 314638 218020 314644
rect 216034 311944 216090 311953
rect 216034 311879 216090 311888
rect 215942 298072 215998 298081
rect 215942 298007 215998 298016
rect 217876 291304 217928 291310
rect 217874 291272 217876 291281
rect 217928 291272 217930 291281
rect 217874 291207 217930 291216
rect 216770 288688 216826 288697
rect 216770 288623 216826 288632
rect 216784 284442 216812 288623
rect 217980 286482 218008 314638
rect 218060 291848 218112 291854
rect 218060 291790 218112 291796
rect 218072 291281 218100 291790
rect 218152 291304 218204 291310
rect 218058 291272 218114 291281
rect 218152 291246 218204 291252
rect 218058 291207 218114 291216
rect 217968 286476 218020 286482
rect 217968 286418 218020 286424
rect 218164 285326 218192 291246
rect 218152 285320 218204 285326
rect 218152 285262 218204 285268
rect 217322 284472 217378 284481
rect 216772 284436 216824 284442
rect 217322 284407 217378 284416
rect 216772 284378 216824 284384
rect 216784 284172 216812 284378
rect 217336 284172 217364 284407
rect 218256 284172 218284 365871
rect 227442 364440 227498 364449
rect 227442 364375 227498 364384
rect 240508 364404 240560 364410
rect 225604 356108 225656 356114
rect 225604 356050 225656 356056
rect 222936 353388 222988 353394
rect 222936 353330 222988 353336
rect 218704 353320 218756 353326
rect 218704 353262 218756 353268
rect 218716 296857 218744 353262
rect 221464 346452 221516 346458
rect 221464 346394 221516 346400
rect 220084 342372 220136 342378
rect 220084 342314 220136 342320
rect 220096 302326 220124 342314
rect 220174 336968 220230 336977
rect 220174 336903 220230 336912
rect 220188 305017 220216 336903
rect 221476 306374 221504 346394
rect 222842 338192 222898 338201
rect 222842 338127 222898 338136
rect 221200 306346 221504 306374
rect 220174 305008 220230 305017
rect 220174 304943 220230 304952
rect 221200 303754 221228 306346
rect 222106 305008 222162 305017
rect 222106 304943 222162 304952
rect 221188 303748 221240 303754
rect 221188 303690 221240 303696
rect 220084 302320 220136 302326
rect 220084 302262 220136 302268
rect 220728 302320 220780 302326
rect 220728 302262 220780 302268
rect 218702 296848 218758 296857
rect 218702 296783 218758 296792
rect 220636 292596 220688 292602
rect 220636 292538 220688 292544
rect 219162 285968 219218 285977
rect 219162 285903 219218 285912
rect 218336 285320 218388 285326
rect 218336 285262 218388 285268
rect 218348 284186 218376 285262
rect 218348 284158 218638 284186
rect 219176 284172 219204 285903
rect 219716 285728 219768 285734
rect 219716 285670 219768 285676
rect 220082 285696 220138 285705
rect 219728 284172 219756 285670
rect 220082 285631 220138 285640
rect 220096 284172 220124 285631
rect 220648 284172 220676 292538
rect 220740 285734 220768 302262
rect 220728 285728 220780 285734
rect 220728 285670 220780 285676
rect 221200 284172 221228 303690
rect 221556 286476 221608 286482
rect 221556 286418 221608 286424
rect 221568 284172 221596 286418
rect 222120 284172 222148 304943
rect 222474 289640 222530 289649
rect 222474 289575 222530 289584
rect 222488 288697 222516 289575
rect 222474 288688 222530 288697
rect 222474 288623 222530 288632
rect 222488 284172 222516 288623
rect 222856 285734 222884 338127
rect 222948 321026 222976 353330
rect 223946 349208 224002 349217
rect 223946 349143 224002 349152
rect 222936 321020 222988 321026
rect 222936 320962 222988 320968
rect 223028 320884 223080 320890
rect 223028 320826 223080 320832
rect 223040 289649 223068 320826
rect 223026 289640 223082 289649
rect 223026 289575 223082 289584
rect 223026 287328 223082 287337
rect 223026 287263 223082 287272
rect 222844 285728 222896 285734
rect 222844 285670 222896 285676
rect 223040 284172 223068 287263
rect 223580 285796 223632 285802
rect 223580 285738 223632 285744
rect 223592 284172 223620 285738
rect 223960 284172 223988 349143
rect 224224 329112 224276 329118
rect 224224 329054 224276 329060
rect 224236 286278 224264 329054
rect 225328 298784 225380 298790
rect 225328 298726 225380 298732
rect 225340 292641 225368 298726
rect 225616 295497 225644 356050
rect 226430 331392 226486 331401
rect 226430 331327 226486 331336
rect 226444 306374 226472 331327
rect 226444 306346 226656 306374
rect 225418 295488 225474 295497
rect 225418 295423 225474 295432
rect 225602 295488 225658 295497
rect 225602 295423 225658 295432
rect 225326 292632 225382 292641
rect 225326 292567 225382 292576
rect 224500 288448 224552 288454
rect 224500 288390 224552 288396
rect 224224 286272 224276 286278
rect 224224 286214 224276 286220
rect 208674 283928 208730 283937
rect 208504 283900 208674 283914
rect 208518 283886 208674 283900
rect 207110 283863 207166 283872
rect 208674 283863 208730 283872
rect 214102 283928 214158 283937
rect 215942 283928 215998 283937
rect 214158 283886 214406 283914
rect 214102 283863 214158 283872
rect 217414 283928 217470 283937
rect 215998 283886 216246 283914
rect 215942 283863 215998 283872
rect 224512 283914 224540 288390
rect 225052 286272 225104 286278
rect 225052 286214 225104 286220
rect 225064 285841 225092 286214
rect 225050 285832 225106 285841
rect 225050 285767 225106 285776
rect 225064 284172 225092 285767
rect 225432 284172 225460 295423
rect 225970 294536 226026 294545
rect 225970 294471 226026 294480
rect 225984 284172 226012 294471
rect 226522 286104 226578 286113
rect 226522 286039 226578 286048
rect 226536 285734 226564 286039
rect 226524 285728 226576 285734
rect 226524 285670 226576 285676
rect 226536 284172 226564 285670
rect 226628 283937 226656 306346
rect 227456 284172 227484 364375
rect 240508 364346 240560 364352
rect 238022 363080 238078 363089
rect 238022 363015 238078 363024
rect 232502 361720 232558 361729
rect 232502 361655 232558 361664
rect 228362 359000 228418 359009
rect 228362 358935 228418 358944
rect 227628 318164 227680 318170
rect 227628 318106 227680 318112
rect 227640 310593 227668 318106
rect 227812 311228 227864 311234
rect 227812 311170 227864 311176
rect 227626 310584 227682 310593
rect 227626 310519 227682 310528
rect 227640 285802 227668 310519
rect 227628 285796 227680 285802
rect 227628 285738 227680 285744
rect 224682 283928 224738 283937
rect 217470 283886 217718 283914
rect 224512 283900 224682 283914
rect 224526 283886 224682 283900
rect 217414 283863 217470 283872
rect 224682 283863 224738 283872
rect 226614 283928 226670 283937
rect 227824 283914 227852 311170
rect 228376 298790 228404 358935
rect 231124 345160 231176 345166
rect 231124 345102 231176 345108
rect 228456 335436 228508 335442
rect 228456 335378 228508 335384
rect 228364 298784 228416 298790
rect 228364 298726 228416 298732
rect 228362 292632 228418 292641
rect 228362 292567 228418 292576
rect 228376 284172 228404 292567
rect 228468 285734 228496 335378
rect 230386 330440 230442 330449
rect 230386 330375 230442 330384
rect 229742 295488 229798 295497
rect 229742 295423 229798 295432
rect 229756 287473 229784 295423
rect 229742 287464 229798 287473
rect 229742 287399 229798 287408
rect 228916 285796 228968 285802
rect 228916 285738 228968 285744
rect 228456 285728 228508 285734
rect 228456 285670 228508 285676
rect 228928 284172 228956 285738
rect 229284 285728 229336 285734
rect 229284 285670 229336 285676
rect 227994 283928 228050 283937
rect 226670 283886 226918 283914
rect 227824 283900 227994 283914
rect 227838 283886 227994 283900
rect 226614 283863 226670 283872
rect 229296 283914 229324 285670
rect 229756 284186 229784 287399
rect 229756 284158 229862 284186
rect 230400 284172 230428 330375
rect 230480 312656 230532 312662
rect 230480 312598 230532 312604
rect 230492 284481 230520 312598
rect 230572 288516 230624 288522
rect 230572 288458 230624 288464
rect 230584 285977 230612 288458
rect 230570 285968 230626 285977
rect 230570 285903 230626 285912
rect 230478 284472 230534 284481
rect 230478 284407 230534 284416
rect 230584 284186 230612 285903
rect 231136 285802 231164 345102
rect 232516 289814 232544 361655
rect 233882 356144 233938 356153
rect 233882 356079 233938 356088
rect 233698 296848 233754 296857
rect 233698 296783 233754 296792
rect 232778 291408 232834 291417
rect 232778 291343 232834 291352
rect 232504 289808 232556 289814
rect 232504 289750 232556 289756
rect 231308 287156 231360 287162
rect 231308 287098 231360 287104
rect 231124 285796 231176 285802
rect 231124 285738 231176 285744
rect 230584 284158 230782 284186
rect 229466 283928 229522 283937
rect 229296 283900 229466 283914
rect 229310 283886 229466 283900
rect 227994 283863 228050 283872
rect 231320 283914 231348 287098
rect 232228 285796 232280 285802
rect 232228 285738 232280 285744
rect 231674 284472 231730 284481
rect 231674 284407 231730 284416
rect 231688 284172 231716 284407
rect 232240 284172 232268 285738
rect 232792 284172 232820 291343
rect 233712 291145 233740 296783
rect 233896 292641 233924 356079
rect 235264 347880 235316 347886
rect 235264 347822 235316 347828
rect 233976 311160 234028 311166
rect 233976 311102 234028 311108
rect 233882 292632 233938 292641
rect 233882 292567 233938 292576
rect 233698 291136 233754 291145
rect 233698 291071 233754 291080
rect 233148 285728 233200 285734
rect 233148 285670 233200 285676
rect 233160 284172 233188 285670
rect 233712 284172 233740 291071
rect 233896 285734 233924 292567
rect 233988 291310 234016 311102
rect 235276 306374 235304 347822
rect 236644 339516 236696 339522
rect 236644 339458 236696 339464
rect 235540 314016 235592 314022
rect 235540 313958 235592 313964
rect 235184 306346 235304 306374
rect 235184 302433 235212 306346
rect 235170 302424 235226 302433
rect 235170 302359 235226 302368
rect 233976 291304 234028 291310
rect 233976 291246 234028 291252
rect 233884 285728 233936 285734
rect 233884 285670 233936 285676
rect 233988 284186 234016 291246
rect 234620 289808 234672 289814
rect 234620 289750 234672 289756
rect 233988 284158 234278 284186
rect 234632 284172 234660 289750
rect 235184 284172 235212 302359
rect 235552 284172 235580 313958
rect 236184 298784 236236 298790
rect 236184 298726 236236 298732
rect 236196 298178 236224 298726
rect 236184 298172 236236 298178
rect 236184 298114 236236 298120
rect 236092 297356 236144 297362
rect 236092 297298 236144 297304
rect 236000 293276 236052 293282
rect 236000 293218 236052 293224
rect 236012 285705 236040 293218
rect 235998 285696 236054 285705
rect 235998 285631 236054 285640
rect 236104 284172 236132 297298
rect 236196 284186 236224 298114
rect 236656 297362 236684 339458
rect 236644 297356 236696 297362
rect 236644 297298 236696 297304
rect 236656 296818 236684 297298
rect 236644 296812 236696 296818
rect 236644 296754 236696 296760
rect 238036 294001 238064 363015
rect 239402 336016 239458 336025
rect 239402 335951 239458 335960
rect 238116 320952 238168 320958
rect 238116 320894 238168 320900
rect 238022 293992 238078 294001
rect 238022 293927 238078 293936
rect 238128 288454 238156 320894
rect 238484 296744 238536 296750
rect 238484 296686 238536 296692
rect 237932 288448 237984 288454
rect 237932 288390 237984 288396
rect 238116 288448 238168 288454
rect 238116 288390 238168 288396
rect 237944 284186 237972 288390
rect 238116 287156 238168 287162
rect 238116 287098 238168 287104
rect 236196 284158 236670 284186
rect 237590 284158 237972 284186
rect 238128 284172 238156 287098
rect 238496 284172 238524 296686
rect 239034 293992 239090 294001
rect 239034 293927 239090 293936
rect 239048 284172 239076 293927
rect 239416 291106 239444 335951
rect 239496 330540 239548 330546
rect 239496 330482 239548 330488
rect 239404 291100 239456 291106
rect 239404 291042 239456 291048
rect 239508 290057 239536 330482
rect 239956 290488 240008 290494
rect 239956 290430 240008 290436
rect 239494 290048 239550 290057
rect 239494 289983 239550 289992
rect 239508 284186 239536 289983
rect 239968 287337 239996 290430
rect 239954 287328 240010 287337
rect 239954 287263 240010 287272
rect 239508 284158 239614 284186
rect 239968 284172 239996 287263
rect 240520 284172 240548 364346
rect 241520 357468 241572 357474
rect 241520 357410 241572 357416
rect 240784 325780 240836 325786
rect 240784 325722 240836 325728
rect 240796 286550 240824 325722
rect 241532 300801 241560 357410
rect 240874 300792 240930 300801
rect 240874 300727 240930 300736
rect 241518 300792 241574 300801
rect 241518 300727 241574 300736
rect 240888 300121 240916 300727
rect 240874 300112 240930 300121
rect 240874 300047 240930 300056
rect 240784 286544 240836 286550
rect 240784 286486 240836 286492
rect 240888 284172 240916 300047
rect 241426 294128 241482 294137
rect 241426 294063 241482 294072
rect 241440 284172 241468 294063
rect 242176 289814 242204 374070
rect 248512 372632 248564 372638
rect 248512 372574 248564 372580
rect 247316 336796 247368 336802
rect 247316 336738 247368 336744
rect 243820 321632 243872 321638
rect 243820 321574 243872 321580
rect 242256 318096 242308 318102
rect 242256 318038 242308 318044
rect 242164 289808 242216 289814
rect 242164 289750 242216 289756
rect 241980 286544 242032 286550
rect 241980 286486 242032 286492
rect 231582 283928 231638 283937
rect 231320 283900 231582 283914
rect 231334 283886 231582 283900
rect 229466 283863 229522 283872
rect 231582 283863 231638 283872
rect 236734 283928 236790 283937
rect 241992 283914 242020 286486
rect 242268 285841 242296 318038
rect 242348 291100 242400 291106
rect 242348 291042 242400 291048
rect 242360 289882 242388 291042
rect 242348 289876 242400 289882
rect 242348 289818 242400 289824
rect 242254 285832 242310 285841
rect 242254 285767 242310 285776
rect 242360 284172 242388 289818
rect 242900 289808 242952 289814
rect 242900 289750 242952 289756
rect 242912 284172 242940 289750
rect 243450 285832 243506 285841
rect 243450 285767 243506 285776
rect 243464 284050 243492 285767
rect 243832 284172 243860 321574
rect 244280 315308 244332 315314
rect 244280 315250 244332 315256
rect 244004 302252 244056 302258
rect 244004 302194 244056 302200
rect 243634 284064 243690 284073
rect 243464 284036 243634 284050
rect 243478 284022 243634 284036
rect 243634 283999 243690 284008
rect 242256 283960 242308 283966
rect 236790 283886 237038 283914
rect 241992 283908 242256 283914
rect 241992 283902 242308 283908
rect 241992 283900 242296 283902
rect 242006 283886 242296 283900
rect 236734 283863 236790 283872
rect 200026 282704 200082 282713
rect 200026 282639 200082 282648
rect 199660 275392 199712 275398
rect 199660 275334 199712 275340
rect 199566 273864 199622 273873
rect 199566 273799 199622 273808
rect 244016 271289 244044 302194
rect 244094 284064 244150 284073
rect 244094 283999 244150 284008
rect 244108 282985 244136 283999
rect 244094 282976 244150 282985
rect 244094 282911 244150 282920
rect 244292 278089 244320 315250
rect 245660 312588 245712 312594
rect 245660 312530 245712 312536
rect 244924 299532 244976 299538
rect 244924 299474 244976 299480
rect 244372 295996 244424 296002
rect 244372 295938 244424 295944
rect 244278 278080 244334 278089
rect 244278 278015 244334 278024
rect 244002 271280 244058 271289
rect 244002 271215 244058 271224
rect 199568 264240 199620 264246
rect 199568 264182 199620 264188
rect 199474 249792 199530 249801
rect 199474 249727 199530 249736
rect 199488 249082 199516 249727
rect 199476 249076 199528 249082
rect 199476 249018 199528 249024
rect 199580 240281 199608 264182
rect 244384 259593 244412 295938
rect 244464 287088 244516 287094
rect 244464 287030 244516 287036
rect 244370 259584 244426 259593
rect 244370 259519 244426 259528
rect 244384 259486 244412 259519
rect 244372 259480 244424 259486
rect 244372 259422 244424 259428
rect 244476 258777 244504 287030
rect 244936 269113 244964 299474
rect 245672 274553 245700 312530
rect 245752 305652 245804 305658
rect 245752 305594 245804 305600
rect 245764 276729 245792 305594
rect 245842 300248 245898 300257
rect 245842 300183 245898 300192
rect 245750 276720 245806 276729
rect 245750 276655 245752 276664
rect 245804 276655 245806 276664
rect 245752 276626 245804 276632
rect 245764 276595 245792 276626
rect 245856 274666 245884 300183
rect 245936 294636 245988 294642
rect 245936 294578 245988 294584
rect 245948 287054 245976 294578
rect 247222 292768 247278 292777
rect 247222 292703 247278 292712
rect 247130 290184 247186 290193
rect 247130 290119 247186 290128
rect 245948 287026 246068 287054
rect 245934 282432 245990 282441
rect 245934 282367 245990 282376
rect 245948 281722 245976 282367
rect 245936 281716 245988 281722
rect 245936 281658 245988 281664
rect 245934 281072 245990 281081
rect 245934 281007 245990 281016
rect 245948 280838 245976 281007
rect 245936 280832 245988 280838
rect 245936 280774 245988 280780
rect 245936 279880 245988 279886
rect 245936 279822 245988 279828
rect 245948 279449 245976 279822
rect 245934 279440 245990 279449
rect 245934 279375 245990 279384
rect 245936 278724 245988 278730
rect 245936 278666 245988 278672
rect 245948 277545 245976 278666
rect 245934 277536 245990 277545
rect 245934 277471 245990 277480
rect 245936 276004 245988 276010
rect 245936 275946 245988 275952
rect 245948 275913 245976 275946
rect 245934 275904 245990 275913
rect 245934 275839 245990 275848
rect 245856 274638 245976 274666
rect 245658 274544 245714 274553
rect 245658 274479 245714 274488
rect 245842 274544 245898 274553
rect 245842 274479 245898 274488
rect 245856 273970 245884 274479
rect 245844 273964 245896 273970
rect 245844 273906 245896 273912
rect 245842 273728 245898 273737
rect 245842 273663 245898 273672
rect 245856 273290 245884 273663
rect 245844 273284 245896 273290
rect 245844 273226 245896 273232
rect 245750 273184 245806 273193
rect 245750 273119 245806 273128
rect 245764 272542 245792 273119
rect 245752 272536 245804 272542
rect 245752 272478 245804 272484
rect 245948 272377 245976 274638
rect 245934 272368 245990 272377
rect 245934 272303 245990 272312
rect 245842 271552 245898 271561
rect 245842 271487 245844 271496
rect 245896 271487 245898 271496
rect 245844 271458 245896 271464
rect 245936 270496 245988 270502
rect 245936 270438 245988 270444
rect 245948 270201 245976 270438
rect 245934 270192 245990 270201
rect 245934 270127 245990 270136
rect 246040 269657 246068 287026
rect 247040 284368 247092 284374
rect 247040 284310 247092 284316
rect 246396 283620 246448 283626
rect 246396 283562 246448 283568
rect 246408 283257 246436 283562
rect 246394 283248 246450 283257
rect 246394 283183 246450 283192
rect 246120 282872 246172 282878
rect 246120 282814 246172 282820
rect 246132 281625 246160 282814
rect 246118 281616 246174 281625
rect 246118 281551 246174 281560
rect 246120 281512 246172 281518
rect 246120 281454 246172 281460
rect 246132 280265 246160 281454
rect 246118 280256 246174 280265
rect 246118 280191 246174 280200
rect 246486 272368 246542 272377
rect 246486 272303 246542 272312
rect 246026 269648 246082 269657
rect 246026 269583 246082 269592
rect 244922 269104 244978 269113
rect 244922 269039 244978 269048
rect 245752 269068 245804 269074
rect 245752 269010 245804 269016
rect 245764 268025 245792 269010
rect 245750 268016 245806 268025
rect 245750 267951 245806 267960
rect 245842 267472 245898 267481
rect 245842 267407 245898 267416
rect 245856 266422 245884 267407
rect 245934 266656 245990 266665
rect 245934 266591 245990 266600
rect 245844 266416 245896 266422
rect 245844 266358 245896 266364
rect 245948 266354 245976 266591
rect 245936 266348 245988 266354
rect 245936 266290 245988 266296
rect 245934 265840 245990 265849
rect 245934 265775 245936 265784
rect 245988 265775 245990 265784
rect 245936 265746 245988 265752
rect 246040 264246 246068 269583
rect 246500 267034 246528 272303
rect 246580 269816 246632 269822
rect 246580 269758 246632 269764
rect 246488 267028 246540 267034
rect 246488 266970 246540 266976
rect 246592 265305 246620 269758
rect 246670 269104 246726 269113
rect 246670 269039 246726 269048
rect 246578 265296 246634 265305
rect 246578 265231 246634 265240
rect 246028 264240 246080 264246
rect 244922 264208 244978 264217
rect 246028 264182 246080 264188
rect 244922 264143 244978 264152
rect 244462 258768 244518 258777
rect 244462 258703 244518 258712
rect 200040 257446 200068 257477
rect 200028 257440 200080 257446
rect 200026 257408 200028 257417
rect 200080 257408 200082 257417
rect 200026 257343 200082 257352
rect 199934 240816 199990 240825
rect 199934 240751 199990 240760
rect 199566 240272 199622 240281
rect 199566 240207 199622 240216
rect 199948 235346 199976 240751
rect 199936 235340 199988 235346
rect 199936 235282 199988 235288
rect 200040 215966 200068 257343
rect 244278 250880 244334 250889
rect 244278 250815 244334 250824
rect 244002 243264 244058 243273
rect 243924 243222 244002 243250
rect 200120 240508 200172 240514
rect 200120 240450 200172 240456
rect 200132 239562 200160 240450
rect 200120 239556 200172 239562
rect 200120 239498 200172 239504
rect 200120 239420 200172 239426
rect 200120 239362 200172 239368
rect 200132 238649 200160 239362
rect 200224 238785 200252 240244
rect 200304 240168 200356 240174
rect 200304 240110 200356 240116
rect 200210 238776 200266 238785
rect 200210 238711 200266 238720
rect 200118 238640 200174 238649
rect 200118 238575 200174 238584
rect 200224 237425 200252 238711
rect 200210 237416 200266 237425
rect 200210 237351 200266 237360
rect 200316 234666 200344 240110
rect 200304 234660 200356 234666
rect 200304 234602 200356 234608
rect 200592 219434 200620 240244
rect 201144 240145 201172 240244
rect 201130 240136 201186 240145
rect 201130 240071 201186 240080
rect 201144 238754 201172 240071
rect 201144 238726 201448 238754
rect 200762 237416 200818 237425
rect 200762 237351 200818 237360
rect 200132 219406 200620 219434
rect 200028 215960 200080 215966
rect 200028 215902 200080 215908
rect 200132 207754 200160 219406
rect 200040 207726 200160 207754
rect 200040 207670 200068 207726
rect 200028 207664 200080 207670
rect 200028 207606 200080 207612
rect 200040 201482 200068 207606
rect 200028 201476 200080 201482
rect 200028 201418 200080 201424
rect 199384 193860 199436 193866
rect 199384 193802 199436 193808
rect 200776 184278 200804 237351
rect 200854 232656 200910 232665
rect 200854 232591 200910 232600
rect 200868 201414 200896 232591
rect 201420 225350 201448 238726
rect 201408 225344 201460 225350
rect 201408 225286 201460 225292
rect 201512 204241 201540 240244
rect 202064 237289 202092 240244
rect 202050 237280 202106 237289
rect 202050 237215 202106 237224
rect 202144 234660 202196 234666
rect 202144 234602 202196 234608
rect 201590 231160 201646 231169
rect 201590 231095 201646 231104
rect 201604 222902 201632 231095
rect 201592 222896 201644 222902
rect 201592 222838 201644 222844
rect 202156 221474 202184 234602
rect 202144 221468 202196 221474
rect 202144 221410 202196 221416
rect 201498 204232 201554 204241
rect 201498 204167 201554 204176
rect 202234 204232 202290 204241
rect 202234 204167 202290 204176
rect 200856 201408 200908 201414
rect 200856 201350 200908 201356
rect 202144 199436 202196 199442
rect 202144 199378 202196 199384
rect 200764 184272 200816 184278
rect 200764 184214 200816 184220
rect 200762 178936 200818 178945
rect 200762 178871 200818 178880
rect 198094 178664 198150 178673
rect 198094 178599 198150 178608
rect 198094 177168 198150 177177
rect 198094 177103 198150 177112
rect 198108 160002 198136 177103
rect 198096 159996 198148 160002
rect 198096 159938 198148 159944
rect 198188 145036 198240 145042
rect 198188 144978 198240 144984
rect 198094 105224 198150 105233
rect 198094 105159 198150 105168
rect 198108 89010 198136 105159
rect 198096 89004 198148 89010
rect 198096 88946 198148 88952
rect 198096 87644 198148 87650
rect 198096 87586 198148 87592
rect 198002 39264 198058 39273
rect 198002 39199 198058 39208
rect 196716 20052 196768 20058
rect 196716 19994 196768 20000
rect 196622 3360 196678 3369
rect 196622 3295 196678 3304
rect 198108 2174 198136 87586
rect 198200 62082 198228 144978
rect 199384 140072 199436 140078
rect 199384 140014 199436 140020
rect 198188 62076 198240 62082
rect 198188 62018 198240 62024
rect 199396 51814 199424 140014
rect 199476 116068 199528 116074
rect 199476 116010 199528 116016
rect 199488 90953 199516 116010
rect 199474 90944 199530 90953
rect 199474 90879 199530 90888
rect 199384 51808 199436 51814
rect 199384 51750 199436 51756
rect 200776 15978 200804 178871
rect 200856 138712 200908 138718
rect 200856 138654 200908 138660
rect 200764 15972 200816 15978
rect 200764 15914 200816 15920
rect 198096 2168 198148 2174
rect 198096 2110 198148 2116
rect 200868 2009 200896 138654
rect 202156 3534 202184 199378
rect 202248 195401 202276 204167
rect 202616 198801 202644 240244
rect 202786 236736 202842 236745
rect 202786 236671 202788 236680
rect 202840 236671 202842 236680
rect 202788 236642 202840 236648
rect 202984 219434 203012 240244
rect 203536 225010 203564 240244
rect 204088 233170 204116 240244
rect 204456 240009 204484 240244
rect 204442 240000 204498 240009
rect 204442 239935 204498 239944
rect 204166 239456 204222 239465
rect 204166 239391 204222 239400
rect 204180 236706 204208 239391
rect 205008 238754 205036 240244
rect 205008 238726 205128 238754
rect 205100 236745 205128 238726
rect 205086 236736 205142 236745
rect 204168 236700 204220 236706
rect 205086 236671 205142 236680
rect 204168 236642 204220 236648
rect 204996 235340 205048 235346
rect 204996 235282 205048 235288
rect 203616 233164 203668 233170
rect 203616 233106 203668 233112
rect 204076 233164 204128 233170
rect 204076 233106 204128 233112
rect 203628 228313 203656 233106
rect 203614 228304 203670 228313
rect 203614 228239 203670 228248
rect 203616 225344 203668 225350
rect 203616 225286 203668 225292
rect 203524 225004 203576 225010
rect 203524 224946 203576 224952
rect 203536 223553 203564 224946
rect 203522 223544 203578 223553
rect 203522 223479 203578 223488
rect 202892 219406 203012 219434
rect 202892 202774 202920 219406
rect 202880 202768 202932 202774
rect 202880 202710 202932 202716
rect 203524 202768 203576 202774
rect 203524 202710 203576 202716
rect 202602 198792 202658 198801
rect 202602 198727 202658 198736
rect 202234 195392 202290 195401
rect 202234 195327 202290 195336
rect 202616 191826 202644 198727
rect 202604 191820 202656 191826
rect 202604 191762 202656 191768
rect 203536 186969 203564 202710
rect 203522 186960 203578 186969
rect 203522 186895 203578 186904
rect 203628 182918 203656 225286
rect 204902 222048 204958 222057
rect 204902 221983 204958 221992
rect 204916 220969 204944 221983
rect 204902 220960 204958 220969
rect 204902 220895 204958 220904
rect 203616 182912 203668 182918
rect 203616 182854 203668 182860
rect 202236 143676 202288 143682
rect 202236 143618 202288 143624
rect 202248 59362 202276 143618
rect 202420 132592 202472 132598
rect 202420 132534 202472 132540
rect 202432 108322 202460 132534
rect 203616 121508 203668 121514
rect 203616 121450 203668 121456
rect 203524 114640 203576 114646
rect 203524 114582 203576 114588
rect 202512 112464 202564 112470
rect 202512 112406 202564 112412
rect 202420 108316 202472 108322
rect 202420 108258 202472 108264
rect 202328 107772 202380 107778
rect 202328 107714 202380 107720
rect 202340 81326 202368 107714
rect 202524 93226 202552 112406
rect 202512 93220 202564 93226
rect 202512 93162 202564 93168
rect 202328 81320 202380 81326
rect 202328 81262 202380 81268
rect 203536 67590 203564 114582
rect 203628 105602 203656 121450
rect 203616 105596 203668 105602
rect 203616 105538 203668 105544
rect 204916 97889 204944 220895
rect 205008 200802 205036 235282
rect 205100 235278 205128 236671
rect 205088 235272 205140 235278
rect 205088 235214 205140 235220
rect 205086 228440 205142 228449
rect 205086 228375 205142 228384
rect 205100 214674 205128 228375
rect 205376 222057 205404 240244
rect 205928 229094 205956 240244
rect 205928 229066 206232 229094
rect 205362 222048 205418 222057
rect 205362 221983 205418 221992
rect 206204 216186 206232 229066
rect 206284 225208 206336 225214
rect 206284 225150 206336 225156
rect 206296 217326 206324 225150
rect 206284 217320 206336 217326
rect 206284 217262 206336 217268
rect 206204 216158 206416 216186
rect 206282 216064 206338 216073
rect 206282 215999 206338 216008
rect 205088 214668 205140 214674
rect 205088 214610 205140 214616
rect 204996 200796 205048 200802
rect 204996 200738 205048 200744
rect 206296 188465 206324 215999
rect 206388 211041 206416 216158
rect 206480 215286 206508 240244
rect 206848 226302 206876 240244
rect 206836 226296 206888 226302
rect 206836 226238 206888 226244
rect 206848 225214 206876 226238
rect 206836 225208 206888 225214
rect 206836 225150 206888 225156
rect 206468 215280 206520 215286
rect 206468 215222 206520 215228
rect 206480 211993 206508 215222
rect 206466 211984 206522 211993
rect 206466 211919 206522 211928
rect 206374 211032 206430 211041
rect 206374 210967 206430 210976
rect 206388 191214 206416 210967
rect 207400 205601 207428 240244
rect 207386 205592 207442 205601
rect 207386 205527 207442 205536
rect 207952 200114 207980 240244
rect 208320 239465 208348 240244
rect 208306 239456 208362 239465
rect 208306 239391 208362 239400
rect 208320 238649 208348 239391
rect 208306 238640 208362 238649
rect 208306 238575 208362 238584
rect 208872 234433 208900 240244
rect 208858 234424 208914 234433
rect 208858 234359 208914 234368
rect 209136 233300 209188 233306
rect 209136 233242 209188 233248
rect 209042 224224 209098 224233
rect 209042 224159 209098 224168
rect 209056 206990 209084 224159
rect 209148 219337 209176 233242
rect 209240 231441 209268 240244
rect 209226 231432 209282 231441
rect 209226 231367 209282 231376
rect 209792 220969 209820 240244
rect 210344 235657 210372 240244
rect 210330 235648 210386 235657
rect 210330 235583 210386 235592
rect 210712 224233 210740 240244
rect 210698 224224 210754 224233
rect 210698 224159 210754 224168
rect 209778 220960 209834 220969
rect 209778 220895 209834 220904
rect 209134 219328 209190 219337
rect 209134 219263 209190 219272
rect 209792 213897 209820 220895
rect 209778 213888 209834 213897
rect 209778 213823 209834 213832
rect 210422 213208 210478 213217
rect 210422 213143 210478 213152
rect 209134 211848 209190 211857
rect 209134 211783 209190 211792
rect 209044 206984 209096 206990
rect 209044 206926 209096 206932
rect 207676 200086 207980 200114
rect 207676 198626 207704 200086
rect 207664 198620 207716 198626
rect 207664 198562 207716 198568
rect 207676 192506 207704 198562
rect 207664 192500 207716 192506
rect 207664 192442 207716 192448
rect 206376 191208 206428 191214
rect 206376 191150 206428 191156
rect 206282 188456 206338 188465
rect 206282 188391 206338 188400
rect 207664 184952 207716 184958
rect 207664 184894 207716 184900
rect 207020 176860 207072 176866
rect 207020 176802 207072 176808
rect 207032 175982 207060 176802
rect 207020 175976 207072 175982
rect 207020 175918 207072 175924
rect 207676 167113 207704 184894
rect 209148 181558 209176 211783
rect 210436 194546 210464 213143
rect 211264 209681 211292 240244
rect 211250 209672 211306 209681
rect 211250 209607 211306 209616
rect 211264 208457 211292 209607
rect 211250 208448 211306 208457
rect 211250 208383 211306 208392
rect 211816 206922 211844 240244
rect 212184 225049 212212 240244
rect 212170 225040 212226 225049
rect 212170 224975 212226 224984
rect 212184 222193 212212 224975
rect 212170 222184 212226 222193
rect 212170 222119 212226 222128
rect 211894 208448 211950 208457
rect 211894 208383 211950 208392
rect 211804 206916 211856 206922
rect 211804 206858 211856 206864
rect 211908 199442 211936 208383
rect 212448 206916 212500 206922
rect 212448 206858 212500 206864
rect 212460 206378 212488 206858
rect 212448 206372 212500 206378
rect 212448 206314 212500 206320
rect 212736 202473 212764 240244
rect 213104 237425 213132 240244
rect 213656 238754 213684 240244
rect 213656 238726 213868 238754
rect 214208 238746 214236 240244
rect 213656 238649 213684 238726
rect 213642 238640 213698 238649
rect 213642 238575 213698 238584
rect 213090 237416 213146 237425
rect 213090 237351 213146 237360
rect 213734 234696 213790 234705
rect 213734 234631 213790 234640
rect 213000 213988 213052 213994
rect 213000 213930 213052 213936
rect 213012 211138 213040 213930
rect 213000 211132 213052 211138
rect 213000 211074 213052 211080
rect 213748 209098 213776 234631
rect 213736 209092 213788 209098
rect 213736 209034 213788 209040
rect 213748 208418 213776 209034
rect 213736 208412 213788 208418
rect 213736 208354 213788 208360
rect 212722 202464 212778 202473
rect 212722 202399 212778 202408
rect 211896 199436 211948 199442
rect 211896 199378 211948 199384
rect 213840 196654 213868 238726
rect 214196 238740 214248 238746
rect 214196 238682 214248 238688
rect 214208 237522 214236 238682
rect 214576 238377 214604 240244
rect 215128 240145 215156 240244
rect 215114 240136 215170 240145
rect 215114 240071 215170 240080
rect 215128 238754 215156 240071
rect 215128 238726 215248 238754
rect 214562 238368 214618 238377
rect 214562 238303 214618 238312
rect 214196 237516 214248 237522
rect 214196 237458 214248 237464
rect 214656 237516 214708 237522
rect 214656 237458 214708 237464
rect 214564 237448 214616 237454
rect 214564 237390 214616 237396
rect 212080 196648 212132 196654
rect 212080 196590 212132 196596
rect 213828 196648 213880 196654
rect 213828 196590 213880 196596
rect 210424 194540 210476 194546
rect 210424 194482 210476 194488
rect 212092 193934 212120 196590
rect 214576 195906 214604 237390
rect 214668 213246 214696 237458
rect 214748 236700 214800 236706
rect 214748 236642 214800 236648
rect 214760 227050 214788 236642
rect 214748 227044 214800 227050
rect 214748 226986 214800 226992
rect 214748 225004 214800 225010
rect 214748 224946 214800 224952
rect 214656 213240 214708 213246
rect 214656 213182 214708 213188
rect 214760 210458 214788 224946
rect 214838 213888 214894 213897
rect 214838 213823 214894 213832
rect 214852 213314 214880 213823
rect 214840 213308 214892 213314
rect 214840 213250 214892 213256
rect 214852 210526 214880 213250
rect 214840 210520 214892 210526
rect 214840 210462 214892 210468
rect 214748 210452 214800 210458
rect 214748 210394 214800 210400
rect 214564 195900 214616 195906
rect 214564 195842 214616 195848
rect 212080 193928 212132 193934
rect 212080 193870 212132 193876
rect 214564 188352 214616 188358
rect 214564 188294 214616 188300
rect 209136 181552 209188 181558
rect 209136 181494 209188 181500
rect 209044 180872 209096 180878
rect 209044 180814 209096 180820
rect 207754 175400 207810 175409
rect 207754 175335 207810 175344
rect 207662 167104 207718 167113
rect 207662 167039 207718 167048
rect 207768 165753 207796 175335
rect 207754 165744 207810 165753
rect 207754 165679 207810 165688
rect 206284 151836 206336 151842
rect 206284 151778 206336 151784
rect 204996 133952 205048 133958
rect 204996 133894 205048 133900
rect 204902 97880 204958 97889
rect 204902 97815 204958 97824
rect 205008 84153 205036 133894
rect 205088 131164 205140 131170
rect 205088 131106 205140 131112
rect 205100 115161 205128 131106
rect 206296 124914 206324 151778
rect 206376 150544 206428 150550
rect 206376 150486 206428 150492
rect 206388 129062 206416 150486
rect 209056 150346 209084 180814
rect 214576 180198 214604 188294
rect 214564 180192 214616 180198
rect 214564 180134 214616 180140
rect 213920 176656 213972 176662
rect 213920 176598 213972 176604
rect 213932 175681 213960 176598
rect 215220 175982 215248 238726
rect 215680 229094 215708 240244
rect 216048 237454 216076 240244
rect 216036 237448 216088 237454
rect 216036 237390 216088 237396
rect 216048 237289 216076 237390
rect 216034 237280 216090 237289
rect 216034 237215 216090 237224
rect 216600 234433 216628 240244
rect 216586 234424 216642 234433
rect 216586 234359 216642 234368
rect 217152 231538 217180 240244
rect 217322 231840 217378 231849
rect 217322 231775 217378 231784
rect 217140 231532 217192 231538
rect 217140 231474 217192 231480
rect 217336 231130 217364 231775
rect 217324 231124 217376 231130
rect 217324 231066 217376 231072
rect 215680 229066 215984 229094
rect 215956 224942 215984 229066
rect 215944 224936 215996 224942
rect 215944 224878 215996 224884
rect 215956 188601 215984 224878
rect 217046 212392 217102 212401
rect 217046 212327 217102 212336
rect 217060 211177 217088 212327
rect 217046 211168 217102 211177
rect 217046 211103 217102 211112
rect 217230 189952 217286 189961
rect 217230 189887 217286 189896
rect 215942 188592 215998 188601
rect 215942 188527 215998 188536
rect 214104 175976 214156 175982
rect 214104 175918 214156 175924
rect 215208 175976 215260 175982
rect 215208 175918 215260 175924
rect 213918 175672 213974 175681
rect 213918 175607 213974 175616
rect 213920 175228 213972 175234
rect 213920 175170 213972 175176
rect 213932 175001 213960 175170
rect 214012 175160 214064 175166
rect 214012 175102 214064 175108
rect 213918 174992 213974 175001
rect 213918 174927 213974 174936
rect 214024 174321 214052 175102
rect 214010 174312 214066 174321
rect 214010 174247 214066 174256
rect 213920 173868 213972 173874
rect 213920 173810 213972 173816
rect 213932 173641 213960 173810
rect 214012 173800 214064 173806
rect 214012 173742 214064 173748
rect 213918 173632 213974 173641
rect 213918 173567 213974 173576
rect 214024 172961 214052 173742
rect 214010 172952 214066 172961
rect 214010 172887 214066 172896
rect 213920 172508 213972 172514
rect 213920 172450 213972 172456
rect 213932 172281 213960 172450
rect 213918 172272 213974 172281
rect 213918 172207 213974 172216
rect 214116 171601 214144 175918
rect 214562 175264 214618 175273
rect 214562 175199 214618 175208
rect 214576 173942 214604 175199
rect 214564 173936 214616 173942
rect 214564 173878 214616 173884
rect 214102 171592 214158 171601
rect 214102 171527 214158 171536
rect 214012 171080 214064 171086
rect 213918 171048 213974 171057
rect 214012 171022 214064 171028
rect 213918 170983 213920 170992
rect 213972 170983 213974 170992
rect 213920 170954 213972 170960
rect 214024 170377 214052 171022
rect 214010 170368 214066 170377
rect 214010 170303 214066 170312
rect 214012 169720 214064 169726
rect 213918 169688 213974 169697
rect 214012 169662 214064 169668
rect 213918 169623 213920 169632
rect 213972 169623 213974 169632
rect 213920 169594 213972 169600
rect 214024 169017 214052 169662
rect 214010 169008 214066 169017
rect 214010 168943 214066 168952
rect 213920 168360 213972 168366
rect 213918 168328 213920 168337
rect 213972 168328 213974 168337
rect 213918 168263 213974 168272
rect 214564 167680 214616 167686
rect 214564 167622 214616 167628
rect 213920 167000 213972 167006
rect 213918 166968 213920 166977
rect 213972 166968 213974 166977
rect 213918 166903 213974 166912
rect 214012 166932 214064 166938
rect 214012 166874 214064 166880
rect 214024 166433 214052 166874
rect 214010 166424 214066 166433
rect 214010 166359 214066 166368
rect 214012 165572 214064 165578
rect 214012 165514 214064 165520
rect 213920 165504 213972 165510
rect 213920 165446 213972 165452
rect 213932 165073 213960 165446
rect 213918 165064 213974 165073
rect 213918 164999 213974 165008
rect 214024 164393 214052 165514
rect 214010 164384 214066 164393
rect 214010 164319 214066 164328
rect 213920 164212 213972 164218
rect 213920 164154 213972 164160
rect 213932 163713 213960 164154
rect 214012 164144 214064 164150
rect 214012 164086 214064 164092
rect 213918 163704 213974 163713
rect 213918 163639 213974 163648
rect 214024 163033 214052 164086
rect 214010 163024 214066 163033
rect 214010 162959 214066 162968
rect 214012 162852 214064 162858
rect 214012 162794 214064 162800
rect 213920 162784 213972 162790
rect 213920 162726 213972 162732
rect 213932 162353 213960 162726
rect 213918 162344 213974 162353
rect 213918 162279 213974 162288
rect 214024 161809 214052 162794
rect 214010 161800 214066 161809
rect 214010 161735 214066 161744
rect 214012 161424 214064 161430
rect 214012 161366 214064 161372
rect 213920 161356 213972 161362
rect 213920 161298 213972 161304
rect 213932 161129 213960 161298
rect 213918 161120 213974 161129
rect 213918 161055 213974 161064
rect 214024 160449 214052 161366
rect 214010 160440 214066 160449
rect 214010 160375 214066 160384
rect 213920 160064 213972 160070
rect 213920 160006 213972 160012
rect 213932 159769 213960 160006
rect 214012 159996 214064 160002
rect 214012 159938 214064 159944
rect 213918 159760 213974 159769
rect 213918 159695 213974 159704
rect 214024 159089 214052 159938
rect 214010 159080 214066 159089
rect 214010 159015 214066 159024
rect 214012 158704 214064 158710
rect 214012 158646 214064 158652
rect 213920 158636 213972 158642
rect 213920 158578 213972 158584
rect 213932 158409 213960 158578
rect 213918 158400 213974 158409
rect 213918 158335 213974 158344
rect 214024 157729 214052 158646
rect 214010 157720 214066 157729
rect 214010 157655 214066 157664
rect 213920 157344 213972 157350
rect 213920 157286 213972 157292
rect 213932 157185 213960 157286
rect 214012 157276 214064 157282
rect 214012 157218 214064 157224
rect 213918 157176 213974 157185
rect 213918 157111 213974 157120
rect 214024 156505 214052 157218
rect 214010 156496 214066 156505
rect 214010 156431 214066 156440
rect 213920 155916 213972 155922
rect 213920 155858 213972 155864
rect 213932 155825 213960 155858
rect 214012 155848 214064 155854
rect 213918 155816 213974 155825
rect 214012 155790 214064 155796
rect 213918 155751 213974 155760
rect 214024 155145 214052 155790
rect 214010 155136 214066 155145
rect 214010 155071 214066 155080
rect 214010 154456 214066 154465
rect 214010 154391 214066 154400
rect 213918 153776 213974 153785
rect 213918 153711 213974 153720
rect 213932 153338 213960 153711
rect 213920 153332 213972 153338
rect 213920 153274 213972 153280
rect 214024 153270 214052 154391
rect 214012 153264 214064 153270
rect 214012 153206 214064 153212
rect 213182 153096 213238 153105
rect 213182 153031 213238 153040
rect 209044 150340 209096 150346
rect 209044 150282 209096 150288
rect 207754 145616 207810 145625
rect 207754 145551 207810 145560
rect 207664 129872 207716 129878
rect 207664 129814 207716 129820
rect 206376 129056 206428 129062
rect 206376 128998 206428 129004
rect 206376 125656 206428 125662
rect 206376 125598 206428 125604
rect 206284 124908 206336 124914
rect 206284 124850 206336 124856
rect 205086 115152 205142 115161
rect 205086 115087 205142 115096
rect 205180 104984 205232 104990
rect 205180 104926 205232 104932
rect 205088 90432 205140 90438
rect 205088 90374 205140 90380
rect 204994 84144 205050 84153
rect 204994 84079 205050 84088
rect 204904 80708 204956 80714
rect 204904 80650 204956 80656
rect 203524 67584 203576 67590
rect 203524 67526 203576 67532
rect 202236 59356 202288 59362
rect 202236 59298 202288 59304
rect 204916 10402 204944 80650
rect 205100 43450 205128 90374
rect 205192 84969 205220 104926
rect 206284 96688 206336 96694
rect 206284 96630 206336 96636
rect 206296 90370 206324 96630
rect 206284 90364 206336 90370
rect 206284 90306 206336 90312
rect 206284 89072 206336 89078
rect 206284 89014 206336 89020
rect 205178 84960 205234 84969
rect 205178 84895 205234 84904
rect 205088 43444 205140 43450
rect 205088 43386 205140 43392
rect 206296 13122 206324 89014
rect 206388 63510 206416 125598
rect 206468 117428 206520 117434
rect 206468 117370 206520 117376
rect 206376 63504 206428 63510
rect 206376 63446 206428 63452
rect 206480 56574 206508 117370
rect 207676 78577 207704 129814
rect 207768 93129 207796 145551
rect 209228 142248 209280 142254
rect 209228 142190 209280 142196
rect 209044 141432 209096 141438
rect 209044 141374 209096 141380
rect 207754 93120 207810 93129
rect 207754 93055 207810 93064
rect 207662 78568 207718 78577
rect 207662 78503 207718 78512
rect 206468 56568 206520 56574
rect 206468 56510 206520 56516
rect 209056 14550 209084 141374
rect 209136 135924 209188 135930
rect 209136 135866 209188 135872
rect 209148 96014 209176 135866
rect 209240 131782 209268 142190
rect 210608 139528 210660 139534
rect 210608 139470 210660 139476
rect 209228 131776 209280 131782
rect 209228 131718 209280 131724
rect 209320 131232 209372 131238
rect 209320 131174 209372 131180
rect 209228 106412 209280 106418
rect 209228 106354 209280 106360
rect 209136 96008 209188 96014
rect 209136 95950 209188 95956
rect 209134 91760 209190 91769
rect 209134 91695 209190 91704
rect 209044 14544 209096 14550
rect 209044 14486 209096 14492
rect 206284 13116 206336 13122
rect 206284 13058 206336 13064
rect 209148 11830 209176 91695
rect 209240 89729 209268 106354
rect 209332 91633 209360 131174
rect 210424 128444 210476 128450
rect 210424 128386 210476 128392
rect 209318 91624 209374 91633
rect 209318 91559 209374 91568
rect 209226 89720 209282 89729
rect 209226 89655 209282 89664
rect 210436 57934 210464 128386
rect 210516 111852 210568 111858
rect 210516 111794 210568 111800
rect 210528 70378 210556 111794
rect 210620 106865 210648 139470
rect 211804 139460 211856 139466
rect 211804 139402 211856 139408
rect 211816 127634 211844 139402
rect 211804 127628 211856 127634
rect 211804 127570 211856 127576
rect 211804 118788 211856 118794
rect 211804 118730 211856 118736
rect 210606 106856 210662 106865
rect 210606 106791 210662 106800
rect 211816 93809 211844 118730
rect 211988 113348 212040 113354
rect 211988 113290 212040 113296
rect 211896 99476 211948 99482
rect 211896 99418 211948 99424
rect 211802 93800 211858 93809
rect 211802 93735 211858 93744
rect 211804 83496 211856 83502
rect 211804 83438 211856 83444
rect 210516 70372 210568 70378
rect 210516 70314 210568 70320
rect 210424 57928 210476 57934
rect 210424 57870 210476 57876
rect 209136 11824 209188 11830
rect 209136 11766 209188 11772
rect 204904 10396 204956 10402
rect 204904 10338 204956 10344
rect 211816 6225 211844 83438
rect 211908 64870 211936 99418
rect 212000 91089 212028 113290
rect 213196 102814 213224 153031
rect 213918 152552 213974 152561
rect 213918 152487 213974 152496
rect 213932 151842 213960 152487
rect 213920 151836 213972 151842
rect 213920 151778 213972 151784
rect 214102 151192 214158 151201
rect 214102 151127 214158 151136
rect 213920 150544 213972 150550
rect 213918 150512 213920 150521
rect 213972 150512 213974 150521
rect 214116 150482 214144 151127
rect 213918 150447 213974 150456
rect 214104 150476 214156 150482
rect 214104 150418 214156 150424
rect 214012 150408 214064 150414
rect 214012 150350 214064 150356
rect 213920 150340 213972 150346
rect 213920 150282 213972 150288
rect 213932 149841 213960 150282
rect 213918 149832 213974 149841
rect 213918 149767 213974 149776
rect 214024 149161 214052 150350
rect 214010 149152 214066 149161
rect 214010 149087 214066 149096
rect 214576 148481 214604 167622
rect 214654 151872 214710 151881
rect 214654 151807 214710 151816
rect 214668 151065 214696 151807
rect 214654 151056 214710 151065
rect 214654 150991 214710 151000
rect 214562 148472 214618 148481
rect 214562 148407 214618 148416
rect 213918 147928 213974 147937
rect 213918 147863 213974 147872
rect 213932 147694 213960 147863
rect 213920 147688 213972 147694
rect 213920 147630 213972 147636
rect 213918 147248 213974 147257
rect 213918 147183 213974 147192
rect 213932 146334 213960 147183
rect 216126 146568 216182 146577
rect 216126 146503 216182 146512
rect 213920 146328 213972 146334
rect 213920 146270 213972 146276
rect 214010 145888 214066 145897
rect 214010 145823 214066 145832
rect 213918 145208 213974 145217
rect 213918 145143 213974 145152
rect 213932 144974 213960 145143
rect 214024 145042 214052 145823
rect 214012 145036 214064 145042
rect 214012 144978 214064 144984
rect 213920 144968 213972 144974
rect 213920 144910 213972 144916
rect 214010 144528 214066 144537
rect 214010 144463 214066 144472
rect 213918 143848 213974 143857
rect 213918 143783 213974 143792
rect 213932 143614 213960 143783
rect 214024 143682 214052 144463
rect 214012 143676 214064 143682
rect 214012 143618 214064 143624
rect 213920 143608 213972 143614
rect 213920 143550 213972 143556
rect 214010 143304 214066 143313
rect 214010 143239 214066 143248
rect 213918 142624 213974 142633
rect 213918 142559 213974 142568
rect 213932 142254 213960 142559
rect 213920 142248 213972 142254
rect 213920 142190 213972 142196
rect 214024 142186 214052 143239
rect 214012 142180 214064 142186
rect 214012 142122 214064 142128
rect 213918 141944 213974 141953
rect 213918 141879 213974 141888
rect 213932 140826 213960 141879
rect 214010 141264 214066 141273
rect 214010 141199 214066 141208
rect 213920 140820 213972 140826
rect 213920 140762 213972 140768
rect 213918 140584 213974 140593
rect 213918 140519 213974 140528
rect 213932 139466 213960 140519
rect 213920 139460 213972 139466
rect 213920 139402 213972 139408
rect 213918 139224 213974 139233
rect 213918 139159 213974 139168
rect 213932 138038 213960 139159
rect 213920 138032 213972 138038
rect 213920 137974 213972 137980
rect 213918 137320 213974 137329
rect 214024 137290 214052 141199
rect 214102 139904 214158 139913
rect 214102 139839 214158 139848
rect 214116 139534 214144 139839
rect 214104 139528 214156 139534
rect 214104 139470 214156 139476
rect 214654 138680 214710 138689
rect 214654 138615 214710 138624
rect 213918 137255 213974 137264
rect 214012 137284 214064 137290
rect 213932 136678 213960 137255
rect 214012 137226 214064 137232
rect 213920 136672 213972 136678
rect 213920 136614 213972 136620
rect 214010 135960 214066 135969
rect 214010 135895 214066 135904
rect 213920 135312 213972 135318
rect 213918 135280 213920 135289
rect 213972 135280 213974 135289
rect 213918 135215 213974 135224
rect 214024 134570 214052 135895
rect 214562 134600 214618 134609
rect 214012 134564 214064 134570
rect 214562 134535 214618 134544
rect 214012 134506 214064 134512
rect 213920 133952 213972 133958
rect 213918 133920 213920 133929
rect 213972 133920 213974 133929
rect 213918 133855 213974 133864
rect 214010 133376 214066 133385
rect 214010 133311 214066 133320
rect 213274 133104 213330 133113
rect 213274 133039 213330 133048
rect 213184 102808 213236 102814
rect 213184 102750 213236 102756
rect 213288 93838 213316 133039
rect 213918 132696 213974 132705
rect 213918 132631 213974 132640
rect 213932 132598 213960 132631
rect 213920 132592 213972 132598
rect 213920 132534 213972 132540
rect 214024 132530 214052 133311
rect 214012 132524 214064 132530
rect 214012 132466 214064 132472
rect 214010 132016 214066 132025
rect 214010 131951 214066 131960
rect 213918 131336 213974 131345
rect 213918 131271 213974 131280
rect 213932 131238 213960 131271
rect 213920 131232 213972 131238
rect 213920 131174 213972 131180
rect 214024 131170 214052 131951
rect 214012 131164 214064 131170
rect 214012 131106 214064 131112
rect 214010 130656 214066 130665
rect 214010 130591 214066 130600
rect 213918 129976 213974 129985
rect 213918 129911 213974 129920
rect 213932 129878 213960 129911
rect 213920 129872 213972 129878
rect 213920 129814 213972 129820
rect 214024 129810 214052 130591
rect 214012 129804 214064 129810
rect 214012 129746 214064 129752
rect 213918 129296 213974 129305
rect 213918 129231 213974 129240
rect 213932 128382 213960 129231
rect 214010 128752 214066 128761
rect 214010 128687 214066 128696
rect 214024 128450 214052 128687
rect 214012 128444 214064 128450
rect 214012 128386 214064 128392
rect 213920 128376 213972 128382
rect 213920 128318 213972 128324
rect 214010 128072 214066 128081
rect 214010 128007 214066 128016
rect 213918 127392 213974 127401
rect 213918 127327 213974 127336
rect 213932 127022 213960 127327
rect 213920 127016 213972 127022
rect 213920 126958 213972 126964
rect 214024 126313 214052 128007
rect 214010 126304 214066 126313
rect 214576 126274 214604 134535
rect 214010 126239 214066 126248
rect 214564 126268 214616 126274
rect 214564 126210 214616 126216
rect 213918 126032 213974 126041
rect 213918 125967 213974 125976
rect 213932 125662 213960 125967
rect 213920 125656 213972 125662
rect 213920 125598 213972 125604
rect 214562 125352 214618 125361
rect 214562 125287 214618 125296
rect 213918 124672 213974 124681
rect 213918 124607 213974 124616
rect 213932 124234 213960 124607
rect 213920 124228 213972 124234
rect 213920 124170 213972 124176
rect 214010 124128 214066 124137
rect 214010 124063 214066 124072
rect 213918 123448 213974 123457
rect 213918 123383 213974 123392
rect 213932 122874 213960 123383
rect 214024 122942 214052 124063
rect 214012 122936 214064 122942
rect 214012 122878 214064 122884
rect 213920 122868 213972 122874
rect 213920 122810 213972 122816
rect 213918 122768 213974 122777
rect 213918 122703 213974 122712
rect 213366 122088 213422 122097
rect 213366 122023 213422 122032
rect 213380 94518 213408 122023
rect 213932 121514 213960 122703
rect 214576 122126 214604 125287
rect 214564 122120 214616 122126
rect 214564 122062 214616 122068
rect 213920 121508 213972 121514
rect 213920 121450 213972 121456
rect 214010 121408 214066 121417
rect 214010 121343 214066 121352
rect 213918 120728 213974 120737
rect 213918 120663 213974 120672
rect 213932 120222 213960 120663
rect 213920 120216 213972 120222
rect 213920 120158 213972 120164
rect 214024 120154 214052 121343
rect 214012 120148 214064 120154
rect 214012 120090 214064 120096
rect 214010 120048 214066 120057
rect 214010 119983 214066 119992
rect 213918 119504 213974 119513
rect 213918 119439 213974 119448
rect 213932 118726 213960 119439
rect 214024 118794 214052 119983
rect 214012 118788 214064 118794
rect 214012 118730 214064 118736
rect 213920 118720 213972 118726
rect 213920 118662 213972 118668
rect 214010 118144 214066 118153
rect 214010 118079 214066 118088
rect 213918 117464 213974 117473
rect 213918 117399 213920 117408
rect 213972 117399 213974 117408
rect 213920 117370 213972 117376
rect 214024 117366 214052 118079
rect 214012 117360 214064 117366
rect 214012 117302 214064 117308
rect 214010 116784 214066 116793
rect 214010 116719 214066 116728
rect 213918 116104 213974 116113
rect 213918 116039 213920 116048
rect 213972 116039 213974 116048
rect 213920 116010 213972 116016
rect 214024 116006 214052 116719
rect 214562 116512 214618 116521
rect 214562 116447 214618 116456
rect 214012 116000 214064 116006
rect 214012 115942 214064 115948
rect 214010 115424 214066 115433
rect 214010 115359 214066 115368
rect 213918 114880 213974 114889
rect 213918 114815 213974 114824
rect 213932 114578 213960 114815
rect 214024 114646 214052 115359
rect 214012 114640 214064 114646
rect 214012 114582 214064 114588
rect 213920 114572 213972 114578
rect 213920 114514 213972 114520
rect 213918 114200 213974 114209
rect 213918 114135 213974 114144
rect 213932 113218 213960 114135
rect 214286 113520 214342 113529
rect 214286 113455 214342 113464
rect 214300 113354 214328 113455
rect 214288 113348 214340 113354
rect 214288 113290 214340 113296
rect 213920 113212 213972 113218
rect 213920 113154 213972 113160
rect 213918 112840 213974 112849
rect 213918 112775 213974 112784
rect 213932 111858 213960 112775
rect 213920 111852 213972 111858
rect 213920 111794 213972 111800
rect 214010 111480 214066 111489
rect 214010 111415 214066 111424
rect 213918 110800 213974 110809
rect 213918 110735 213974 110744
rect 213932 110566 213960 110735
rect 213920 110560 213972 110566
rect 213920 110502 213972 110508
rect 214024 110498 214052 111415
rect 214012 110492 214064 110498
rect 214012 110434 214064 110440
rect 214010 110256 214066 110265
rect 214010 110191 214066 110200
rect 213918 109576 213974 109585
rect 213918 109511 213974 109520
rect 213932 109138 213960 109511
rect 213920 109132 213972 109138
rect 213920 109074 213972 109080
rect 214024 109070 214052 110191
rect 214012 109064 214064 109070
rect 214012 109006 214064 109012
rect 214010 108896 214066 108905
rect 214010 108831 214066 108840
rect 213918 108216 213974 108225
rect 213918 108151 213974 108160
rect 213932 107778 213960 108151
rect 213920 107772 213972 107778
rect 213920 107714 213972 107720
rect 214024 107710 214052 108831
rect 214012 107704 214064 107710
rect 214012 107646 214064 107652
rect 214010 107536 214066 107545
rect 214010 107471 214066 107480
rect 213918 106856 213974 106865
rect 213918 106791 213974 106800
rect 213932 106350 213960 106791
rect 214024 106418 214052 107471
rect 214012 106412 214064 106418
rect 214012 106354 214064 106360
rect 213920 106344 213972 106350
rect 213920 106286 213972 106292
rect 214010 106176 214066 106185
rect 214010 106111 214066 106120
rect 213920 104984 213972 104990
rect 213918 104952 213920 104961
rect 213972 104952 213974 104961
rect 214024 104922 214052 106111
rect 213918 104887 213974 104896
rect 214012 104916 214064 104922
rect 214012 104858 214064 104864
rect 214010 104272 214066 104281
rect 214010 104207 214066 104216
rect 214024 103630 214052 104207
rect 214012 103624 214064 103630
rect 213918 103592 213974 103601
rect 214012 103566 214064 103572
rect 213918 103527 213920 103536
rect 213972 103527 213974 103536
rect 213920 103498 213972 103504
rect 213458 102232 213514 102241
rect 213458 102167 213514 102176
rect 213368 94512 213420 94518
rect 213368 94454 213420 94460
rect 213276 93832 213328 93838
rect 213276 93774 213328 93780
rect 211986 91080 212042 91089
rect 211986 91015 212042 91024
rect 213184 87712 213236 87718
rect 213184 87654 213236 87660
rect 211896 64864 211948 64870
rect 211896 64806 211948 64812
rect 213196 28286 213224 87654
rect 213274 87544 213330 87553
rect 213274 87479 213330 87488
rect 213288 71233 213316 87479
rect 213472 82793 213500 102167
rect 214194 101552 214250 101561
rect 214194 101487 214250 101496
rect 213918 101008 213974 101017
rect 213918 100943 213974 100952
rect 213932 100774 213960 100943
rect 213920 100768 213972 100774
rect 213920 100710 213972 100716
rect 214010 100328 214066 100337
rect 214010 100263 214066 100272
rect 213918 99648 213974 99657
rect 213918 99583 213974 99592
rect 213932 99414 213960 99583
rect 214024 99482 214052 100263
rect 214012 99476 214064 99482
rect 214012 99418 214064 99424
rect 213920 99408 213972 99414
rect 213920 99350 213972 99356
rect 214102 98968 214158 98977
rect 214102 98903 214158 98912
rect 213918 98288 213974 98297
rect 213918 98223 213974 98232
rect 213932 98054 213960 98223
rect 213920 98048 213972 98054
rect 213920 97990 213972 97996
rect 213918 97608 213974 97617
rect 213918 97543 213974 97552
rect 213932 96694 213960 97543
rect 213920 96688 213972 96694
rect 213920 96630 213972 96636
rect 214010 96384 214066 96393
rect 214010 96319 214066 96328
rect 214024 88233 214052 96319
rect 214116 95946 214144 98903
rect 214104 95940 214156 95946
rect 214104 95882 214156 95888
rect 214208 95849 214236 101487
rect 214470 97880 214526 97889
rect 214470 97815 214526 97824
rect 214484 96694 214512 97815
rect 214472 96688 214524 96694
rect 214472 96630 214524 96636
rect 214194 95840 214250 95849
rect 214194 95775 214250 95784
rect 214010 88224 214066 88233
rect 214010 88159 214066 88168
rect 213458 82784 213514 82793
rect 213458 82719 213514 82728
rect 213274 71224 213330 71233
rect 213274 71159 213330 71168
rect 213184 28280 213236 28286
rect 213184 28222 213236 28228
rect 214576 13122 214604 116447
rect 214668 103514 214696 138615
rect 216034 138000 216090 138009
rect 216034 137935 216090 137944
rect 215942 136640 215998 136649
rect 215942 136575 215998 136584
rect 214746 126712 214802 126721
rect 214746 126647 214802 126656
rect 214760 112470 214788 126647
rect 215956 113801 215984 136575
rect 215942 113792 215998 113801
rect 215942 113727 215998 113736
rect 214748 112464 214800 112470
rect 214748 112406 214800 112412
rect 214668 103486 214880 103514
rect 214852 97306 214880 103486
rect 214840 97300 214892 97306
rect 214840 97242 214892 97248
rect 214746 96928 214802 96937
rect 214746 96863 214802 96872
rect 214656 91860 214708 91866
rect 214656 91802 214708 91808
rect 214564 13116 214616 13122
rect 214564 13058 214616 13064
rect 211802 6216 211858 6225
rect 211802 6151 211858 6160
rect 202144 3528 202196 3534
rect 202144 3470 202196 3476
rect 214668 3466 214696 91802
rect 214760 66230 214788 96863
rect 215942 93256 215998 93265
rect 215942 93191 215998 93200
rect 214748 66224 214800 66230
rect 214748 66166 214800 66172
rect 215956 33862 215984 93191
rect 216048 92313 216076 137935
rect 216140 93673 216168 146503
rect 216218 94480 216274 94489
rect 216218 94415 216274 94424
rect 216126 93664 216182 93673
rect 216126 93599 216182 93608
rect 216034 92304 216090 92313
rect 216034 92239 216090 92248
rect 216232 51785 216260 94415
rect 217244 93770 217272 189887
rect 217336 177449 217364 231066
rect 217520 212401 217548 240244
rect 217506 212392 217562 212401
rect 217506 212327 217562 212336
rect 218072 208321 218100 240244
rect 218152 240168 218204 240174
rect 218152 240110 218204 240116
rect 218164 238746 218192 240110
rect 218152 238740 218204 238746
rect 218152 238682 218204 238688
rect 218440 229094 218468 240244
rect 218992 233170 219020 240244
rect 219544 238649 219572 240244
rect 219912 238754 219940 240244
rect 219912 238726 220216 238754
rect 219912 238678 219940 238726
rect 219900 238672 219952 238678
rect 219530 238640 219586 238649
rect 219900 238614 219952 238620
rect 219530 238575 219586 238584
rect 218980 233164 219032 233170
rect 218980 233106 219032 233112
rect 219532 231872 219584 231878
rect 219532 231814 219584 231820
rect 218440 229066 218836 229094
rect 218808 216617 218836 229066
rect 219544 217977 219572 231814
rect 220084 227792 220136 227798
rect 220084 227734 220136 227740
rect 219530 217968 219586 217977
rect 219530 217903 219586 217912
rect 218794 216608 218850 216617
rect 218794 216543 218850 216552
rect 218058 208312 218114 208321
rect 218058 208247 218114 208256
rect 218072 207097 218100 208247
rect 218058 207088 218114 207097
rect 218058 207023 218114 207032
rect 218702 207088 218758 207097
rect 218702 207023 218758 207032
rect 218716 181665 218744 207023
rect 218808 204950 218836 216543
rect 218888 205012 218940 205018
rect 218888 204954 218940 204960
rect 218796 204944 218848 204950
rect 218796 204886 218848 204892
rect 218900 195294 218928 204954
rect 218888 195288 218940 195294
rect 218888 195230 218940 195236
rect 218702 181656 218758 181665
rect 218702 181591 218758 181600
rect 217322 177440 217378 177449
rect 217322 177375 217378 177384
rect 220096 176050 220124 227734
rect 220188 206310 220216 238726
rect 220360 233164 220412 233170
rect 220360 233106 220412 233112
rect 220372 231878 220400 233106
rect 220360 231872 220412 231878
rect 220360 231814 220412 231820
rect 220464 229090 220492 240244
rect 221016 233306 221044 240244
rect 221094 240136 221150 240145
rect 221094 240071 221150 240080
rect 221108 238678 221136 240071
rect 221096 238672 221148 238678
rect 221096 238614 221148 238620
rect 221004 233300 221056 233306
rect 221004 233242 221056 233248
rect 221384 232665 221412 240244
rect 221936 232801 221964 240244
rect 222108 233300 222160 233306
rect 222108 233242 222160 233248
rect 221922 232792 221978 232801
rect 221922 232727 221978 232736
rect 221370 232656 221426 232665
rect 221370 232591 221426 232600
rect 221554 232520 221610 232529
rect 221554 232455 221610 232464
rect 221464 231532 221516 231538
rect 221464 231474 221516 231480
rect 220452 229084 220504 229090
rect 220452 229026 220504 229032
rect 220268 227860 220320 227866
rect 220268 227802 220320 227808
rect 220280 213761 220308 227802
rect 220464 227798 220492 229026
rect 220452 227792 220504 227798
rect 220452 227734 220504 227740
rect 220266 213752 220322 213761
rect 220266 213687 220322 213696
rect 220266 211168 220322 211177
rect 220266 211103 220322 211112
rect 220176 206304 220228 206310
rect 220176 206246 220228 206252
rect 220280 185638 220308 211103
rect 220728 189780 220780 189786
rect 220728 189722 220780 189728
rect 220740 187105 220768 189722
rect 221476 189174 221504 231474
rect 221568 197305 221596 232455
rect 222120 231169 222148 233242
rect 222106 231160 222162 231169
rect 222106 231095 222162 231104
rect 222304 213858 222332 240244
rect 222856 230382 222884 240244
rect 222844 230376 222896 230382
rect 222844 230318 222896 230324
rect 222292 213852 222344 213858
rect 222292 213794 222344 213800
rect 221554 197296 221610 197305
rect 221554 197231 221610 197240
rect 221464 189168 221516 189174
rect 221464 189110 221516 189116
rect 221476 187678 221504 189110
rect 221464 187672 221516 187678
rect 221464 187614 221516 187620
rect 222106 187640 222162 187649
rect 222106 187575 222162 187584
rect 220726 187096 220782 187105
rect 220726 187031 220782 187040
rect 222120 186386 222148 187575
rect 222108 186380 222160 186386
rect 222108 186322 222160 186328
rect 220268 185632 220320 185638
rect 220268 185574 220320 185580
rect 220266 179480 220322 179489
rect 220266 179415 220322 179424
rect 220280 176633 220308 179415
rect 222856 177410 222884 230318
rect 223408 219366 223436 240244
rect 223776 220726 223804 240244
rect 224328 237386 224356 240244
rect 224316 237380 224368 237386
rect 224316 237322 224368 237328
rect 224328 236706 224356 237322
rect 224316 236700 224368 236706
rect 224316 236642 224368 236648
rect 224880 224874 224908 240244
rect 224960 240168 225012 240174
rect 224958 240136 224960 240145
rect 225012 240136 225014 240145
rect 224958 240071 225014 240080
rect 225248 237153 225276 240244
rect 225800 238754 225828 240244
rect 225524 238726 225828 238754
rect 225234 237144 225290 237153
rect 225234 237079 225290 237088
rect 224316 224868 224368 224874
rect 224316 224810 224368 224816
rect 224868 224868 224920 224874
rect 224868 224810 224920 224816
rect 223764 220720 223816 220726
rect 223764 220662 223816 220668
rect 223776 219978 223804 220662
rect 223764 219972 223816 219978
rect 223764 219914 223816 219920
rect 224224 219972 224276 219978
rect 224224 219914 224276 219920
rect 223396 219360 223448 219366
rect 223396 219302 223448 219308
rect 223408 218142 223436 219302
rect 222936 218136 222988 218142
rect 222936 218078 222988 218084
rect 223396 218136 223448 218142
rect 223396 218078 223448 218084
rect 222844 177404 222896 177410
rect 222844 177346 222896 177352
rect 222948 176633 222976 218078
rect 223028 213852 223080 213858
rect 223028 213794 223080 213800
rect 223040 199510 223068 213794
rect 223028 199504 223080 199510
rect 223028 199446 223080 199452
rect 223028 196036 223080 196042
rect 223028 195978 223080 195984
rect 223040 189038 223068 195978
rect 223028 189032 223080 189038
rect 223028 188974 223080 188980
rect 224236 180794 224264 219914
rect 224328 188358 224356 224810
rect 225524 219434 225552 238726
rect 225696 236088 225748 236094
rect 225696 236030 225748 236036
rect 225604 234660 225656 234666
rect 225604 234602 225656 234608
rect 225616 226137 225644 234602
rect 225708 227497 225736 236030
rect 226168 234666 226196 240244
rect 226720 238513 226748 240244
rect 226706 238504 226762 238513
rect 226706 238439 226762 238448
rect 226156 234660 226208 234666
rect 226156 234602 226208 234608
rect 227272 228478 227300 240244
rect 227640 238678 227668 240244
rect 227812 240168 227864 240174
rect 227812 240110 227864 240116
rect 227628 238672 227680 238678
rect 227628 238614 227680 238620
rect 227260 228472 227312 228478
rect 227260 228414 227312 228420
rect 227272 227866 227300 228414
rect 227260 227860 227312 227866
rect 227260 227802 227312 227808
rect 225694 227488 225750 227497
rect 225694 227423 225750 227432
rect 225602 226128 225658 226137
rect 225602 226063 225658 226072
rect 226984 222896 227036 222902
rect 226984 222838 227036 222844
rect 224972 219406 225552 219434
rect 224408 218748 224460 218754
rect 224408 218690 224460 218696
rect 224420 200025 224448 218690
rect 224972 215257 225000 219406
rect 224958 215248 225014 215257
rect 224958 215183 225014 215192
rect 224972 214849 225000 215183
rect 224958 214840 225014 214849
rect 224958 214775 225014 214784
rect 225694 214840 225750 214849
rect 225694 214775 225750 214784
rect 225602 202328 225658 202337
rect 225602 202263 225658 202272
rect 224406 200016 224462 200025
rect 224406 199951 224462 199960
rect 224316 188352 224368 188358
rect 224316 188294 224368 188300
rect 225616 184385 225644 202263
rect 225708 200870 225736 214775
rect 226996 211857 227024 222838
rect 227824 212498 227852 240110
rect 228192 233209 228220 240244
rect 228744 239737 228772 240244
rect 228730 239728 228786 239737
rect 228730 239663 228786 239672
rect 229006 239728 229062 239737
rect 229006 239663 229062 239672
rect 228178 233200 228234 233209
rect 228178 233135 228234 233144
rect 229020 224262 229048 239663
rect 229112 238134 229140 240244
rect 229100 238128 229152 238134
rect 229100 238070 229152 238076
rect 229664 236094 229692 240244
rect 229742 240136 229798 240145
rect 229742 240071 229798 240080
rect 229652 236088 229704 236094
rect 229652 236030 229704 236036
rect 229008 224256 229060 224262
rect 229008 224198 229060 224204
rect 227812 212492 227864 212498
rect 227812 212434 227864 212440
rect 228364 212492 228416 212498
rect 228364 212434 228416 212440
rect 226982 211848 227038 211857
rect 226982 211783 227038 211792
rect 225878 205048 225934 205057
rect 225878 204983 225934 204992
rect 225696 200864 225748 200870
rect 225696 200806 225748 200812
rect 225892 194041 225920 204983
rect 226984 196648 227036 196654
rect 226984 196590 227036 196596
rect 226338 196072 226394 196081
rect 226338 196007 226394 196016
rect 226352 195974 226380 196007
rect 226340 195968 226392 195974
rect 226340 195910 226392 195916
rect 225694 194032 225750 194041
rect 225694 193967 225750 193976
rect 225878 194032 225934 194041
rect 225878 193967 225934 193976
rect 225602 184376 225658 184385
rect 225602 184311 225658 184320
rect 224236 180766 224356 180794
rect 224224 180124 224276 180130
rect 224224 180066 224276 180072
rect 224236 179314 224264 180066
rect 224328 179450 224356 180766
rect 225708 180169 225736 193967
rect 225694 180160 225750 180169
rect 225694 180095 225750 180104
rect 224316 179444 224368 179450
rect 224316 179386 224368 179392
rect 224224 179308 224276 179314
rect 224224 179250 224276 179256
rect 226996 177313 227024 196590
rect 228376 189825 228404 212434
rect 228454 196072 228510 196081
rect 228454 196007 228510 196016
rect 228362 189816 228418 189825
rect 228362 189751 228418 189760
rect 227718 177440 227774 177449
rect 227718 177375 227774 177384
rect 224958 177304 225014 177313
rect 224958 177239 225014 177248
rect 226982 177304 227038 177313
rect 226982 177239 227038 177248
rect 220266 176624 220322 176633
rect 220266 176559 220322 176568
rect 222934 176624 222990 176633
rect 222934 176559 222990 176568
rect 220084 176044 220136 176050
rect 220084 175986 220136 175992
rect 224972 175846 225000 177239
rect 227732 176225 227760 177375
rect 227718 176216 227774 176225
rect 227718 176151 227774 176160
rect 228468 176089 228496 196007
rect 229468 179444 229520 179450
rect 229468 179386 229520 179392
rect 229376 177336 229428 177342
rect 229376 177278 229428 177284
rect 228454 176080 228510 176089
rect 228454 176015 228510 176024
rect 229192 175976 229244 175982
rect 229192 175918 229244 175924
rect 224960 175840 225012 175846
rect 224960 175782 225012 175788
rect 229098 175128 229154 175137
rect 229098 175063 229154 175072
rect 229112 173777 229140 175063
rect 229098 173768 229154 173777
rect 229098 173703 229154 173712
rect 229100 173664 229152 173670
rect 229100 173606 229152 173612
rect 229112 146849 229140 173606
rect 229204 164393 229232 175918
rect 229284 175228 229336 175234
rect 229284 175170 229336 175176
rect 229296 175001 229324 175170
rect 229282 174992 229338 175001
rect 229282 174927 229338 174936
rect 229388 167657 229416 177278
rect 229480 173670 229508 179386
rect 229756 176769 229784 240071
rect 230216 219201 230244 240244
rect 230584 240145 230612 240244
rect 230570 240136 230626 240145
rect 230570 240071 230626 240080
rect 230480 238128 230532 238134
rect 230480 238070 230532 238076
rect 230492 233238 230520 238070
rect 230584 237425 230612 240071
rect 231136 238610 231164 240244
rect 231124 238604 231176 238610
rect 231124 238546 231176 238552
rect 230570 237416 230626 237425
rect 230570 237351 230626 237360
rect 230480 233232 230532 233238
rect 230480 233174 230532 233180
rect 231504 231305 231532 240244
rect 232056 238754 232084 240244
rect 232056 238726 232176 238754
rect 231766 237960 231822 237969
rect 231766 237895 231822 237904
rect 231674 237416 231730 237425
rect 231780 237386 231808 237895
rect 231674 237351 231730 237360
rect 231768 237380 231820 237386
rect 231490 231296 231546 231305
rect 231490 231231 231546 231240
rect 231688 229094 231716 237351
rect 231768 237322 231820 237328
rect 231768 233232 231820 233238
rect 231768 233174 231820 233180
rect 231780 231130 231808 233174
rect 231768 231124 231820 231130
rect 231768 231066 231820 231072
rect 231688 229066 231808 229094
rect 230202 219192 230258 219201
rect 230202 219127 230258 219136
rect 230480 215960 230532 215966
rect 230480 215902 230532 215908
rect 229928 179308 229980 179314
rect 229928 179250 229980 179256
rect 229742 176760 229798 176769
rect 229742 176695 229798 176704
rect 229940 175234 229968 179250
rect 229928 175228 229980 175234
rect 229928 175170 229980 175176
rect 229468 173664 229520 173670
rect 229468 173606 229520 173612
rect 229744 167680 229796 167686
rect 229374 167648 229430 167657
rect 229744 167622 229796 167628
rect 229374 167583 229430 167592
rect 229190 164384 229246 164393
rect 229190 164319 229246 164328
rect 229756 148209 229784 167622
rect 230492 166326 230520 215902
rect 231124 206372 231176 206378
rect 231124 206314 231176 206320
rect 230572 193860 230624 193866
rect 230572 193802 230624 193808
rect 230584 171134 230612 193802
rect 231136 176186 231164 206314
rect 231780 196081 231808 229066
rect 232148 204270 232176 238726
rect 232608 224777 232636 240244
rect 232594 224768 232650 224777
rect 232594 224703 232650 224712
rect 232136 204264 232188 204270
rect 232136 204206 232188 204212
rect 231952 203720 232004 203726
rect 231952 203662 232004 203668
rect 231766 196072 231822 196081
rect 231766 196007 231822 196016
rect 231216 185700 231268 185706
rect 231216 185642 231268 185648
rect 231228 177342 231256 185642
rect 231216 177336 231268 177342
rect 231216 177278 231268 177284
rect 231124 176180 231176 176186
rect 231124 176122 231176 176128
rect 231860 176044 231912 176050
rect 231860 175986 231912 175992
rect 231766 175944 231822 175953
rect 231766 175879 231822 175888
rect 231780 175273 231808 175879
rect 231766 175264 231822 175273
rect 230848 175228 230900 175234
rect 230848 175170 230900 175176
rect 231124 175228 231176 175234
rect 231766 175199 231822 175208
rect 231124 175170 231176 175176
rect 230860 171134 230888 175170
rect 231136 174729 231164 175170
rect 231122 174720 231178 174729
rect 231122 174655 231178 174664
rect 231584 173868 231636 173874
rect 231584 173810 231636 173816
rect 231596 172825 231624 173810
rect 231766 173224 231822 173233
rect 231766 173159 231822 173168
rect 231582 172816 231638 172825
rect 231582 172751 231638 172760
rect 231584 172508 231636 172514
rect 231584 172450 231636 172456
rect 231596 171465 231624 172450
rect 231780 171873 231808 173159
rect 231766 171864 231822 171873
rect 231766 171799 231822 171808
rect 231582 171456 231638 171465
rect 231582 171391 231638 171400
rect 230584 171106 230704 171134
rect 230480 166320 230532 166326
rect 230480 166262 230532 166268
rect 230110 162208 230166 162217
rect 230110 162143 230166 162152
rect 229742 148200 229798 148209
rect 229742 148135 229798 148144
rect 229098 146840 229154 146849
rect 229098 146775 229154 146784
rect 229928 138712 229980 138718
rect 229928 138654 229980 138660
rect 229742 138408 229798 138417
rect 229742 138343 229798 138352
rect 219164 96076 219216 96082
rect 219164 96018 219216 96024
rect 219256 96076 219308 96082
rect 219256 96018 219308 96024
rect 219176 95849 219204 96018
rect 219268 95985 219296 96018
rect 220084 96008 220136 96014
rect 219254 95976 219310 95985
rect 220084 95950 220136 95956
rect 226982 95976 227038 95985
rect 219254 95911 219310 95920
rect 219162 95840 219218 95849
rect 219162 95775 219218 95784
rect 217324 94512 217376 94518
rect 217324 94454 217376 94460
rect 217232 93764 217284 93770
rect 217232 93706 217284 93712
rect 216218 51776 216274 51785
rect 216218 51711 216274 51720
rect 215944 33856 215996 33862
rect 215944 33798 215996 33804
rect 217336 21486 217364 94454
rect 218704 90364 218756 90370
rect 218704 90306 218756 90312
rect 218716 47598 218744 90306
rect 218704 47592 218756 47598
rect 218704 47534 218756 47540
rect 217324 21480 217376 21486
rect 217324 21422 217376 21428
rect 220096 6225 220124 95950
rect 226982 95911 227038 95920
rect 224408 95260 224460 95266
rect 224408 95202 224460 95208
rect 224222 91896 224278 91905
rect 224222 91831 224278 91840
rect 223028 86352 223080 86358
rect 223028 86294 223080 86300
rect 220174 86184 220230 86193
rect 220174 86119 220230 86128
rect 220188 15910 220216 86119
rect 222844 83564 222896 83570
rect 222844 83506 222896 83512
rect 221462 50416 221518 50425
rect 221462 50351 221518 50360
rect 221476 25634 221504 50351
rect 221464 25628 221516 25634
rect 221464 25570 221516 25576
rect 222856 24138 222884 83506
rect 222936 47660 222988 47666
rect 222936 47602 222988 47608
rect 222844 24132 222896 24138
rect 222844 24074 222896 24080
rect 220176 15904 220228 15910
rect 220176 15846 220228 15852
rect 220082 6216 220138 6225
rect 220082 6151 220138 6160
rect 214656 3460 214708 3466
rect 214656 3402 214708 3408
rect 222948 2786 222976 47602
rect 223040 47598 223068 86294
rect 223028 47592 223080 47598
rect 223028 47534 223080 47540
rect 224236 18698 224264 91831
rect 224420 79529 224448 95202
rect 225604 84924 225656 84930
rect 225604 84866 225656 84872
rect 224406 79520 224462 79529
rect 224406 79455 224462 79464
rect 224316 79348 224368 79354
rect 224316 79290 224368 79296
rect 224224 18692 224276 18698
rect 224224 18634 224276 18640
rect 224328 6254 224356 79290
rect 225616 26897 225644 84866
rect 225602 26888 225658 26897
rect 225602 26823 225658 26832
rect 226996 14482 227024 95911
rect 227718 95296 227774 95305
rect 227718 95231 227720 95240
rect 227772 95231 227774 95240
rect 227720 95202 227772 95208
rect 228364 93900 228416 93906
rect 228364 93842 228416 93848
rect 227076 89004 227128 89010
rect 227076 88946 227128 88952
rect 227088 50289 227116 88946
rect 227074 50280 227130 50289
rect 227074 50215 227130 50224
rect 227076 46300 227128 46306
rect 227076 46242 227128 46248
rect 226984 14476 227036 14482
rect 226984 14418 227036 14424
rect 227088 7585 227116 46242
rect 228376 9042 228404 93842
rect 229756 13190 229784 138343
rect 229834 120456 229890 120465
rect 229834 120391 229890 120400
rect 229848 93906 229876 120391
rect 229836 93900 229888 93906
rect 229836 93842 229888 93848
rect 229940 75206 229968 138654
rect 230124 138281 230152 162143
rect 230480 153196 230532 153202
rect 230480 153138 230532 153144
rect 230492 151609 230520 153138
rect 230478 151600 230534 151609
rect 230478 151535 230534 151544
rect 230572 150408 230624 150414
rect 230572 150350 230624 150356
rect 230294 149288 230350 149297
rect 230294 149223 230350 149232
rect 230308 138825 230336 149223
rect 230584 149161 230612 150350
rect 230570 149152 230626 149161
rect 230570 149087 230626 149096
rect 230386 148064 230442 148073
rect 230386 147999 230442 148008
rect 230294 138816 230350 138825
rect 230294 138751 230350 138760
rect 230110 138272 230166 138281
rect 230110 138207 230166 138216
rect 230400 118810 230428 147999
rect 230676 147801 230704 171106
rect 230768 171106 230888 171134
rect 230768 166161 230796 171106
rect 231124 171080 231176 171086
rect 231124 171022 231176 171028
rect 231136 170921 231164 171022
rect 231122 170912 231178 170921
rect 231122 170847 231178 170856
rect 231676 169040 231728 169046
rect 231676 168982 231728 168988
rect 231766 169008 231822 169017
rect 230848 166320 230900 166326
rect 230848 166262 230900 166268
rect 230754 166152 230810 166161
rect 230754 166087 230810 166096
rect 230754 162072 230810 162081
rect 230754 162007 230810 162016
rect 230768 159089 230796 162007
rect 230754 159080 230810 159089
rect 230754 159015 230810 159024
rect 230860 157729 230888 166262
rect 231492 165572 231544 165578
rect 231492 165514 231544 165520
rect 231124 164892 231176 164898
rect 231124 164834 231176 164840
rect 231136 162489 231164 164834
rect 231504 164801 231532 165514
rect 231490 164792 231546 164801
rect 231490 164727 231546 164736
rect 231688 162897 231716 168982
rect 231872 168994 231900 175986
rect 231964 170513 231992 203662
rect 232504 193928 232556 193934
rect 232504 193870 232556 193876
rect 232516 180266 232544 193870
rect 232976 193225 233004 240244
rect 233528 233889 233556 240244
rect 234080 238754 234108 240244
rect 233988 238726 234108 238754
rect 233514 233880 233570 233889
rect 233514 233815 233570 233824
rect 233988 233306 234016 238726
rect 233976 233300 234028 233306
rect 233976 233242 234028 233248
rect 233988 230450 234016 233242
rect 233976 230444 234028 230450
rect 233976 230386 234028 230392
rect 234448 214402 234476 240244
rect 234712 238604 234764 238610
rect 234712 238546 234764 238552
rect 234724 219434 234752 238546
rect 235000 226273 235028 240244
rect 235368 238377 235396 240244
rect 235920 238649 235948 240244
rect 235906 238640 235962 238649
rect 235906 238575 235962 238584
rect 235354 238368 235410 238377
rect 235354 238303 235410 238312
rect 236472 235793 236500 240244
rect 236736 239556 236788 239562
rect 236736 239498 236788 239504
rect 236458 235784 236514 235793
rect 236458 235719 236514 235728
rect 234986 226264 235042 226273
rect 234986 226199 235042 226208
rect 234632 219406 234752 219434
rect 234632 216714 234660 219406
rect 236748 217326 236776 239498
rect 236840 229094 236868 240244
rect 236840 229066 236960 229094
rect 236932 220794 236960 229066
rect 237392 228857 237420 240244
rect 237944 240145 237972 240244
rect 237930 240136 237986 240145
rect 237930 240071 237986 240080
rect 238022 239456 238078 239465
rect 238022 239391 238078 239400
rect 237378 228848 237434 228857
rect 237378 228783 237434 228792
rect 237392 227769 237420 228783
rect 237378 227760 237434 227769
rect 237378 227695 237434 227704
rect 236920 220788 236972 220794
rect 236920 220730 236972 220736
rect 236932 220114 236960 220730
rect 236920 220108 236972 220114
rect 236920 220050 236972 220056
rect 236644 217320 236696 217326
rect 236644 217262 236696 217268
rect 236736 217320 236788 217326
rect 236736 217262 236788 217268
rect 234620 216708 234672 216714
rect 234620 216650 234672 216656
rect 233240 214396 233292 214402
rect 233240 214338 233292 214344
rect 234436 214396 234488 214402
rect 234436 214338 234488 214344
rect 233252 213994 233280 214338
rect 233240 213988 233292 213994
rect 233240 213930 233292 213936
rect 233148 204264 233200 204270
rect 233148 204206 233200 204212
rect 233160 203590 233188 204206
rect 233148 203584 233200 203590
rect 233148 203526 233200 203532
rect 232962 193216 233018 193225
rect 232962 193151 233018 193160
rect 232504 180260 232556 180266
rect 232504 180202 232556 180208
rect 233148 180192 233200 180198
rect 233148 180134 233200 180140
rect 232136 177404 232188 177410
rect 232136 177346 232188 177352
rect 232042 175128 232098 175137
rect 232042 175063 232098 175072
rect 231950 170504 232006 170513
rect 231950 170439 232006 170448
rect 231822 168966 231900 168994
rect 231766 168943 231822 168952
rect 231768 168360 231820 168366
rect 231768 168302 231820 168308
rect 231780 168065 231808 168302
rect 231766 168056 231822 168065
rect 231766 167991 231822 168000
rect 231768 166728 231820 166734
rect 231766 166696 231768 166705
rect 231820 166696 231822 166705
rect 231766 166631 231822 166640
rect 231768 164008 231820 164014
rect 231768 163950 231820 163956
rect 231780 163849 231808 163950
rect 231766 163840 231822 163849
rect 231766 163775 231822 163784
rect 231674 162888 231730 162897
rect 231674 162823 231730 162832
rect 231308 162580 231360 162586
rect 231308 162522 231360 162528
rect 231122 162480 231178 162489
rect 231122 162415 231178 162424
rect 231320 161945 231348 162522
rect 231306 161936 231362 161945
rect 231306 161871 231362 161880
rect 232056 161474 232084 175063
rect 231872 161446 232084 161474
rect 231768 161424 231820 161430
rect 231768 161366 231820 161372
rect 230940 161016 230992 161022
rect 231780 160993 231808 161366
rect 230940 160958 230992 160964
rect 231766 160984 231822 160993
rect 230952 160585 230980 160958
rect 231766 160919 231822 160928
rect 230938 160576 230994 160585
rect 230938 160511 230994 160520
rect 231768 160064 231820 160070
rect 231768 160006 231820 160012
rect 231780 159633 231808 160006
rect 231766 159624 231822 159633
rect 231766 159559 231822 159568
rect 231766 158672 231822 158681
rect 231216 158636 231268 158642
rect 231872 158658 231900 161446
rect 231822 158630 231900 158658
rect 231766 158607 231822 158616
rect 231216 158578 231268 158584
rect 231228 158137 231256 158578
rect 231214 158128 231270 158137
rect 231214 158063 231270 158072
rect 231490 157992 231546 158001
rect 231490 157927 231546 157936
rect 230846 157720 230902 157729
rect 230846 157655 230902 157664
rect 230940 157004 230992 157010
rect 230940 156946 230992 156952
rect 230952 156233 230980 156946
rect 230938 156224 230994 156233
rect 230938 156159 230994 156168
rect 230848 155916 230900 155922
rect 230848 155858 230900 155864
rect 230860 155281 230888 155858
rect 230846 155272 230902 155281
rect 230846 155207 230902 155216
rect 231308 154420 231360 154426
rect 231308 154362 231360 154368
rect 231320 153921 231348 154362
rect 231306 153912 231362 153921
rect 231306 153847 231362 153856
rect 230846 153776 230902 153785
rect 230846 153711 230902 153720
rect 230662 147792 230718 147801
rect 230662 147727 230718 147736
rect 230860 145897 230888 153711
rect 231504 152969 231532 157927
rect 231674 157448 231730 157457
rect 231674 157383 231730 157392
rect 231688 154329 231716 157383
rect 231674 154320 231730 154329
rect 231674 154255 231730 154264
rect 231490 152960 231546 152969
rect 231490 152895 231546 152904
rect 232148 151814 232176 177346
rect 233160 176050 233188 180134
rect 233148 176044 233200 176050
rect 233148 175986 233200 175992
rect 232780 165640 232832 165646
rect 232780 165582 232832 165588
rect 232594 162888 232650 162897
rect 232594 162823 232650 162832
rect 231780 151786 232176 151814
rect 231584 151156 231636 151162
rect 231584 151098 231636 151104
rect 231596 150113 231624 151098
rect 231780 150657 231808 151786
rect 231766 150648 231822 150657
rect 231766 150583 231822 150592
rect 231582 150104 231638 150113
rect 231582 150039 231638 150048
rect 231674 149696 231730 149705
rect 231674 149631 231730 149640
rect 231124 146872 231176 146878
rect 231124 146814 231176 146820
rect 230846 145888 230902 145897
rect 230846 145823 230902 145832
rect 230572 144220 230624 144226
rect 230572 144162 230624 144168
rect 230584 142089 230612 144162
rect 230570 142080 230626 142089
rect 230570 142015 230626 142024
rect 230940 141432 230992 141438
rect 230940 141374 230992 141380
rect 230952 135425 230980 141374
rect 230938 135416 230994 135425
rect 230938 135351 230994 135360
rect 230756 133204 230808 133210
rect 230756 133146 230808 133152
rect 230768 132494 230796 133146
rect 230676 132466 230796 132494
rect 230480 131368 230532 131374
rect 230480 131310 230532 131316
rect 230492 131209 230520 131310
rect 230478 131200 230534 131209
rect 230478 131135 230534 131144
rect 230676 127401 230704 132466
rect 230940 132456 230992 132462
rect 230940 132398 230992 132404
rect 230952 132161 230980 132398
rect 230938 132152 230994 132161
rect 230938 132087 230994 132096
rect 231136 130257 231164 146814
rect 231308 146600 231360 146606
rect 231308 146542 231360 146548
rect 231216 145580 231268 145586
rect 231216 145522 231268 145528
rect 231228 132569 231256 145522
rect 231320 134065 231348 146542
rect 231688 144945 231716 149631
rect 231768 149048 231820 149054
rect 231768 148990 231820 148996
rect 231780 148753 231808 148990
rect 231766 148744 231822 148753
rect 231766 148679 231822 148688
rect 231674 144936 231730 144945
rect 231674 144871 231730 144880
rect 231768 144084 231820 144090
rect 231768 144026 231820 144032
rect 231780 143993 231808 144026
rect 231766 143984 231822 143993
rect 231766 143919 231822 143928
rect 231768 143540 231820 143546
rect 231768 143482 231820 143488
rect 231780 143449 231808 143482
rect 231766 143440 231822 143449
rect 231766 143375 231822 143384
rect 231766 143304 231822 143313
rect 231766 143239 231822 143248
rect 231780 142497 231808 143239
rect 231766 142488 231822 142497
rect 231766 142423 231822 142432
rect 231768 140752 231820 140758
rect 231766 140720 231768 140729
rect 231820 140720 231822 140729
rect 231766 140655 231822 140664
rect 231492 137964 231544 137970
rect 231492 137906 231544 137912
rect 231504 136921 231532 137906
rect 231768 137896 231820 137902
rect 231766 137864 231768 137873
rect 231820 137864 231822 137873
rect 231766 137799 231822 137808
rect 231490 136912 231546 136921
rect 231490 136847 231546 136856
rect 231768 136604 231820 136610
rect 231768 136546 231820 136552
rect 231676 136536 231728 136542
rect 231676 136478 231728 136484
rect 231688 135969 231716 136478
rect 231780 136377 231808 136546
rect 231766 136368 231822 136377
rect 231766 136303 231822 136312
rect 231674 135960 231730 135969
rect 231674 135895 231730 135904
rect 231768 135244 231820 135250
rect 231768 135186 231820 135192
rect 231676 135176 231728 135182
rect 231676 135118 231728 135124
rect 231688 134473 231716 135118
rect 231780 135017 231808 135186
rect 231766 135008 231822 135017
rect 231766 134943 231822 134952
rect 231674 134464 231730 134473
rect 231674 134399 231730 134408
rect 231306 134056 231362 134065
rect 231306 133991 231362 134000
rect 231492 133884 231544 133890
rect 231492 133826 231544 133832
rect 231504 133113 231532 133826
rect 231490 133104 231546 133113
rect 231490 133039 231546 133048
rect 231214 132560 231270 132569
rect 231214 132495 231270 132504
rect 231768 131096 231820 131102
rect 231768 131038 231820 131044
rect 231492 131028 231544 131034
rect 231492 130970 231544 130976
rect 231306 130384 231362 130393
rect 231306 130319 231362 130328
rect 231122 130248 231178 130257
rect 231122 130183 231178 130192
rect 230754 129024 230810 129033
rect 230754 128959 230810 128968
rect 230662 127392 230718 127401
rect 230662 127327 230718 127336
rect 230768 126993 230796 128959
rect 230754 126984 230810 126993
rect 230754 126919 230810 126928
rect 231214 126304 231270 126313
rect 231124 126268 231176 126274
rect 231214 126239 231270 126248
rect 231124 126210 231176 126216
rect 230848 124976 230900 124982
rect 230848 124918 230900 124924
rect 230664 123480 230716 123486
rect 230664 123422 230716 123428
rect 230676 118969 230704 123422
rect 230756 122528 230808 122534
rect 230756 122470 230808 122476
rect 230768 122233 230796 122470
rect 230754 122224 230810 122233
rect 230754 122159 230810 122168
rect 230662 118960 230718 118969
rect 230662 118895 230718 118904
rect 230400 118782 230520 118810
rect 230492 106185 230520 118782
rect 230860 116113 230888 124918
rect 230940 124908 230992 124914
rect 230940 124850 230992 124856
rect 230952 123185 230980 124850
rect 230938 123176 230994 123185
rect 230938 123111 230994 123120
rect 230846 116104 230902 116113
rect 230846 116039 230902 116048
rect 230572 114640 230624 114646
rect 231136 114617 231164 126210
rect 231228 120737 231256 126239
rect 231320 125089 231348 130319
rect 231504 129849 231532 130970
rect 231780 130665 231808 131038
rect 231766 130656 231822 130665
rect 231766 130591 231822 130600
rect 231490 129840 231546 129849
rect 231490 129775 231546 129784
rect 231768 129736 231820 129742
rect 231768 129678 231820 129684
rect 231492 129600 231544 129606
rect 231492 129542 231544 129548
rect 231504 128897 231532 129542
rect 231780 129305 231808 129678
rect 231766 129296 231822 129305
rect 231766 129231 231822 129240
rect 231490 128888 231546 128897
rect 231490 128823 231546 128832
rect 231766 128344 231822 128353
rect 231766 128279 231768 128288
rect 231820 128279 231822 128288
rect 231768 128250 231820 128256
rect 231676 128240 231728 128246
rect 231676 128182 231728 128188
rect 231688 127945 231716 128182
rect 231674 127936 231730 127945
rect 231674 127871 231730 127880
rect 231768 126948 231820 126954
rect 231768 126890 231820 126896
rect 231780 126041 231808 126890
rect 231766 126032 231822 126041
rect 231766 125967 231822 125976
rect 232502 126032 232558 126041
rect 232502 125967 232558 125976
rect 231306 125080 231362 125089
rect 231306 125015 231362 125024
rect 231768 123888 231820 123894
rect 231768 123830 231820 123836
rect 231780 123593 231808 123830
rect 231766 123584 231822 123593
rect 231766 123519 231822 123528
rect 231584 122732 231636 122738
rect 231584 122674 231636 122680
rect 231596 121689 231624 122674
rect 231582 121680 231638 121689
rect 231582 121615 231638 121624
rect 231768 121440 231820 121446
rect 231768 121382 231820 121388
rect 231780 121281 231808 121382
rect 231766 121272 231822 121281
rect 231766 121207 231822 121216
rect 231676 120964 231728 120970
rect 231676 120906 231728 120912
rect 231214 120728 231270 120737
rect 231214 120663 231270 120672
rect 231688 120329 231716 120906
rect 231674 120320 231730 120329
rect 231674 120255 231730 120264
rect 231768 120080 231820 120086
rect 231768 120022 231820 120028
rect 231780 119377 231808 120022
rect 231766 119368 231822 119377
rect 231766 119303 231822 119312
rect 231216 118720 231268 118726
rect 231216 118662 231268 118668
rect 230572 114582 230624 114588
rect 231122 114608 231178 114617
rect 230584 113665 230612 114582
rect 231122 114543 231178 114552
rect 230846 113792 230902 113801
rect 230846 113727 230902 113736
rect 230570 113656 230626 113665
rect 230570 113591 230626 113600
rect 230756 111784 230808 111790
rect 230756 111726 230808 111732
rect 230768 110809 230796 111726
rect 230754 110800 230810 110809
rect 230754 110735 230810 110744
rect 230860 109449 230888 113727
rect 231228 111353 231256 118662
rect 231400 118652 231452 118658
rect 231400 118594 231452 118600
rect 231412 118017 231440 118594
rect 231398 118008 231454 118017
rect 231398 117943 231454 117952
rect 231492 117700 231544 117706
rect 231492 117642 231544 117648
rect 231504 117473 231532 117642
rect 231490 117464 231546 117473
rect 231490 117399 231546 117408
rect 231768 117292 231820 117298
rect 231768 117234 231820 117240
rect 231780 117065 231808 117234
rect 231766 117056 231822 117065
rect 231766 116991 231822 117000
rect 231676 116884 231728 116890
rect 231676 116826 231728 116832
rect 231688 116521 231716 116826
rect 231674 116512 231730 116521
rect 231674 116447 231730 116456
rect 231492 115932 231544 115938
rect 231492 115874 231544 115880
rect 231504 115161 231532 115874
rect 231490 115152 231546 115161
rect 231490 115087 231546 115096
rect 231768 114504 231820 114510
rect 231768 114446 231820 114452
rect 231492 114436 231544 114442
rect 231492 114378 231544 114384
rect 231504 113257 231532 114378
rect 231780 114209 231808 114446
rect 231766 114200 231822 114209
rect 231766 114135 231822 114144
rect 231490 113248 231546 113257
rect 231490 113183 231546 113192
rect 231768 113144 231820 113150
rect 231768 113086 231820 113092
rect 231400 113076 231452 113082
rect 231400 113018 231452 113024
rect 231412 112305 231440 113018
rect 231780 112713 231808 113086
rect 231766 112704 231822 112713
rect 231766 112639 231822 112648
rect 231398 112296 231454 112305
rect 231398 112231 231454 112240
rect 231214 111344 231270 111353
rect 231214 111279 231270 111288
rect 231584 111104 231636 111110
rect 231490 111072 231546 111081
rect 231584 111046 231636 111052
rect 231490 111007 231546 111016
rect 231504 109857 231532 111007
rect 231490 109848 231546 109857
rect 231490 109783 231546 109792
rect 231400 109744 231452 109750
rect 231400 109686 231452 109692
rect 230846 109440 230902 109449
rect 230846 109375 230902 109384
rect 231308 107636 231360 107642
rect 231308 107578 231360 107584
rect 231320 107137 231348 107578
rect 231306 107128 231362 107137
rect 231306 107063 231362 107072
rect 231412 106570 231440 109686
rect 231596 109154 231624 111046
rect 231768 110424 231820 110430
rect 231766 110392 231768 110401
rect 231820 110392 231822 110401
rect 231766 110327 231822 110336
rect 231320 106542 231440 106570
rect 231504 109126 231624 109154
rect 230478 106176 230534 106185
rect 230478 106111 230534 106120
rect 231214 105496 231270 105505
rect 231214 105431 231270 105440
rect 231124 104372 231176 104378
rect 231124 104314 231176 104320
rect 231136 103737 231164 104314
rect 231122 103728 231178 103737
rect 231122 103663 231178 103672
rect 231032 102808 231084 102814
rect 231032 102750 231084 102756
rect 230572 102060 230624 102066
rect 230572 102002 230624 102008
rect 230584 101833 230612 102002
rect 230570 101824 230626 101833
rect 230570 101759 230626 101768
rect 230572 100700 230624 100706
rect 230572 100642 230624 100648
rect 230584 100473 230612 100642
rect 230570 100464 230626 100473
rect 230570 100399 230626 100408
rect 230478 97064 230534 97073
rect 230478 96999 230534 97008
rect 230492 95690 230520 96999
rect 230570 96248 230626 96257
rect 230570 96183 230626 96192
rect 230584 95878 230612 96183
rect 230572 95872 230624 95878
rect 230572 95814 230624 95820
rect 230492 95662 230612 95690
rect 230584 95266 230612 95662
rect 230572 95260 230624 95266
rect 230572 95202 230624 95208
rect 230584 93854 230612 95202
rect 230492 93826 230612 93854
rect 231044 93854 231072 102750
rect 231124 100632 231176 100638
rect 231124 100574 231176 100580
rect 231136 99521 231164 100574
rect 231122 99512 231178 99521
rect 231122 99447 231178 99456
rect 231124 99340 231176 99346
rect 231124 99282 231176 99288
rect 231136 98569 231164 99282
rect 231122 98560 231178 98569
rect 231122 98495 231178 98504
rect 231044 93826 231164 93854
rect 230492 93770 230520 93826
rect 230480 93764 230532 93770
rect 230480 93706 230532 93712
rect 229928 75200 229980 75206
rect 229928 75142 229980 75148
rect 230492 39438 230520 93706
rect 230480 39432 230532 39438
rect 230480 39374 230532 39380
rect 231136 22778 231164 93826
rect 231228 57254 231256 105431
rect 231320 99929 231348 106542
rect 231400 106276 231452 106282
rect 231400 106218 231452 106224
rect 231412 105641 231440 106218
rect 231398 105632 231454 105641
rect 231398 105567 231454 105576
rect 231504 103514 231532 109126
rect 231584 108996 231636 109002
rect 231584 108938 231636 108944
rect 231596 107953 231624 108938
rect 231768 108588 231820 108594
rect 231768 108530 231820 108536
rect 231780 108497 231808 108530
rect 231766 108488 231822 108497
rect 231766 108423 231822 108432
rect 231582 107944 231638 107953
rect 231582 107879 231638 107888
rect 231768 107568 231820 107574
rect 231768 107510 231820 107516
rect 231780 106593 231808 107510
rect 231766 106584 231822 106593
rect 231766 106519 231822 106528
rect 231768 106208 231820 106214
rect 231768 106150 231820 106156
rect 231780 105233 231808 106150
rect 231766 105224 231822 105233
rect 231766 105159 231822 105168
rect 231768 104780 231820 104786
rect 231768 104722 231820 104728
rect 231780 104281 231808 104722
rect 231766 104272 231822 104281
rect 231766 104207 231822 104216
rect 231412 103486 231532 103514
rect 231768 103488 231820 103494
rect 231412 102377 231440 103486
rect 231768 103430 231820 103436
rect 231780 102785 231808 103430
rect 231766 102776 231822 102785
rect 231766 102711 231822 102720
rect 231398 102368 231454 102377
rect 231398 102303 231454 102312
rect 231676 102128 231728 102134
rect 231676 102070 231728 102076
rect 231766 102096 231822 102105
rect 231688 100881 231716 102070
rect 231766 102031 231822 102040
rect 231780 101425 231808 102031
rect 231766 101416 231822 101425
rect 231766 101351 231822 101360
rect 231674 100872 231730 100881
rect 231674 100807 231730 100816
rect 231306 99920 231362 99929
rect 231306 99855 231362 99864
rect 231676 98660 231728 98666
rect 231676 98602 231728 98608
rect 231688 96665 231716 98602
rect 231768 97980 231820 97986
rect 231768 97922 231820 97928
rect 231780 97617 231808 97922
rect 231766 97608 231822 97617
rect 231766 97543 231822 97552
rect 231674 96656 231730 96665
rect 231674 96591 231730 96600
rect 231216 57248 231268 57254
rect 231216 57190 231268 57196
rect 231216 43444 231268 43450
rect 231216 43386 231268 43392
rect 231124 22772 231176 22778
rect 231124 22714 231176 22720
rect 229744 13184 229796 13190
rect 229744 13126 229796 13132
rect 228364 9036 228416 9042
rect 228364 8978 228416 8984
rect 227074 7576 227130 7585
rect 227074 7511 227130 7520
rect 224316 6248 224368 6254
rect 224316 6190 224368 6196
rect 222936 2780 222988 2786
rect 222936 2722 222988 2728
rect 231228 2106 231256 43386
rect 232516 35193 232544 125967
rect 232608 122534 232636 162823
rect 232686 155000 232742 155009
rect 232686 154935 232742 154944
rect 232596 122528 232648 122534
rect 232596 122470 232648 122476
rect 232700 114646 232728 154935
rect 232792 126449 232820 165582
rect 233252 161022 233280 213930
rect 233332 181552 233384 181558
rect 233332 181494 233384 181500
rect 233240 161016 233292 161022
rect 233240 160958 233292 160964
rect 233344 155961 233372 181494
rect 233422 180160 233478 180169
rect 233422 180095 233478 180104
rect 233436 157010 233464 180095
rect 233514 176080 233570 176089
rect 233514 176015 233570 176024
rect 233528 171086 233556 176015
rect 233516 171080 233568 171086
rect 233516 171022 233568 171028
rect 233976 169788 234028 169794
rect 233976 169730 234028 169736
rect 233884 158772 233936 158778
rect 233884 158714 233936 158720
rect 233424 157004 233476 157010
rect 233424 156946 233476 156952
rect 233330 155952 233386 155961
rect 233330 155887 233386 155896
rect 232872 151088 232924 151094
rect 232872 151030 232924 151036
rect 232778 126440 232834 126449
rect 232778 126375 232834 126384
rect 232884 124545 232912 151030
rect 232870 124536 232926 124545
rect 232870 124471 232926 124480
rect 232778 121816 232834 121825
rect 232778 121751 232834 121760
rect 232688 114640 232740 114646
rect 232688 114582 232740 114588
rect 232686 109712 232742 109721
rect 232686 109647 232742 109656
rect 232596 95872 232648 95878
rect 232596 95814 232648 95820
rect 232502 35184 232558 35193
rect 232502 35119 232558 35128
rect 232608 5574 232636 95814
rect 232700 84930 232728 109647
rect 232792 90438 232820 121751
rect 233896 118425 233924 158714
rect 233988 131374 234016 169730
rect 234160 153876 234212 153882
rect 234160 153818 234212 153824
rect 234068 148368 234120 148374
rect 234068 148310 234120 148316
rect 233976 131368 234028 131374
rect 233976 131310 234028 131316
rect 233882 118416 233938 118425
rect 233882 118351 233938 118360
rect 233882 116240 233938 116249
rect 233882 116175 233938 116184
rect 232780 90432 232832 90438
rect 232780 90374 232832 90380
rect 232688 84924 232740 84930
rect 232688 84866 232740 84872
rect 233896 7614 233924 116175
rect 234080 111790 234108 148310
rect 234172 125497 234200 153818
rect 234632 153202 234660 216650
rect 234712 189168 234764 189174
rect 234712 189110 234764 189116
rect 234724 165753 234752 189110
rect 236092 188352 236144 188358
rect 236092 188294 236144 188300
rect 236000 184272 236052 184278
rect 236000 184214 236052 184220
rect 236012 181558 236040 184214
rect 236000 181552 236052 181558
rect 236000 181494 236052 181500
rect 234802 177304 234858 177313
rect 234802 177239 234858 177248
rect 234710 165744 234766 165753
rect 234710 165679 234766 165688
rect 234816 157457 234844 177239
rect 236000 176180 236052 176186
rect 236000 176122 236052 176128
rect 234894 168736 234950 168745
rect 234894 168671 234950 168680
rect 234908 166734 234936 168671
rect 234896 166728 234948 166734
rect 234896 166670 234948 166676
rect 235540 162920 235592 162926
rect 235540 162862 235592 162868
rect 234802 157448 234858 157457
rect 234802 157383 234858 157392
rect 235264 157412 235316 157418
rect 235264 157354 235316 157360
rect 234620 153196 234672 153202
rect 234620 153138 234672 153144
rect 234158 125488 234214 125497
rect 234158 125423 234214 125432
rect 234158 117872 234214 117881
rect 234158 117807 234214 117816
rect 234068 111784 234120 111790
rect 234068 111726 234120 111732
rect 233974 104000 234030 104009
rect 233974 103935 234030 103944
rect 233988 29646 234016 103935
rect 234172 89078 234200 117807
rect 235276 116890 235304 157354
rect 235356 144968 235408 144974
rect 235356 144910 235408 144916
rect 235264 116884 235316 116890
rect 235264 116826 235316 116832
rect 235262 114880 235318 114889
rect 235262 114815 235318 114824
rect 234160 89072 234212 89078
rect 234160 89014 234212 89020
rect 233976 29640 234028 29646
rect 233976 29582 234028 29588
rect 235276 21418 235304 114815
rect 235368 104378 235396 144910
rect 235446 124672 235502 124681
rect 235446 124607 235502 124616
rect 235356 104372 235408 104378
rect 235356 104314 235408 104320
rect 235354 98696 235410 98705
rect 235354 98631 235410 98640
rect 235368 42090 235396 98631
rect 235460 80714 235488 124607
rect 235552 123894 235580 162862
rect 236012 155922 236040 176122
rect 236104 169561 236132 188294
rect 236182 178800 236238 178809
rect 236182 178735 236238 178744
rect 236090 169552 236146 169561
rect 236090 169487 236146 169496
rect 236092 166320 236144 166326
rect 236092 166262 236144 166268
rect 236104 164014 236132 166262
rect 236092 164008 236144 164014
rect 236092 163950 236144 163956
rect 236196 163441 236224 178735
rect 236656 176089 236684 217262
rect 237380 211200 237432 211206
rect 237380 211142 237432 211148
rect 237392 210905 237420 211142
rect 237378 210896 237434 210905
rect 237378 210831 237434 210840
rect 236734 198792 236790 198801
rect 236734 198727 236790 198736
rect 236748 188358 236776 198727
rect 237472 195288 237524 195294
rect 237472 195230 237524 195236
rect 237380 192568 237432 192574
rect 237380 192510 237432 192516
rect 236736 188352 236788 188358
rect 236736 188294 236788 188300
rect 236642 176080 236698 176089
rect 236642 176015 236698 176024
rect 236828 169856 236880 169862
rect 236828 169798 236880 169804
rect 236182 163432 236238 163441
rect 236182 163367 236238 163376
rect 236736 162172 236788 162178
rect 236736 162114 236788 162120
rect 236644 156664 236696 156670
rect 236644 156606 236696 156612
rect 236000 155916 236052 155922
rect 236000 155858 236052 155864
rect 235540 123888 235592 123894
rect 235540 123830 235592 123836
rect 236656 117706 236684 156606
rect 236748 129606 236776 162114
rect 236840 146878 236868 169798
rect 237392 154426 237420 192510
rect 237484 169969 237512 195230
rect 238036 193866 238064 239391
rect 238114 227760 238170 227769
rect 238114 227695 238170 227704
rect 238128 214606 238156 227695
rect 238116 214600 238168 214606
rect 238116 214542 238168 214548
rect 238312 211206 238340 240244
rect 238760 239488 238812 239494
rect 238760 239430 238812 239436
rect 238772 238678 238800 239430
rect 238760 238672 238812 238678
rect 238760 238614 238812 238620
rect 238864 218754 238892 240244
rect 239232 240009 239260 240244
rect 239218 240000 239274 240009
rect 239218 239935 239274 239944
rect 238942 236600 238998 236609
rect 238942 236535 238998 236544
rect 238852 218748 238904 218754
rect 238852 218690 238904 218696
rect 238300 211200 238352 211206
rect 238300 211142 238352 211148
rect 238116 208412 238168 208418
rect 238116 208354 238168 208360
rect 238024 193860 238076 193866
rect 238024 193802 238076 193808
rect 238128 187241 238156 208354
rect 238114 187232 238170 187241
rect 238114 187167 238170 187176
rect 237564 186992 237616 186998
rect 237564 186934 237616 186940
rect 237470 169960 237526 169969
rect 237470 169895 237526 169904
rect 237576 162586 237604 186934
rect 238760 182912 238812 182918
rect 238760 182854 238812 182860
rect 238208 172576 238260 172582
rect 238208 172518 238260 172524
rect 237564 162580 237616 162586
rect 237564 162522 237616 162528
rect 238024 160132 238076 160138
rect 238024 160074 238076 160080
rect 237380 154420 237432 154426
rect 237380 154362 237432 154368
rect 236918 150104 236974 150113
rect 236918 150039 236974 150048
rect 236828 146872 236880 146878
rect 236828 146814 236880 146820
rect 236828 140820 236880 140826
rect 236828 140762 236880 140768
rect 236736 129600 236788 129606
rect 236736 129542 236788 129548
rect 236644 117700 236696 117706
rect 236644 117642 236696 117648
rect 236644 116000 236696 116006
rect 236644 115942 236696 115948
rect 235448 80708 235500 80714
rect 235448 80650 235500 80656
rect 236656 49026 236684 115942
rect 236736 108316 236788 108322
rect 236736 108258 236788 108264
rect 236644 49020 236696 49026
rect 236644 48962 236696 48968
rect 236748 44946 236776 108258
rect 236840 99346 236868 140762
rect 236932 108594 236960 150039
rect 238036 120970 238064 160074
rect 238116 151836 238168 151842
rect 238116 151778 238168 151784
rect 238024 120964 238076 120970
rect 238024 120906 238076 120912
rect 238022 119096 238078 119105
rect 238022 119031 238078 119040
rect 236920 108588 236972 108594
rect 236920 108530 236972 108536
rect 236918 100056 236974 100065
rect 236918 99991 236974 100000
rect 236828 99340 236880 99346
rect 236828 99282 236880 99288
rect 236932 86290 236960 99991
rect 236920 86284 236972 86290
rect 236920 86226 236972 86232
rect 236736 44940 236788 44946
rect 236736 44882 236788 44888
rect 235356 42084 235408 42090
rect 235356 42026 235408 42032
rect 235264 21412 235316 21418
rect 235264 21354 235316 21360
rect 238036 7682 238064 119031
rect 238128 118726 238156 151778
rect 238220 146606 238248 172518
rect 238392 169108 238444 169114
rect 238392 169050 238444 169056
rect 238208 146600 238260 146606
rect 238208 146542 238260 146548
rect 238298 146432 238354 146441
rect 238298 146367 238354 146376
rect 238208 142180 238260 142186
rect 238208 142122 238260 142128
rect 238116 118720 238168 118726
rect 238116 118662 238168 118668
rect 238116 103556 238168 103562
rect 238116 103498 238168 103504
rect 238128 26994 238156 103498
rect 238220 100638 238248 142122
rect 238312 104786 238340 146367
rect 238404 144090 238432 169050
rect 238772 153377 238800 182854
rect 238852 177336 238904 177342
rect 238852 177278 238904 177284
rect 238864 153785 238892 177278
rect 238850 153776 238906 153785
rect 238850 153711 238906 153720
rect 238758 153368 238814 153377
rect 238758 153303 238814 153312
rect 238392 144084 238444 144090
rect 238392 144026 238444 144032
rect 238956 141137 238984 236535
rect 239784 224913 239812 240244
rect 240140 238808 240192 238814
rect 240140 238750 240192 238756
rect 240152 234598 240180 238750
rect 240336 238746 240364 240244
rect 240324 238740 240376 238746
rect 240324 238682 240376 238688
rect 240336 237454 240364 238682
rect 240324 237448 240376 237454
rect 240324 237390 240376 237396
rect 240140 234592 240192 234598
rect 240140 234534 240192 234540
rect 240704 226302 240732 240244
rect 240874 239864 240930 239873
rect 240874 239799 240930 239808
rect 240784 237448 240836 237454
rect 240784 237390 240836 237396
rect 240692 226296 240744 226302
rect 240692 226238 240744 226244
rect 239770 224904 239826 224913
rect 239770 224839 239826 224848
rect 240138 213344 240194 213353
rect 240138 213279 240194 213288
rect 239404 180124 239456 180130
rect 239404 180066 239456 180072
rect 239034 173904 239090 173913
rect 239416 173874 239444 180066
rect 239034 173839 239090 173848
rect 239404 173868 239456 173874
rect 239048 167686 239076 173839
rect 239404 173810 239456 173816
rect 239036 167680 239088 167686
rect 239036 167622 239088 167628
rect 239496 167068 239548 167074
rect 239496 167010 239548 167016
rect 238942 141128 238998 141137
rect 238942 141063 238998 141072
rect 239402 137184 239458 137193
rect 239402 137119 239458 137128
rect 238392 117972 238444 117978
rect 238392 117914 238444 117920
rect 238300 104780 238352 104786
rect 238300 104722 238352 104728
rect 238208 100632 238260 100638
rect 238208 100574 238260 100580
rect 238404 79354 238432 117914
rect 238392 79348 238444 79354
rect 238392 79290 238444 79296
rect 239416 50386 239444 137119
rect 239508 133210 239536 167010
rect 240152 158642 240180 213279
rect 240230 204232 240286 204241
rect 240230 204167 240286 204176
rect 240244 172514 240272 204167
rect 240796 188426 240824 237390
rect 240888 206961 240916 239799
rect 241256 238814 241284 240244
rect 241244 238808 241296 238814
rect 241244 238750 241296 238756
rect 241808 238746 241836 240244
rect 241796 238740 241848 238746
rect 241796 238682 241848 238688
rect 241808 237862 241836 238682
rect 242176 238649 242204 240244
rect 242256 240100 242308 240106
rect 242256 240042 242308 240048
rect 242162 238640 242218 238649
rect 242162 238575 242218 238584
rect 241796 237856 241848 237862
rect 241796 237798 241848 237804
rect 242176 237425 242204 238575
rect 241610 237416 241666 237425
rect 241610 237351 241666 237360
rect 242162 237416 242218 237425
rect 242162 237351 242218 237360
rect 240968 225004 241020 225010
rect 240968 224946 241020 224952
rect 240874 206952 240930 206961
rect 240874 206887 240930 206896
rect 240980 204241 241008 224946
rect 241520 216640 241572 216646
rect 241520 216582 241572 216588
rect 240966 204232 241022 204241
rect 240966 204167 241022 204176
rect 240784 188420 240836 188426
rect 240784 188362 240836 188368
rect 241426 187776 241482 187785
rect 241426 187711 241482 187720
rect 240874 172816 240930 172825
rect 240874 172751 240930 172760
rect 240232 172508 240284 172514
rect 240232 172450 240284 172456
rect 240232 171828 240284 171834
rect 240232 171770 240284 171776
rect 240244 168366 240272 171770
rect 240784 171148 240836 171154
rect 240784 171090 240836 171096
rect 240232 168360 240284 168366
rect 240232 168302 240284 168308
rect 240140 158636 240192 158642
rect 240140 158578 240192 158584
rect 239586 153232 239642 153241
rect 239586 153167 239642 153176
rect 239496 133204 239548 133210
rect 239496 133146 239548 133152
rect 239494 112160 239550 112169
rect 239494 112095 239550 112104
rect 239508 68377 239536 112095
rect 239600 111761 239628 153167
rect 239680 146940 239732 146946
rect 239680 146882 239732 146888
rect 239586 111752 239642 111761
rect 239586 111687 239642 111696
rect 239692 107574 239720 146882
rect 240796 145586 240824 171090
rect 240888 155281 240916 172751
rect 241440 172417 241468 187711
rect 241426 172408 241482 172417
rect 241426 172343 241482 172352
rect 241152 157480 241204 157486
rect 241152 157422 241204 157428
rect 240874 155272 240930 155281
rect 240874 155207 240930 155216
rect 241060 154624 241112 154630
rect 241060 154566 241112 154572
rect 240784 145580 240836 145586
rect 240784 145522 240836 145528
rect 240968 145036 241020 145042
rect 240968 144978 241020 144984
rect 240784 140072 240836 140078
rect 240784 140014 240836 140020
rect 240796 126313 240824 140014
rect 240782 126304 240838 126313
rect 240782 126239 240838 126248
rect 240876 122868 240928 122874
rect 240876 122810 240928 122816
rect 240784 116068 240836 116074
rect 240784 116010 240836 116016
rect 239680 107568 239732 107574
rect 239680 107510 239732 107516
rect 239586 106856 239642 106865
rect 239586 106791 239642 106800
rect 239600 83502 239628 106791
rect 240140 95260 240192 95266
rect 240140 95202 240192 95208
rect 240152 93770 240180 95202
rect 240140 93764 240192 93770
rect 240140 93706 240192 93712
rect 239588 83496 239640 83502
rect 239588 83438 239640 83444
rect 239494 68368 239550 68377
rect 239494 68303 239550 68312
rect 240140 51808 240192 51814
rect 240140 51750 240192 51756
rect 239404 50380 239456 50386
rect 239404 50322 239456 50328
rect 238116 26988 238168 26994
rect 238116 26930 238168 26936
rect 238024 7676 238076 7682
rect 238024 7618 238076 7624
rect 233884 7608 233936 7614
rect 233884 7550 233936 7556
rect 239310 6216 239366 6225
rect 239310 6151 239366 6160
rect 232596 5568 232648 5574
rect 232596 5510 232648 5516
rect 235816 5568 235868 5574
rect 235816 5510 235868 5516
rect 231216 2100 231268 2106
rect 231216 2042 231268 2048
rect 200854 2000 200910 2009
rect 200854 1935 200910 1944
rect 235828 480 235856 5510
rect 239324 480 239352 6151
rect 240152 490 240180 51750
rect 240796 4826 240824 116010
rect 240888 76566 240916 122810
rect 240980 103494 241008 144978
rect 241072 114442 241100 154566
rect 241164 117298 241192 157422
rect 241532 150414 241560 216582
rect 241624 169114 241652 237351
rect 242268 216646 242296 240042
rect 242440 237856 242492 237862
rect 242440 237798 242492 237804
rect 242256 216640 242308 216646
rect 242256 216582 242308 216588
rect 242452 187785 242480 237798
rect 242728 235929 242756 240244
rect 242808 240168 242860 240174
rect 242808 240110 242860 240116
rect 242820 238513 242848 240110
rect 242806 238504 242862 238513
rect 242806 238439 242862 238448
rect 242714 235920 242770 235929
rect 242714 235855 242770 235864
rect 243280 225010 243308 240244
rect 243648 231810 243676 240244
rect 243924 238678 243952 243222
rect 244002 243199 244058 243208
rect 244002 241360 244058 241369
rect 244002 241295 244058 241304
rect 244016 239873 244044 241295
rect 244002 239864 244058 239873
rect 244002 239799 244058 239808
rect 243912 238672 243964 238678
rect 243912 238614 243964 238620
rect 243636 231804 243688 231810
rect 243636 231746 243688 231752
rect 243268 225004 243320 225010
rect 243268 224946 243320 224952
rect 243648 219434 243676 231746
rect 243726 228304 243782 228313
rect 243726 228239 243782 228248
rect 243556 219406 243676 219434
rect 242438 187776 242494 187785
rect 242438 187711 242494 187720
rect 241704 180260 241756 180266
rect 241704 180202 241756 180208
rect 241612 169108 241664 169114
rect 241612 169050 241664 169056
rect 241716 160070 241744 180202
rect 243556 178702 243584 219406
rect 242900 178696 242952 178702
rect 242900 178638 242952 178644
rect 243544 178696 243596 178702
rect 243544 178638 243596 178644
rect 242256 168428 242308 168434
rect 242256 168370 242308 168376
rect 241704 160064 241756 160070
rect 241704 160006 241756 160012
rect 242164 151904 242216 151910
rect 242164 151846 242216 151852
rect 241520 150408 241572 150414
rect 241520 150350 241572 150356
rect 241152 117292 241204 117298
rect 241152 117234 241204 117240
rect 241060 114436 241112 114442
rect 241060 114378 241112 114384
rect 242176 110430 242204 151846
rect 242268 131034 242296 168370
rect 242440 155984 242492 155990
rect 242440 155926 242492 155932
rect 242348 143608 242400 143614
rect 242348 143550 242400 143556
rect 242256 131028 242308 131034
rect 242256 130970 242308 130976
rect 242164 110424 242216 110430
rect 242164 110366 242216 110372
rect 242256 109064 242308 109070
rect 242256 109006 242308 109012
rect 240968 103488 241020 103494
rect 240968 103430 241020 103436
rect 241060 102876 241112 102882
rect 241060 102818 241112 102824
rect 241072 93265 241100 102818
rect 242162 101144 242218 101153
rect 242162 101079 242218 101088
rect 241058 93256 241114 93265
rect 241058 93191 241114 93200
rect 240876 76560 240928 76566
rect 240876 76502 240928 76508
rect 241520 43512 241572 43518
rect 241520 43454 241572 43460
rect 241532 16574 241560 43454
rect 242176 37942 242204 101079
rect 242268 54534 242296 109006
rect 242360 102066 242388 143550
rect 242452 124982 242480 155926
rect 242912 137902 242940 178638
rect 243740 175953 243768 228239
rect 244292 205630 244320 250815
rect 244462 247344 244518 247353
rect 244462 247279 244518 247288
rect 244370 240816 244426 240825
rect 244370 240751 244426 240760
rect 244384 229094 244412 240751
rect 244476 230353 244504 247279
rect 244462 230344 244518 230353
rect 244462 230279 244518 230288
rect 244384 229066 244504 229094
rect 244476 209778 244504 229066
rect 244464 209772 244516 209778
rect 244464 209714 244516 209720
rect 244280 205624 244332 205630
rect 244280 205566 244332 205572
rect 244292 205193 244320 205566
rect 244278 205184 244334 205193
rect 244278 205119 244334 205128
rect 244280 198552 244332 198558
rect 244280 198494 244332 198500
rect 243820 183796 243872 183802
rect 243820 183738 243872 183744
rect 243726 175944 243782 175953
rect 243726 175879 243782 175888
rect 243636 175296 243688 175302
rect 243636 175238 243688 175244
rect 242992 173936 243044 173942
rect 242992 173878 243044 173884
rect 243004 161430 243032 173878
rect 242992 161424 243044 161430
rect 242992 161366 243044 161372
rect 242900 137896 242952 137902
rect 242900 137838 242952 137844
rect 242440 124976 242492 124982
rect 242440 124918 242492 124924
rect 243544 124228 243596 124234
rect 243544 124170 243596 124176
rect 242348 102060 242400 102066
rect 242348 102002 242400 102008
rect 242256 54528 242308 54534
rect 242256 54470 242308 54476
rect 242164 37936 242216 37942
rect 242164 37878 242216 37884
rect 243556 32502 243584 124170
rect 243648 111217 243676 175238
rect 243832 143546 243860 183738
rect 244292 172281 244320 198494
rect 244476 176089 244504 209714
rect 244936 198558 244964 264143
rect 245842 263120 245898 263129
rect 245842 263055 245898 263064
rect 245014 258768 245070 258777
rect 245014 258703 245070 258712
rect 245028 246362 245056 258703
rect 245658 256592 245714 256601
rect 245658 256527 245714 256536
rect 245672 256086 245700 256527
rect 245660 256080 245712 256086
rect 245660 256022 245712 256028
rect 245660 253224 245712 253230
rect 245660 253166 245712 253172
rect 245672 253065 245700 253166
rect 245658 253056 245714 253065
rect 245658 252991 245714 253000
rect 245660 250504 245712 250510
rect 245660 250446 245712 250452
rect 245672 250345 245700 250446
rect 245658 250336 245714 250345
rect 245658 250271 245714 250280
rect 245750 248704 245806 248713
rect 245750 248639 245806 248648
rect 245016 246356 245068 246362
rect 245016 246298 245068 246304
rect 245658 245168 245714 245177
rect 245658 245103 245714 245112
rect 245672 240106 245700 245103
rect 245660 240100 245712 240106
rect 245660 240042 245712 240048
rect 245660 214668 245712 214674
rect 245660 214610 245712 214616
rect 244924 198552 244976 198558
rect 244924 198494 244976 198500
rect 244462 176080 244518 176089
rect 244372 176044 244424 176050
rect 244462 176015 244518 176024
rect 244372 175986 244424 175992
rect 244278 172272 244334 172281
rect 244278 172207 244334 172216
rect 244384 165578 244412 175986
rect 245016 173936 245068 173942
rect 245016 173878 245068 173884
rect 244922 171592 244978 171601
rect 244922 171527 244978 171536
rect 244372 165572 244424 165578
rect 244372 165514 244424 165520
rect 243912 158840 243964 158846
rect 243912 158782 243964 158788
rect 243820 143540 243872 143546
rect 243820 143482 243872 143488
rect 243728 136672 243780 136678
rect 243728 136614 243780 136620
rect 243634 111208 243690 111217
rect 243634 111143 243690 111152
rect 243740 80889 243768 136614
rect 243924 123486 243952 158782
rect 244936 132462 244964 171527
rect 245028 136542 245056 173878
rect 245106 167104 245162 167113
rect 245106 167039 245162 167048
rect 245016 136536 245068 136542
rect 245016 136478 245068 136484
rect 244924 132456 244976 132462
rect 244924 132398 244976 132404
rect 245014 131472 245070 131481
rect 245014 131407 245070 131416
rect 244924 128376 244976 128382
rect 244924 128318 244976 128324
rect 243912 123480 243964 123486
rect 243912 123422 243964 123428
rect 243818 123176 243874 123185
rect 243818 123111 243874 123120
rect 243832 82113 243860 123111
rect 243818 82104 243874 82113
rect 243818 82039 243874 82048
rect 243726 80880 243782 80889
rect 243726 80815 243782 80824
rect 244936 44849 244964 128318
rect 245028 55865 245056 131407
rect 245120 129033 245148 167039
rect 245292 160744 245344 160750
rect 245292 160686 245344 160692
rect 245200 131164 245252 131170
rect 245200 131106 245252 131112
rect 245106 129024 245162 129033
rect 245106 128959 245162 128968
rect 245106 102232 245162 102241
rect 245106 102167 245162 102176
rect 245014 55856 245070 55865
rect 245014 55791 245070 55800
rect 244922 44840 244978 44849
rect 244922 44775 244978 44784
rect 244278 33824 244334 33833
rect 244278 33759 244334 33768
rect 243544 32496 243596 32502
rect 243544 32438 243596 32444
rect 244292 16574 244320 33759
rect 245120 31074 245148 102167
rect 245212 94489 245240 131106
rect 245304 126954 245332 160686
rect 245672 141681 245700 214610
rect 245764 212430 245792 248639
rect 245856 223009 245884 263055
rect 246684 262886 246712 269039
rect 247052 263242 247080 284310
rect 247144 263362 247172 290119
rect 247236 267734 247264 292703
rect 247328 283626 247356 336738
rect 248420 284436 248472 284442
rect 248420 284378 248472 284384
rect 247316 283620 247368 283626
rect 247316 283562 247368 283568
rect 247236 267706 247356 267734
rect 247132 263356 247184 263362
rect 247132 263298 247184 263304
rect 247052 263214 247264 263242
rect 247040 263152 247092 263158
rect 247040 263094 247092 263100
rect 246672 262880 246724 262886
rect 246672 262822 246724 262828
rect 245934 262304 245990 262313
rect 245934 262239 245936 262248
rect 245988 262239 245990 262248
rect 245936 262210 245988 262216
rect 246396 261520 246448 261526
rect 246396 261462 246448 261468
rect 246408 260953 246436 261462
rect 246394 260944 246450 260953
rect 246394 260879 246450 260888
rect 245936 260228 245988 260234
rect 245936 260170 245988 260176
rect 245948 260137 245976 260170
rect 245934 260128 245990 260137
rect 245934 260063 245990 260072
rect 245936 259412 245988 259418
rect 245936 259354 245988 259360
rect 245948 258233 245976 259354
rect 245934 258224 245990 258233
rect 245934 258159 245990 258168
rect 246946 256048 247002 256057
rect 247052 256034 247080 263094
rect 247236 258074 247264 263214
rect 247328 261526 247356 267706
rect 247316 261520 247368 261526
rect 247316 261462 247368 261468
rect 247144 258046 247264 258074
rect 247144 257417 247172 258046
rect 247130 257408 247186 257417
rect 247130 257343 247186 257352
rect 247002 256006 247080 256034
rect 247144 256018 247172 257343
rect 247132 256012 247184 256018
rect 246946 255983 247002 255992
rect 247132 255954 247184 255960
rect 246946 255232 247002 255241
rect 247002 255190 247080 255218
rect 246946 255167 247002 255176
rect 245936 253904 245988 253910
rect 245934 253872 245936 253881
rect 245988 253872 245990 253881
rect 245934 253807 245990 253816
rect 246028 252544 246080 252550
rect 246028 252486 246080 252492
rect 245936 252476 245988 252482
rect 245936 252418 245988 252424
rect 245948 252249 245976 252418
rect 245934 252240 245990 252249
rect 245934 252175 245990 252184
rect 246040 251705 246068 252486
rect 246026 251696 246082 251705
rect 246026 251631 246082 251640
rect 245934 248160 245990 248169
rect 245934 248095 245990 248104
rect 245948 247722 245976 248095
rect 245936 247716 245988 247722
rect 245936 247658 245988 247664
rect 245936 246424 245988 246430
rect 245936 246366 245988 246372
rect 245948 245993 245976 246366
rect 245934 245984 245990 245993
rect 245934 245919 245990 245928
rect 245934 243808 245990 243817
rect 245934 243743 245990 243752
rect 245948 242962 245976 243743
rect 245936 242956 245988 242962
rect 245936 242898 245988 242904
rect 246394 242448 246450 242457
rect 246394 242383 246450 242392
rect 246408 241534 246436 242383
rect 246396 241528 246448 241534
rect 246396 241470 246448 241476
rect 245842 223000 245898 223009
rect 245842 222935 245898 222944
rect 247052 222154 247080 255190
rect 247130 244624 247186 244633
rect 247130 244559 247186 244568
rect 247040 222148 247092 222154
rect 247040 222090 247092 222096
rect 245752 212424 245804 212430
rect 245752 212366 245804 212372
rect 245764 183802 245792 212366
rect 246304 211200 246356 211206
rect 246304 211142 246356 211148
rect 245752 183796 245804 183802
rect 245752 183738 245804 183744
rect 245752 181484 245804 181490
rect 245752 181426 245804 181432
rect 245658 141672 245714 141681
rect 245658 141607 245714 141616
rect 245764 140758 245792 181426
rect 245842 179480 245898 179489
rect 245842 179415 245898 179424
rect 245856 158001 245884 179415
rect 246316 175982 246344 211142
rect 246304 175976 246356 175982
rect 246304 175918 246356 175924
rect 245842 157992 245898 158001
rect 245842 157927 245898 157936
rect 245752 140752 245804 140758
rect 245752 140694 245804 140700
rect 245292 126948 245344 126954
rect 245292 126890 245344 126896
rect 246316 98666 246344 175918
rect 247052 169046 247080 222090
rect 247144 208350 247172 244559
rect 247224 241528 247276 241534
rect 247224 241470 247276 241476
rect 247236 237386 247264 241470
rect 247224 237380 247276 237386
rect 247224 237322 247276 237328
rect 247132 208344 247184 208350
rect 247132 208286 247184 208292
rect 247040 169040 247092 169046
rect 247040 168982 247092 168988
rect 247144 167249 247172 208286
rect 247222 175944 247278 175953
rect 247222 175879 247278 175888
rect 247130 167240 247186 167249
rect 247130 167175 247186 167184
rect 246580 154692 246632 154698
rect 246580 154634 246632 154640
rect 246394 139768 246450 139777
rect 246394 139703 246450 139712
rect 246408 108322 246436 139703
rect 246486 127392 246542 127401
rect 246486 127327 246542 127336
rect 246396 108316 246448 108322
rect 246396 108258 246448 108264
rect 246396 100768 246448 100774
rect 246396 100710 246448 100716
rect 246304 98660 246356 98666
rect 246304 98602 246356 98608
rect 245198 94480 245254 94489
rect 245198 94415 245254 94424
rect 246408 47569 246436 100710
rect 246500 87553 246528 127327
rect 246592 126274 246620 154634
rect 247236 149054 247264 175879
rect 248432 171834 248460 284378
rect 248524 280838 248552 372574
rect 306748 368552 306800 368558
rect 306748 368494 306800 368500
rect 305000 365764 305052 365770
rect 305000 365706 305052 365712
rect 259458 360904 259514 360913
rect 259458 360839 259514 360848
rect 252558 353424 252614 353433
rect 252558 353359 252614 353368
rect 251180 342304 251232 342310
rect 251180 342246 251232 342252
rect 249984 338156 250036 338162
rect 249984 338098 250036 338104
rect 248604 327820 248656 327826
rect 248604 327762 248656 327768
rect 248616 283801 248644 327762
rect 249890 307864 249946 307873
rect 249890 307799 249946 307808
rect 248696 294024 248748 294030
rect 248696 293966 248748 293972
rect 248602 283792 248658 283801
rect 248602 283727 248658 283736
rect 248512 280832 248564 280838
rect 248512 280774 248564 280780
rect 248604 271516 248656 271522
rect 248604 271458 248656 271464
rect 248510 261760 248566 261769
rect 248510 261695 248566 261704
rect 248524 223582 248552 261695
rect 248616 236609 248644 271458
rect 248708 260234 248736 293966
rect 249798 287464 249854 287473
rect 249798 287399 249854 287408
rect 248696 260228 248748 260234
rect 248696 260170 248748 260176
rect 248696 247716 248748 247722
rect 248696 247658 248748 247664
rect 248602 236600 248658 236609
rect 248602 236535 248658 236544
rect 248512 223576 248564 223582
rect 248512 223518 248564 223524
rect 248420 171828 248472 171834
rect 248420 171770 248472 171776
rect 247776 168496 247828 168502
rect 247776 168438 247828 168444
rect 247224 149048 247276 149054
rect 247224 148990 247276 148996
rect 247682 135416 247738 135425
rect 247682 135351 247738 135360
rect 246580 126268 246632 126274
rect 246580 126210 246632 126216
rect 246580 98048 246632 98054
rect 246580 97990 246632 97996
rect 246486 87544 246542 87553
rect 246486 87479 246542 87488
rect 246592 76537 246620 97990
rect 246578 76528 246634 76537
rect 246578 76463 246634 76472
rect 247696 61577 247724 135351
rect 247788 129742 247816 168438
rect 248052 167136 248104 167142
rect 248052 167078 248104 167084
rect 247960 146328 248012 146334
rect 247960 146270 248012 146276
rect 247776 129736 247828 129742
rect 247776 129678 247828 129684
rect 247868 127628 247920 127634
rect 247868 127570 247920 127576
rect 247776 110492 247828 110498
rect 247776 110434 247828 110440
rect 247682 61568 247738 61577
rect 247682 61503 247738 61512
rect 247788 49094 247816 110434
rect 247880 82142 247908 127570
rect 247972 106214 248000 146270
rect 248064 128246 248092 167078
rect 248524 164898 248552 223518
rect 248708 220833 248736 247658
rect 248694 220824 248750 220833
rect 248694 220759 248750 220768
rect 249064 212832 249116 212838
rect 249064 212774 249116 212780
rect 248512 164892 248564 164898
rect 248512 164834 248564 164840
rect 249076 144226 249104 212774
rect 249154 174040 249210 174049
rect 249154 173975 249210 173984
rect 249064 144220 249116 144226
rect 249064 144162 249116 144168
rect 249168 135182 249196 173975
rect 249812 157185 249840 287399
rect 249904 279886 249932 307799
rect 249892 279880 249944 279886
rect 249892 279822 249944 279828
rect 249892 273284 249944 273290
rect 249892 273226 249944 273232
rect 249904 196042 249932 273226
rect 249996 265810 250024 338098
rect 250076 281716 250128 281722
rect 250076 281658 250128 281664
rect 249984 265804 250036 265810
rect 249984 265746 250036 265752
rect 249996 265713 250024 265746
rect 249982 265704 250038 265713
rect 249982 265639 250038 265648
rect 250088 229094 250116 281658
rect 251088 279880 251140 279886
rect 251088 279822 251140 279828
rect 251100 279478 251128 279822
rect 251088 279472 251140 279478
rect 251088 279414 251140 279420
rect 251192 270502 251220 342246
rect 251364 330608 251416 330614
rect 251364 330550 251416 330556
rect 251270 296984 251326 296993
rect 251270 296919 251326 296928
rect 251180 270496 251232 270502
rect 251180 270438 251232 270444
rect 251180 261520 251232 261526
rect 251180 261462 251232 261468
rect 249996 229066 250116 229094
rect 249996 227730 250024 229066
rect 249984 227724 250036 227730
rect 249984 227666 250036 227672
rect 249892 196036 249944 196042
rect 249892 195978 249944 195984
rect 249904 175234 249932 195978
rect 249892 175228 249944 175234
rect 249892 175170 249944 175176
rect 249996 162081 250024 227666
rect 250536 172644 250588 172650
rect 250536 172586 250588 172592
rect 249982 162072 250038 162081
rect 249982 162007 250038 162016
rect 249798 157176 249854 157185
rect 249798 157111 249854 157120
rect 250442 156496 250498 156505
rect 250442 156431 250498 156440
rect 249248 149728 249300 149734
rect 249248 149670 249300 149676
rect 249156 135176 249208 135182
rect 249156 135118 249208 135124
rect 248052 128240 248104 128246
rect 248052 128182 248104 128188
rect 249156 125656 249208 125662
rect 249156 125598 249208 125604
rect 249168 117978 249196 125598
rect 249156 117972 249208 117978
rect 249156 117914 249208 117920
rect 249064 117360 249116 117366
rect 249064 117302 249116 117308
rect 247960 106208 248012 106214
rect 247960 106150 248012 106156
rect 247868 82136 247920 82142
rect 247868 82078 247920 82084
rect 247776 49088 247828 49094
rect 247776 49030 247828 49036
rect 246394 47560 246450 47569
rect 246394 47495 246450 47504
rect 249076 42158 249104 117302
rect 249156 114572 249208 114578
rect 249156 114514 249208 114520
rect 249168 66881 249196 114514
rect 249260 113082 249288 149670
rect 249338 142488 249394 142497
rect 249338 142423 249394 142432
rect 249248 113076 249300 113082
rect 249248 113018 249300 113024
rect 249246 109848 249302 109857
rect 249246 109783 249302 109792
rect 249260 83570 249288 109783
rect 249352 109750 249380 142423
rect 250456 115841 250484 156431
rect 250548 133890 250576 172586
rect 250628 162988 250680 162994
rect 250628 162930 250680 162936
rect 250536 133884 250588 133890
rect 250536 133826 250588 133832
rect 250640 124914 250668 162930
rect 251192 144809 251220 261462
rect 251284 212838 251312 296919
rect 251376 252482 251404 330550
rect 251824 285796 251876 285802
rect 251824 285738 251876 285744
rect 251456 262268 251508 262274
rect 251456 262210 251508 262216
rect 251364 252476 251416 252482
rect 251364 252418 251416 252424
rect 251272 212832 251324 212838
rect 251272 212774 251324 212780
rect 251272 210520 251324 210526
rect 251272 210462 251324 210468
rect 251284 151162 251312 210462
rect 251468 202842 251496 262210
rect 251836 261526 251864 285738
rect 252572 282878 252600 353359
rect 255412 347812 255464 347818
rect 255412 347754 255464 347760
rect 252652 321020 252704 321026
rect 252652 320962 252704 320968
rect 252560 282872 252612 282878
rect 252560 282814 252612 282820
rect 252664 272542 252692 320962
rect 253938 303648 253994 303657
rect 253938 303583 253994 303592
rect 252744 298240 252796 298246
rect 252744 298182 252796 298188
rect 252652 272536 252704 272542
rect 252652 272478 252704 272484
rect 252652 270496 252704 270502
rect 252652 270438 252704 270444
rect 251824 261520 251876 261526
rect 251824 261462 251876 261468
rect 251456 202836 251508 202842
rect 251456 202778 251508 202784
rect 251468 200114 251496 202778
rect 251376 200086 251496 200114
rect 251376 173233 251404 200086
rect 252664 180130 252692 270438
rect 252756 250510 252784 298182
rect 252836 283620 252888 283626
rect 252836 283562 252888 283568
rect 252744 250504 252796 250510
rect 252744 250446 252796 250452
rect 252652 180124 252704 180130
rect 252652 180066 252704 180072
rect 251362 173224 251418 173233
rect 251362 173159 251418 173168
rect 251824 164280 251876 164286
rect 251824 164222 251876 164228
rect 251272 151156 251324 151162
rect 251272 151098 251324 151104
rect 251178 144800 251234 144809
rect 251178 144735 251234 144744
rect 250812 143676 250864 143682
rect 250812 143618 250864 143624
rect 250628 124908 250680 124914
rect 250628 124850 250680 124856
rect 250720 123480 250772 123486
rect 250720 123422 250772 123428
rect 250442 115832 250498 115841
rect 250442 115767 250498 115776
rect 250442 113248 250498 113257
rect 250442 113183 250498 113192
rect 249340 109744 249392 109750
rect 249340 109686 249392 109692
rect 249248 83564 249300 83570
rect 249248 83506 249300 83512
rect 249154 66872 249210 66881
rect 249154 66807 249210 66816
rect 249064 42152 249116 42158
rect 249064 42094 249116 42100
rect 248420 36644 248472 36650
rect 248420 36586 248472 36592
rect 245108 31068 245160 31074
rect 245108 31010 245160 31016
rect 241532 16546 241744 16574
rect 244292 16546 245240 16574
rect 240784 4820 240836 4826
rect 240784 4762 240836 4768
rect 240336 598 240548 626
rect 240336 490 240364 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 462 240364 490
rect 240520 480 240548 598
rect 241716 480 241744 16546
rect 244094 10296 244150 10305
rect 244094 10231 244150 10240
rect 242898 4992 242954 5001
rect 242898 4927 242954 4936
rect 242912 480 242940 4927
rect 244108 480 244136 10231
rect 245212 480 245240 16546
rect 247590 3496 247646 3505
rect 247590 3431 247646 3440
rect 246394 3360 246450 3369
rect 246394 3295 246450 3304
rect 246408 480 246436 3295
rect 247604 480 247632 3431
rect 248432 490 248460 36586
rect 249800 32428 249852 32434
rect 249800 32370 249852 32376
rect 249812 16574 249840 32370
rect 250456 17338 250484 113183
rect 250626 112024 250682 112033
rect 250626 111959 250682 111968
rect 250536 107704 250588 107710
rect 250536 107646 250588 107652
rect 250548 55894 250576 107646
rect 250640 71058 250668 111959
rect 250732 87650 250760 123422
rect 250824 111110 250852 143618
rect 251836 124137 251864 164222
rect 251914 157992 251970 158001
rect 251914 157927 251970 157936
rect 251822 124128 251878 124137
rect 251822 124063 251878 124072
rect 251928 118658 251956 157927
rect 252098 144120 252154 144129
rect 252098 144055 252154 144064
rect 252008 124296 252060 124302
rect 252008 124238 252060 124244
rect 251916 118652 251968 118658
rect 251916 118594 251968 118600
rect 250812 111104 250864 111110
rect 250812 111046 250864 111052
rect 251824 109132 251876 109138
rect 251824 109074 251876 109080
rect 250720 87644 250772 87650
rect 250720 87586 250772 87592
rect 250628 71052 250680 71058
rect 250628 70994 250680 71000
rect 250536 55888 250588 55894
rect 250536 55830 250588 55836
rect 250444 17332 250496 17338
rect 250444 17274 250496 17280
rect 249812 16546 250024 16574
rect 248616 598 248828 626
rect 248616 490 248644 598
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 462 248644 490
rect 248800 480 248828 598
rect 249996 480 250024 16546
rect 251180 11756 251232 11762
rect 251180 11698 251232 11704
rect 251192 480 251220 11698
rect 251836 10334 251864 109074
rect 251914 107944 251970 107953
rect 251914 107879 251970 107888
rect 251928 44878 251956 107879
rect 252020 73846 252048 124238
rect 252112 109041 252140 144055
rect 252848 143041 252876 283562
rect 253952 276010 253980 303583
rect 254030 292904 254086 292913
rect 254030 292839 254086 292848
rect 253940 276004 253992 276010
rect 253940 275946 253992 275952
rect 253848 272536 253900 272542
rect 253848 272478 253900 272484
rect 253860 271810 253888 272478
rect 253860 271782 253980 271810
rect 253020 250504 253072 250510
rect 253020 250446 253072 250452
rect 253032 249082 253060 250446
rect 253020 249076 253072 249082
rect 253020 249018 253072 249024
rect 253294 168464 253350 168473
rect 253294 168399 253350 168408
rect 253202 160440 253258 160449
rect 253202 160375 253258 160384
rect 252834 143032 252890 143041
rect 252834 142967 252890 142976
rect 253216 120057 253244 160375
rect 253308 128314 253336 168399
rect 253952 160041 253980 271782
rect 254044 246430 254072 292839
rect 255320 292596 255372 292602
rect 255320 292538 255372 292544
rect 254122 291272 254178 291281
rect 254122 291207 254178 291216
rect 254136 278730 254164 291207
rect 254124 278724 254176 278730
rect 254124 278666 254176 278672
rect 254136 278050 254164 278666
rect 254124 278044 254176 278050
rect 254124 277986 254176 277992
rect 254032 246424 254084 246430
rect 254032 246366 254084 246372
rect 254044 245682 254072 246366
rect 254032 245676 254084 245682
rect 254032 245618 254084 245624
rect 254584 245676 254636 245682
rect 254584 245618 254636 245624
rect 254596 217326 254624 245618
rect 254032 217320 254084 217326
rect 254032 217262 254084 217268
rect 254584 217320 254636 217326
rect 254584 217262 254636 217268
rect 253938 160032 253994 160041
rect 253938 159967 253994 159976
rect 254044 137970 254072 217262
rect 255332 168609 255360 292538
rect 255424 238377 255452 347754
rect 258172 340944 258224 340950
rect 258172 340886 258224 340892
rect 255504 324964 255556 324970
rect 255504 324906 255556 324912
rect 255516 254153 255544 324906
rect 258080 318844 258132 318850
rect 258080 318786 258132 318792
rect 256698 316160 256754 316169
rect 256698 316095 256754 316104
rect 255502 254144 255558 254153
rect 255502 254079 255558 254088
rect 255410 238368 255466 238377
rect 255410 238303 255466 238312
rect 255424 237969 255452 238303
rect 255410 237960 255466 237969
rect 255410 237895 255466 237904
rect 256146 174312 256202 174321
rect 256146 174247 256202 174256
rect 255318 168600 255374 168609
rect 255318 168535 255374 168544
rect 255962 161800 256018 161809
rect 255962 161735 256018 161744
rect 254584 161492 254636 161498
rect 254584 161434 254636 161440
rect 254032 137964 254084 137970
rect 254032 137906 254084 137912
rect 253388 129804 253440 129810
rect 253388 129746 253440 129752
rect 253296 128308 253348 128314
rect 253296 128250 253348 128256
rect 253296 125724 253348 125730
rect 253296 125666 253348 125672
rect 253202 120048 253258 120057
rect 253202 119983 253258 119992
rect 252098 109032 252154 109041
rect 252098 108967 252154 108976
rect 252100 106344 252152 106350
rect 252100 106286 252152 106292
rect 252008 73840 252060 73846
rect 252008 73782 252060 73788
rect 252112 58682 252140 106286
rect 253202 92576 253258 92585
rect 253202 92511 253258 92520
rect 252100 58676 252152 58682
rect 252100 58618 252152 58624
rect 251916 44872 251968 44878
rect 251916 44814 251968 44820
rect 253216 35222 253244 92511
rect 253308 83473 253336 125666
rect 253400 109721 253428 129746
rect 254596 122738 254624 161434
rect 254768 142248 254820 142254
rect 254768 142190 254820 142196
rect 254584 122732 254636 122738
rect 254584 122674 254636 122680
rect 253480 121508 253532 121514
rect 253480 121450 253532 121456
rect 253386 109712 253442 109721
rect 253386 109647 253442 109656
rect 253388 98116 253440 98122
rect 253388 98058 253440 98064
rect 253294 83464 253350 83473
rect 253294 83399 253350 83408
rect 253400 64161 253428 98058
rect 253492 94518 253520 121450
rect 254584 117428 254636 117434
rect 254584 117370 254636 117376
rect 253572 104916 253624 104922
rect 253572 104858 253624 104864
rect 253480 94512 253532 94518
rect 253480 94454 253532 94460
rect 253584 91798 253612 104858
rect 253572 91792 253624 91798
rect 253572 91734 253624 91740
rect 253386 64152 253442 64161
rect 253386 64087 253442 64096
rect 254596 39370 254624 117370
rect 254674 110392 254730 110401
rect 254674 110327 254730 110336
rect 254688 68338 254716 110327
rect 254780 102134 254808 142190
rect 254858 129976 254914 129985
rect 254858 129911 254914 129920
rect 254768 102128 254820 102134
rect 254768 102070 254820 102076
rect 254872 92585 254900 129911
rect 255976 121446 256004 161735
rect 256056 149116 256108 149122
rect 256056 149058 256108 149064
rect 255964 121440 256016 121446
rect 255964 121382 256016 121388
rect 255964 118720 256016 118726
rect 255964 118662 256016 118668
rect 254858 92576 254914 92585
rect 254858 92511 254914 92520
rect 255976 76673 256004 118662
rect 256068 109002 256096 149058
rect 256160 135250 256188 174247
rect 256712 136610 256740 316095
rect 256882 298208 256938 298217
rect 256882 298143 256938 298152
rect 256792 291236 256844 291242
rect 256792 291178 256844 291184
rect 256804 253230 256832 291178
rect 256896 270502 256924 298143
rect 256884 270496 256936 270502
rect 256884 270438 256936 270444
rect 256896 269822 256924 270438
rect 256884 269816 256936 269822
rect 256884 269758 256936 269764
rect 256792 253224 256844 253230
rect 256792 253166 256844 253172
rect 256804 250510 256832 253166
rect 256792 250504 256844 250510
rect 256792 250446 256844 250452
rect 257436 238808 257488 238814
rect 257436 238750 257488 238756
rect 257342 209128 257398 209137
rect 257342 209063 257398 209072
rect 256700 136604 256752 136610
rect 256700 136546 256752 136552
rect 256240 135312 256292 135318
rect 256240 135254 256292 135260
rect 256148 135244 256200 135250
rect 256148 135186 256200 135192
rect 256056 108996 256108 109002
rect 256056 108938 256108 108944
rect 256054 106312 256110 106321
rect 256054 106247 256110 106256
rect 255962 76664 256018 76673
rect 255962 76599 256018 76608
rect 256068 73953 256096 106247
rect 256252 105505 256280 135254
rect 256330 107808 256386 107817
rect 256330 107743 256386 107752
rect 256238 105496 256294 105505
rect 256238 105431 256294 105440
rect 256344 102814 256372 107743
rect 256332 102808 256384 102814
rect 256332 102750 256384 102756
rect 256148 102196 256200 102202
rect 256148 102138 256200 102144
rect 256160 90370 256188 102138
rect 256148 90364 256200 90370
rect 256148 90306 256200 90312
rect 256054 73944 256110 73953
rect 256054 73879 256110 73888
rect 255318 71088 255374 71097
rect 255318 71023 255374 71032
rect 254676 68332 254728 68338
rect 254676 68274 254728 68280
rect 254584 39364 254636 39370
rect 254584 39306 254636 39312
rect 253204 35216 253256 35222
rect 253204 35158 253256 35164
rect 255332 16574 255360 71023
rect 255332 16546 255912 16574
rect 253480 15972 253532 15978
rect 253480 15914 253532 15920
rect 251824 10328 251876 10334
rect 251824 10270 251876 10276
rect 252374 3496 252430 3505
rect 252374 3431 252430 3440
rect 252388 480 252416 3431
rect 253492 480 253520 15914
rect 254674 2000 254730 2009
rect 254674 1935 254730 1944
rect 254688 480 254716 1935
rect 255884 480 255912 16546
rect 257068 3528 257120 3534
rect 257068 3470 257120 3476
rect 257080 480 257108 3470
rect 257356 3466 257384 209063
rect 257448 180130 257476 238750
rect 257436 180124 257488 180130
rect 257436 180066 257488 180072
rect 258092 166326 258120 318786
rect 258184 238746 258212 340886
rect 258356 325032 258408 325038
rect 258356 324974 258408 324980
rect 258264 299600 258316 299606
rect 258264 299542 258316 299548
rect 258276 253910 258304 299542
rect 258368 281518 258396 324974
rect 258356 281512 258408 281518
rect 258356 281454 258408 281460
rect 259368 281512 259420 281518
rect 259368 281454 259420 281460
rect 259380 280906 259408 281454
rect 259368 280900 259420 280906
rect 259368 280842 259420 280848
rect 258264 253904 258316 253910
rect 258264 253846 258316 253852
rect 259368 253904 259420 253910
rect 259368 253846 259420 253852
rect 259380 253230 259408 253846
rect 259368 253224 259420 253230
rect 259368 253166 259420 253172
rect 259472 252550 259500 360839
rect 262218 358864 262274 358873
rect 262218 358799 262274 358808
rect 260840 309188 260892 309194
rect 260840 309130 260892 309136
rect 260102 301064 260158 301073
rect 260102 300999 260158 301008
rect 259552 295384 259604 295390
rect 259552 295326 259604 295332
rect 259564 259418 259592 295326
rect 259552 259412 259604 259418
rect 259552 259354 259604 259360
rect 259460 252544 259512 252550
rect 259460 252486 259512 252492
rect 258172 238740 258224 238746
rect 258172 238682 258224 238688
rect 258816 171284 258868 171290
rect 258816 171226 258868 171232
rect 258080 166320 258132 166326
rect 258080 166262 258132 166268
rect 257620 164348 257672 164354
rect 257620 164290 257672 164296
rect 257528 136740 257580 136746
rect 257528 136682 257580 136688
rect 257436 133952 257488 133958
rect 257436 133894 257488 133900
rect 257448 64297 257476 133894
rect 257540 100065 257568 136682
rect 257632 130393 257660 164290
rect 258722 160304 258778 160313
rect 258722 160239 258778 160248
rect 257618 130384 257674 130393
rect 257618 130319 257674 130328
rect 258736 120086 258764 160239
rect 258828 140049 258856 171226
rect 259092 147688 259144 147694
rect 259092 147630 259144 147636
rect 258814 140040 258870 140049
rect 258814 139975 258870 139984
rect 259000 139528 259052 139534
rect 259000 139470 259052 139476
rect 258814 123040 258870 123049
rect 258814 122975 258870 122984
rect 258724 120080 258776 120086
rect 258724 120022 258776 120028
rect 258078 114744 258134 114753
rect 258078 114679 258134 114688
rect 258092 110401 258120 114679
rect 258078 110392 258134 110401
rect 258078 110327 258134 110336
rect 258724 107772 258776 107778
rect 258724 107714 258776 107720
rect 257526 100056 257582 100065
rect 257526 99991 257582 100000
rect 257620 99408 257672 99414
rect 257620 99350 257672 99356
rect 257632 89010 257660 99350
rect 257620 89004 257672 89010
rect 257620 88946 257672 88952
rect 257434 64288 257490 64297
rect 257434 64223 257490 64232
rect 258080 28348 258132 28354
rect 258080 28290 258132 28296
rect 258092 16574 258120 28290
rect 258736 26926 258764 107714
rect 258828 75313 258856 122975
rect 258908 106412 258960 106418
rect 258908 106354 258960 106360
rect 258814 75304 258870 75313
rect 258814 75239 258870 75248
rect 258920 60042 258948 106354
rect 259012 97986 259040 139470
rect 259104 107642 259132 147630
rect 259092 107636 259144 107642
rect 259092 107578 259144 107584
rect 259000 97980 259052 97986
rect 259000 97922 259052 97928
rect 259092 96688 259144 96694
rect 259092 96630 259144 96636
rect 259104 80753 259132 96630
rect 260116 95198 260144 300999
rect 260748 259412 260800 259418
rect 260748 259354 260800 259360
rect 260760 258738 260788 259354
rect 260748 258732 260800 258738
rect 260748 258674 260800 258680
rect 260196 257372 260248 257378
rect 260196 257314 260248 257320
rect 260208 237289 260236 257314
rect 260852 256086 260880 309130
rect 260840 256080 260892 256086
rect 260840 256022 260892 256028
rect 260852 254590 260880 256022
rect 260840 254584 260892 254590
rect 260840 254526 260892 254532
rect 260748 252544 260800 252550
rect 260748 252486 260800 252492
rect 260760 251870 260788 252486
rect 260748 251864 260800 251870
rect 260748 251806 260800 251812
rect 262232 240145 262260 358799
rect 263598 351928 263654 351937
rect 263598 351863 263654 351872
rect 262862 302288 262918 302297
rect 262862 302223 262918 302232
rect 262218 240136 262274 240145
rect 262218 240071 262274 240080
rect 260194 237280 260250 237289
rect 260194 237215 260250 237224
rect 262876 181529 262904 302223
rect 263612 269074 263640 351863
rect 267738 346488 267794 346497
rect 267738 346423 267794 346432
rect 267002 310584 267058 310593
rect 267002 310519 267058 310528
rect 265624 309256 265676 309262
rect 265624 309198 265676 309204
rect 264244 289876 264296 289882
rect 264244 289818 264296 289824
rect 263600 269068 263652 269074
rect 263600 269010 263652 269016
rect 263612 268394 263640 269010
rect 263600 268388 263652 268394
rect 263600 268330 263652 268336
rect 262862 181520 262918 181529
rect 262862 181455 262918 181464
rect 263140 174004 263192 174010
rect 263140 173946 263192 173952
rect 260286 170232 260342 170241
rect 260286 170167 260342 170176
rect 260194 151328 260250 151337
rect 260194 151263 260250 151272
rect 260208 111081 260236 151263
rect 260300 131102 260328 170167
rect 262864 165708 262916 165714
rect 262864 165650 262916 165656
rect 262876 160750 262904 165650
rect 262864 160744 262916 160750
rect 262864 160686 262916 160692
rect 262956 153264 263008 153270
rect 262956 153206 263008 153212
rect 261484 150476 261536 150482
rect 261484 150418 261536 150424
rect 260288 131096 260340 131102
rect 260288 131038 260340 131044
rect 260288 120148 260340 120154
rect 260288 120090 260340 120096
rect 260194 111072 260250 111081
rect 260194 111007 260250 111016
rect 260194 105224 260250 105233
rect 260194 105159 260250 105168
rect 260104 95192 260156 95198
rect 260104 95134 260156 95140
rect 259090 80744 259146 80753
rect 259090 80679 259146 80688
rect 258908 60036 258960 60042
rect 258908 59978 258960 59984
rect 260208 38010 260236 105159
rect 260300 77897 260328 120090
rect 261496 113801 261524 150418
rect 262862 147792 262918 147801
rect 262862 147727 262918 147736
rect 261760 134020 261812 134026
rect 261760 133962 261812 133968
rect 261576 128444 261628 128450
rect 261576 128386 261628 128392
rect 261482 113792 261538 113801
rect 261482 113727 261538 113736
rect 260380 111852 260432 111858
rect 260380 111794 260432 111800
rect 260392 87718 260420 111794
rect 261484 110560 261536 110566
rect 261484 110502 261536 110508
rect 260380 87712 260432 87718
rect 260380 87654 260432 87660
rect 260286 77888 260342 77897
rect 260286 77823 260342 77832
rect 260196 38004 260248 38010
rect 260196 37946 260248 37952
rect 261496 35290 261524 110502
rect 261588 62801 261616 128386
rect 261668 113620 261720 113626
rect 261668 113562 261720 113568
rect 261680 69601 261708 113562
rect 261772 109857 261800 133962
rect 262770 133240 262826 133249
rect 262770 133175 262826 133184
rect 262784 132841 262812 133175
rect 262770 132832 262826 132841
rect 262770 132767 262826 132776
rect 262770 127664 262826 127673
rect 262770 127599 262826 127608
rect 262784 127265 262812 127599
rect 262770 127256 262826 127265
rect 262770 127191 262826 127200
rect 261758 109848 261814 109857
rect 261758 109783 261814 109792
rect 262876 106282 262904 147727
rect 262968 113150 262996 153206
rect 263152 141438 263180 173946
rect 263230 161528 263286 161537
rect 263230 161463 263286 161472
rect 263140 141432 263192 141438
rect 263140 141374 263192 141380
rect 263048 140888 263100 140894
rect 263048 140830 263100 140836
rect 262956 113144 263008 113150
rect 262956 113086 263008 113092
rect 262864 106276 262916 106282
rect 262864 106218 262916 106224
rect 262956 104984 263008 104990
rect 262956 104926 263008 104932
rect 262772 102264 262824 102270
rect 262772 102206 262824 102212
rect 262784 93854 262812 102206
rect 262862 99648 262918 99657
rect 262862 99583 262918 99592
rect 262876 95985 262904 99583
rect 262862 95976 262918 95985
rect 262862 95911 262918 95920
rect 262784 93826 262904 93854
rect 262218 69728 262274 69737
rect 262218 69663 262274 69672
rect 261666 69592 261722 69601
rect 261666 69527 261722 69536
rect 261574 62792 261630 62801
rect 261574 62727 261630 62736
rect 261484 35284 261536 35290
rect 261484 35226 261536 35232
rect 258724 26920 258776 26926
rect 258724 26862 258776 26868
rect 259458 21312 259514 21321
rect 259458 21247 259514 21256
rect 258092 16546 258304 16574
rect 257344 3460 257396 3466
rect 257344 3402 257396 3408
rect 258276 480 258304 16546
rect 259472 480 259500 21247
rect 262232 16574 262260 69663
rect 262876 46238 262904 93826
rect 262968 61441 262996 104926
rect 263060 100706 263088 140830
rect 263244 140078 263272 161463
rect 263232 140072 263284 140078
rect 263232 140014 263284 140020
rect 263140 139460 263192 139466
rect 263140 139402 263192 139408
rect 263152 123486 263180 139402
rect 264256 131646 264284 289818
rect 264336 288448 264388 288454
rect 264336 288390 264388 288396
rect 264348 274038 264376 288390
rect 264336 274032 264388 274038
rect 264336 273974 264388 273980
rect 265636 242282 265664 309198
rect 265624 242276 265676 242282
rect 265624 242218 265676 242224
rect 267016 189786 267044 310519
rect 267096 287156 267148 287162
rect 267096 287098 267148 287104
rect 267004 189780 267056 189786
rect 267004 189722 267056 189728
rect 267108 179489 267136 287098
rect 267752 266354 267780 346423
rect 302240 314696 302292 314702
rect 302240 314638 302292 314644
rect 286324 307896 286376 307902
rect 286324 307838 286376 307844
rect 280896 306468 280948 306474
rect 280896 306410 280948 306416
rect 271236 303748 271288 303754
rect 271236 303690 271288 303696
rect 269762 298344 269818 298353
rect 269762 298279 269818 298288
rect 267740 266348 267792 266354
rect 267740 266290 267792 266296
rect 269028 266348 269080 266354
rect 269028 266290 269080 266296
rect 269040 265674 269068 266290
rect 269028 265668 269080 265674
rect 269028 265610 269080 265616
rect 268384 241528 268436 241534
rect 268384 241470 268436 241476
rect 266358 179480 266414 179489
rect 266358 179415 266414 179424
rect 267094 179480 267150 179489
rect 267094 179415 267150 179424
rect 266372 177993 266400 179415
rect 266358 177984 266414 177993
rect 266358 177919 266414 177928
rect 268396 177342 268424 241470
rect 269776 185609 269804 298279
rect 269854 286104 269910 286113
rect 269854 286039 269910 286048
rect 269762 185600 269818 185609
rect 269762 185535 269818 185544
rect 269868 181490 269896 286039
rect 271144 280900 271196 280906
rect 271144 280842 271196 280848
rect 269856 181484 269908 181490
rect 269856 181426 269908 181432
rect 271156 177410 271184 280842
rect 271248 242214 271276 303690
rect 276664 300892 276716 300898
rect 276664 300834 276716 300840
rect 273904 280832 273956 280838
rect 273904 280774 273956 280780
rect 271328 242956 271380 242962
rect 271328 242898 271380 242904
rect 271236 242208 271288 242214
rect 271236 242150 271288 242156
rect 271340 182918 271368 242898
rect 272524 227044 272576 227050
rect 272524 226986 272576 226992
rect 271328 182912 271380 182918
rect 271328 182854 271380 182860
rect 272536 180198 272564 226986
rect 272524 180192 272576 180198
rect 272524 180134 272576 180140
rect 273916 178809 273944 280774
rect 276020 266416 276072 266422
rect 276020 266358 276072 266364
rect 276032 201385 276060 266358
rect 276676 227050 276704 300834
rect 278044 276684 278096 276690
rect 278044 276626 278096 276632
rect 276664 227044 276716 227050
rect 276664 226986 276716 226992
rect 276662 211848 276718 211857
rect 276662 211783 276718 211792
rect 276018 201376 276074 201385
rect 276018 201311 276074 201320
rect 274548 181552 274600 181558
rect 274548 181494 274600 181500
rect 274560 178945 274588 181494
rect 274546 178936 274602 178945
rect 274546 178871 274602 178880
rect 273902 178800 273958 178809
rect 273902 178735 273958 178744
rect 271144 177404 271196 177410
rect 271144 177346 271196 177352
rect 268384 177336 268436 177342
rect 268384 177278 268436 177284
rect 276676 176050 276704 211783
rect 276754 201376 276810 201385
rect 276754 201311 276810 201320
rect 276768 177449 276796 201311
rect 278056 178770 278084 276626
rect 280804 274032 280856 274038
rect 280804 273974 280856 273980
rect 278872 242276 278924 242282
rect 278872 242218 278924 242224
rect 278134 198112 278190 198121
rect 278134 198047 278190 198056
rect 278044 178764 278096 178770
rect 278044 178706 278096 178712
rect 276754 177440 276810 177449
rect 276754 177375 276810 177384
rect 278148 177313 278176 198047
rect 278134 177304 278190 177313
rect 278134 177239 278190 177248
rect 278884 177041 278912 242218
rect 279056 199504 279108 199510
rect 279056 199446 279108 199452
rect 278870 177032 278926 177041
rect 278870 176967 278926 176976
rect 276664 176044 276716 176050
rect 276664 175986 276716 175992
rect 278780 175976 278832 175982
rect 273350 175944 273406 175953
rect 273350 175879 273406 175888
rect 278778 175944 278780 175953
rect 278832 175944 278834 175953
rect 278778 175879 278834 175888
rect 273364 175846 273392 175879
rect 273352 175840 273404 175846
rect 273352 175782 273404 175788
rect 264978 175672 265034 175681
rect 264978 175607 265034 175616
rect 264992 175302 265020 175607
rect 264980 175296 265032 175302
rect 264980 175238 265032 175244
rect 265070 175264 265126 175273
rect 265070 175199 265126 175208
rect 264978 174856 265034 174865
rect 264978 174791 265034 174800
rect 264992 174010 265020 174791
rect 264980 174004 265032 174010
rect 264980 173946 265032 173952
rect 265084 173942 265112 175199
rect 265072 173936 265124 173942
rect 265072 173878 265124 173884
rect 265070 173632 265126 173641
rect 265070 173567 265126 173576
rect 264978 172680 265034 172689
rect 264978 172615 264980 172624
rect 265032 172615 265034 172624
rect 264980 172586 265032 172592
rect 265084 172582 265112 173567
rect 265072 172576 265124 172582
rect 265072 172518 265124 172524
rect 265070 172272 265126 172281
rect 265070 172207 265126 172216
rect 264978 171456 265034 171465
rect 264978 171391 265034 171400
rect 264992 171290 265020 171391
rect 264980 171284 265032 171290
rect 264980 171226 265032 171232
rect 265084 171154 265112 172207
rect 265072 171148 265124 171154
rect 265072 171090 265124 171096
rect 265070 171048 265126 171057
rect 265070 170983 265126 170992
rect 264978 170096 265034 170105
rect 264978 170031 265034 170040
rect 264992 169862 265020 170031
rect 264980 169856 265032 169862
rect 264980 169798 265032 169804
rect 265084 169794 265112 170983
rect 265072 169788 265124 169794
rect 265072 169730 265124 169736
rect 265070 169688 265126 169697
rect 265070 169623 265126 169632
rect 264978 169280 265034 169289
rect 264978 169215 265034 169224
rect 264992 168502 265020 169215
rect 264980 168496 265032 168502
rect 264980 168438 265032 168444
rect 265084 168434 265112 169623
rect 265162 168872 265218 168881
rect 265162 168807 265218 168816
rect 265072 168428 265124 168434
rect 265072 168370 265124 168376
rect 264978 167920 265034 167929
rect 264978 167855 265034 167864
rect 264992 167142 265020 167855
rect 265070 167512 265126 167521
rect 265070 167447 265126 167456
rect 264980 167136 265032 167142
rect 264980 167078 265032 167084
rect 265084 167074 265112 167447
rect 265072 167068 265124 167074
rect 265072 167010 265124 167016
rect 264978 166696 265034 166705
rect 264978 166631 265034 166640
rect 264992 165646 265020 166631
rect 264980 165640 265032 165646
rect 264980 165582 265032 165588
rect 265070 165336 265126 165345
rect 265070 165271 265126 165280
rect 264978 164520 265034 164529
rect 264978 164455 265034 164464
rect 264992 164286 265020 164455
rect 265084 164354 265112 165271
rect 265072 164348 265124 164354
rect 265072 164290 265124 164296
rect 264980 164280 265032 164286
rect 264980 164222 265032 164228
rect 265070 164112 265126 164121
rect 265070 164047 265126 164056
rect 264978 163704 265034 163713
rect 264978 163639 265034 163648
rect 264518 163296 264574 163305
rect 264518 163231 264574 163240
rect 264334 156360 264390 156369
rect 264334 156295 264390 156304
rect 264244 131640 264296 131646
rect 264244 131582 264296 131588
rect 264242 128480 264298 128489
rect 264242 128415 264298 128424
rect 263140 123480 263192 123486
rect 263140 123422 263192 123428
rect 263140 118788 263192 118794
rect 263140 118730 263192 118736
rect 263152 102882 263180 118730
rect 263140 102876 263192 102882
rect 263140 102818 263192 102824
rect 263048 100700 263100 100706
rect 263048 100642 263100 100648
rect 263140 99476 263192 99482
rect 263140 99418 263192 99424
rect 263152 72457 263180 99418
rect 263138 72448 263194 72457
rect 263138 72383 263194 72392
rect 262954 61432 263010 61441
rect 262954 61367 263010 61376
rect 262864 46232 262916 46238
rect 262864 46174 262916 46180
rect 264256 42129 264284 128415
rect 264348 115938 264376 156295
rect 264426 146976 264482 146985
rect 264426 146911 264482 146920
rect 264336 115932 264388 115938
rect 264336 115874 264388 115880
rect 264334 110800 264390 110809
rect 264334 110735 264390 110744
rect 264348 51746 264376 110735
rect 264440 104825 264468 146911
rect 264532 122777 264560 163231
rect 264992 162994 265020 163639
rect 264980 162988 265032 162994
rect 264980 162930 265032 162936
rect 265084 162926 265112 164047
rect 265072 162920 265124 162926
rect 265072 162862 265124 162868
rect 264978 162344 265034 162353
rect 264978 162279 265034 162288
rect 264992 161498 265020 162279
rect 265176 162178 265204 168807
rect 265346 166288 265402 166297
rect 265346 166223 265402 166232
rect 265360 165714 265388 166223
rect 265714 165880 265770 165889
rect 265714 165815 265770 165824
rect 265348 165708 265400 165714
rect 265348 165650 265400 165656
rect 265622 164928 265678 164937
rect 265622 164863 265678 164872
rect 265164 162172 265216 162178
rect 265164 162114 265216 162120
rect 264980 161492 265032 161498
rect 264980 161434 265032 161440
rect 264978 161120 265034 161129
rect 264978 161055 265034 161064
rect 264992 160138 265020 161055
rect 264980 160132 265032 160138
rect 264980 160074 265032 160080
rect 265070 159760 265126 159769
rect 265070 159695 265126 159704
rect 264978 159352 265034 159361
rect 264978 159287 265034 159296
rect 264992 158778 265020 159287
rect 265084 158846 265112 159695
rect 265162 158944 265218 158953
rect 265162 158879 265218 158888
rect 265072 158840 265124 158846
rect 265072 158782 265124 158788
rect 264980 158772 265032 158778
rect 264980 158714 265032 158720
rect 265070 158128 265126 158137
rect 265070 158063 265126 158072
rect 264978 157720 265034 157729
rect 264978 157655 265034 157664
rect 264992 157418 265020 157655
rect 265084 157486 265112 158063
rect 265176 158001 265204 158879
rect 265254 158536 265310 158545
rect 265254 158471 265310 158480
rect 265162 157992 265218 158001
rect 265162 157927 265218 157936
rect 265072 157480 265124 157486
rect 265072 157422 265124 157428
rect 264980 157412 265032 157418
rect 264980 157354 265032 157360
rect 264978 157176 265034 157185
rect 264978 157111 265034 157120
rect 264992 155990 265020 157111
rect 265268 156670 265296 158471
rect 265256 156664 265308 156670
rect 265256 156606 265308 156612
rect 264980 155984 265032 155990
rect 264980 155926 265032 155932
rect 265070 155952 265126 155961
rect 265070 155887 265126 155896
rect 265084 154698 265112 155887
rect 265072 154692 265124 154698
rect 265072 154634 265124 154640
rect 264980 154624 265032 154630
rect 264978 154592 264980 154601
rect 265032 154592 265034 154601
rect 264978 154527 265034 154536
rect 265346 154184 265402 154193
rect 265346 154119 265402 154128
rect 265162 153776 265218 153785
rect 265162 153711 265218 153720
rect 265070 152960 265126 152969
rect 265070 152895 265126 152904
rect 264978 152008 265034 152017
rect 264978 151943 265034 151952
rect 264992 151910 265020 151943
rect 264980 151904 265032 151910
rect 264980 151846 265032 151852
rect 265084 151842 265112 152895
rect 265072 151836 265124 151842
rect 265072 151778 265124 151784
rect 264978 151192 265034 151201
rect 264978 151127 265034 151136
rect 264992 150482 265020 151127
rect 264980 150476 265032 150482
rect 264980 150418 265032 150424
rect 264978 149968 265034 149977
rect 264978 149903 265034 149912
rect 264992 149122 265020 149903
rect 265176 149734 265204 153711
rect 265360 153270 265388 154119
rect 265348 153264 265400 153270
rect 265348 153206 265400 153212
rect 265254 152552 265310 152561
rect 265254 152487 265310 152496
rect 265164 149728 265216 149734
rect 265164 149670 265216 149676
rect 264980 149116 265032 149122
rect 264980 149058 265032 149064
rect 264978 149016 265034 149025
rect 264978 148951 265034 148960
rect 264992 147694 265020 148951
rect 265070 148608 265126 148617
rect 265070 148543 265126 148552
rect 264980 147688 265032 147694
rect 264980 147630 265032 147636
rect 264978 147384 265034 147393
rect 264978 147319 265034 147328
rect 264992 146334 265020 147319
rect 265084 146946 265112 148543
rect 265268 148374 265296 152487
rect 265636 151094 265664 164863
rect 265728 153882 265756 165815
rect 279068 155938 279096 199446
rect 279148 188420 279200 188426
rect 279148 188362 279200 188368
rect 279160 161474 279188 188362
rect 280816 187678 280844 273974
rect 280908 244934 280936 306410
rect 282920 296812 282972 296818
rect 282920 296754 282972 296760
rect 281908 261520 281960 261526
rect 281908 261462 281960 261468
rect 280896 244928 280948 244934
rect 280896 244870 280948 244876
rect 281724 193860 281776 193866
rect 281724 193802 281776 193808
rect 280804 187672 280856 187678
rect 280804 187614 280856 187620
rect 280250 186960 280306 186969
rect 280250 186895 280306 186904
rect 279330 185736 279386 185745
rect 279330 185671 279386 185680
rect 279344 170649 279372 185671
rect 280160 185632 280212 185638
rect 280160 185574 280212 185580
rect 279424 175228 279476 175234
rect 279424 175170 279476 175176
rect 279436 174457 279464 175170
rect 279422 174448 279478 174457
rect 279422 174383 279478 174392
rect 279330 170640 279386 170649
rect 279330 170575 279386 170584
rect 280068 167068 280120 167074
rect 280068 167010 280120 167016
rect 280080 164937 280108 167010
rect 280066 164928 280122 164937
rect 280066 164863 280122 164872
rect 279160 161446 279372 161474
rect 279344 161401 279372 161446
rect 279330 161392 279386 161401
rect 279330 161327 279386 161336
rect 279330 155952 279386 155961
rect 279068 155910 279330 155938
rect 279330 155887 279386 155896
rect 267094 155544 267150 155553
rect 267094 155479 267150 155488
rect 265716 153876 265768 153882
rect 265716 153818 265768 153824
rect 265624 151088 265676 151094
rect 265624 151030 265676 151036
rect 265346 150784 265402 150793
rect 265346 150719 265402 150728
rect 265256 148368 265308 148374
rect 265256 148310 265308 148316
rect 265072 146940 265124 146946
rect 265072 146882 265124 146888
rect 264980 146328 265032 146334
rect 264980 146270 265032 146276
rect 265070 146024 265126 146033
rect 265070 145959 265126 145968
rect 264978 145208 265034 145217
rect 264978 145143 265034 145152
rect 264992 145042 265020 145143
rect 264980 145036 265032 145042
rect 264980 144978 265032 144984
rect 265084 144974 265112 145959
rect 265072 144968 265124 144974
rect 265072 144910 265124 144916
rect 265070 144800 265126 144809
rect 265070 144735 265126 144744
rect 264978 144392 265034 144401
rect 264978 144327 265034 144336
rect 264992 143614 265020 144327
rect 265084 143682 265112 144735
rect 265360 144129 265388 150719
rect 265898 149560 265954 149569
rect 265898 149495 265954 149504
rect 265346 144120 265402 144129
rect 265346 144055 265402 144064
rect 265162 143848 265218 143857
rect 265162 143783 265218 143792
rect 265072 143676 265124 143682
rect 265072 143618 265124 143624
rect 264980 143608 265032 143614
rect 264980 143550 265032 143556
rect 265070 143440 265126 143449
rect 265070 143375 265126 143384
rect 265084 142254 265112 143375
rect 265072 142248 265124 142254
rect 264978 142216 265034 142225
rect 265072 142190 265124 142196
rect 264978 142151 264980 142160
rect 265032 142151 265034 142160
rect 264980 142122 265032 142128
rect 264978 141808 265034 141817
rect 264978 141743 265034 141752
rect 264992 140826 265020 141743
rect 265176 141409 265204 143783
rect 265254 143032 265310 143041
rect 265254 142967 265310 142976
rect 265162 141400 265218 141409
rect 265162 141335 265218 141344
rect 265070 141264 265126 141273
rect 265070 141199 265126 141208
rect 264980 140820 265032 140826
rect 264980 140762 265032 140768
rect 264978 139632 265034 139641
rect 264978 139567 265034 139576
rect 264992 139466 265020 139567
rect 264980 139460 265032 139466
rect 264980 139402 265032 139408
rect 265084 138961 265112 141199
rect 265268 140894 265296 142967
rect 265256 140888 265308 140894
rect 265162 140856 265218 140865
rect 265256 140830 265308 140836
rect 265162 140791 265218 140800
rect 265176 139534 265204 140791
rect 265164 139528 265216 139534
rect 265164 139470 265216 139476
rect 265070 138952 265126 138961
rect 265070 138887 265126 138896
rect 264980 138712 265032 138718
rect 264980 138654 265032 138660
rect 265806 138680 265862 138689
rect 264992 138281 265020 138654
rect 265806 138615 265862 138624
rect 264978 138272 265034 138281
rect 264978 138207 265034 138216
rect 265070 137864 265126 137873
rect 265070 137799 265126 137808
rect 264978 137048 265034 137057
rect 264978 136983 265034 136992
rect 264992 136746 265020 136983
rect 264980 136740 265032 136746
rect 264980 136682 265032 136688
rect 265084 136678 265112 137799
rect 265072 136672 265124 136678
rect 265072 136614 265124 136620
rect 264978 136232 265034 136241
rect 264978 136167 265034 136176
rect 264992 135318 265020 136167
rect 264980 135312 265032 135318
rect 264980 135254 265032 135260
rect 265070 134872 265126 134881
rect 265070 134807 265126 134816
rect 264978 134056 265034 134065
rect 265084 134026 265112 134807
rect 265622 134192 265678 134201
rect 265622 134127 265678 134136
rect 264978 133991 265034 134000
rect 265072 134020 265124 134026
rect 264992 133958 265020 133991
rect 265072 133962 265124 133968
rect 264980 133952 265032 133958
rect 264980 133894 265032 133900
rect 265070 132288 265126 132297
rect 265070 132223 265126 132232
rect 264978 131880 265034 131889
rect 264978 131815 265034 131824
rect 264992 131170 265020 131815
rect 264980 131164 265032 131170
rect 264980 131106 265032 131112
rect 264978 130520 265034 130529
rect 264978 130455 265034 130464
rect 264992 129810 265020 130455
rect 264980 129804 265032 129810
rect 264980 129746 265032 129752
rect 264978 129296 265034 129305
rect 264978 129231 265034 129240
rect 264992 128382 265020 129231
rect 264980 128376 265032 128382
rect 264980 128318 265032 128324
rect 265084 127634 265112 132223
rect 265162 128888 265218 128897
rect 265162 128823 265218 128832
rect 265176 128450 265204 128823
rect 265164 128444 265216 128450
rect 265164 128386 265216 128392
rect 265072 127628 265124 127634
rect 265072 127570 265124 127576
rect 265070 126304 265126 126313
rect 265070 126239 265126 126248
rect 264978 125896 265034 125905
rect 264978 125831 265034 125840
rect 264992 125662 265020 125831
rect 265084 125730 265112 126239
rect 265072 125724 265124 125730
rect 265072 125666 265124 125672
rect 264980 125656 265032 125662
rect 264980 125598 265032 125604
rect 265070 125352 265126 125361
rect 265070 125287 265126 125296
rect 264978 124536 265034 124545
rect 264978 124471 265034 124480
rect 264992 124234 265020 124471
rect 265084 124302 265112 125287
rect 265072 124296 265124 124302
rect 265072 124238 265124 124244
rect 264980 124228 265032 124234
rect 264980 124170 265032 124176
rect 264978 124128 265034 124137
rect 264978 124063 265034 124072
rect 264992 122874 265020 124063
rect 264980 122868 265032 122874
rect 264980 122810 265032 122816
rect 264518 122768 264574 122777
rect 264518 122703 264574 122712
rect 264978 122360 265034 122369
rect 264978 122295 265034 122304
rect 264610 121544 264666 121553
rect 264992 121514 265020 122295
rect 264610 121479 264666 121488
rect 264980 121508 265032 121514
rect 264426 104816 264482 104825
rect 264426 104751 264482 104760
rect 264426 102640 264482 102649
rect 264426 102575 264482 102584
rect 264440 73817 264468 102575
rect 264624 84833 264652 121479
rect 264980 121450 265032 121456
rect 264978 120320 265034 120329
rect 264978 120255 265034 120264
rect 264992 120154 265020 120255
rect 264980 120148 265032 120154
rect 264980 120090 265032 120096
rect 264978 119776 265034 119785
rect 264978 119711 265034 119720
rect 264992 118726 265020 119711
rect 265438 118960 265494 118969
rect 265438 118895 265494 118904
rect 265452 118794 265480 118895
rect 265440 118788 265492 118794
rect 265440 118730 265492 118736
rect 264980 118720 265032 118726
rect 264980 118662 265032 118668
rect 265070 118144 265126 118153
rect 265070 118079 265126 118088
rect 264978 117736 265034 117745
rect 264978 117671 265034 117680
rect 264992 117434 265020 117671
rect 264980 117428 265032 117434
rect 264980 117370 265032 117376
rect 265084 117366 265112 118079
rect 265072 117360 265124 117366
rect 265072 117302 265124 117308
rect 265070 116784 265126 116793
rect 265070 116719 265126 116728
rect 265084 116074 265112 116719
rect 265072 116068 265124 116074
rect 265072 116010 265124 116016
rect 264980 116000 265032 116006
rect 264978 115968 264980 115977
rect 265032 115968 265034 115977
rect 264978 115903 265034 115912
rect 264978 115560 265034 115569
rect 264978 115495 265034 115504
rect 264992 114578 265020 115495
rect 264980 114572 265032 114578
rect 264980 114514 265032 114520
rect 264978 114200 265034 114209
rect 264978 114135 265034 114144
rect 264992 113626 265020 114135
rect 264980 113620 265032 113626
rect 264980 113562 265032 113568
rect 264978 112568 265034 112577
rect 264978 112503 265034 112512
rect 264992 111858 265020 112503
rect 264980 111852 265032 111858
rect 264980 111794 265032 111800
rect 264978 111616 265034 111625
rect 264978 111551 265034 111560
rect 264992 110498 265020 111551
rect 265070 111208 265126 111217
rect 265070 111143 265126 111152
rect 265084 110566 265112 111143
rect 265072 110560 265124 110566
rect 265072 110502 265124 110508
rect 264980 110492 265032 110498
rect 264980 110434 265032 110440
rect 265070 110392 265126 110401
rect 265070 110327 265126 110336
rect 264978 109576 265034 109585
rect 264978 109511 265034 109520
rect 264992 109070 265020 109511
rect 265084 109138 265112 110327
rect 265072 109132 265124 109138
rect 265072 109074 265124 109080
rect 264980 109064 265032 109070
rect 264980 109006 265032 109012
rect 265070 109032 265126 109041
rect 265070 108967 265126 108976
rect 264978 108624 265034 108633
rect 264978 108559 265034 108568
rect 264992 107710 265020 108559
rect 265084 107778 265112 108967
rect 265072 107772 265124 107778
rect 265072 107714 265124 107720
rect 264980 107704 265032 107710
rect 264980 107646 265032 107652
rect 264978 107400 265034 107409
rect 264978 107335 265034 107344
rect 264992 106350 265020 107335
rect 265070 106992 265126 107001
rect 265070 106927 265126 106936
rect 265084 106418 265112 106927
rect 265072 106412 265124 106418
rect 265072 106354 265124 106360
rect 264980 106344 265032 106350
rect 264980 106286 265032 106292
rect 264978 106040 265034 106049
rect 264978 105975 265034 105984
rect 264992 104922 265020 105975
rect 265070 105632 265126 105641
rect 265070 105567 265126 105576
rect 265084 104990 265112 105567
rect 265072 104984 265124 104990
rect 265072 104926 265124 104932
rect 264980 104916 265032 104922
rect 264980 104858 265032 104864
rect 264978 103864 265034 103873
rect 264978 103799 265034 103808
rect 264992 103562 265020 103799
rect 264980 103556 265032 103562
rect 264980 103498 265032 103504
rect 264978 103456 265034 103465
rect 264978 103391 265034 103400
rect 264992 102202 265020 103391
rect 265162 103048 265218 103057
rect 265162 102983 265218 102992
rect 265176 102270 265204 102983
rect 265164 102264 265216 102270
rect 265164 102206 265216 102212
rect 264980 102196 265032 102202
rect 264980 102138 265032 102144
rect 264978 101824 265034 101833
rect 264978 101759 265034 101768
rect 264992 100774 265020 101759
rect 264980 100768 265032 100774
rect 264980 100710 265032 100716
rect 264978 100464 265034 100473
rect 264978 100399 265034 100408
rect 264992 99414 265020 100399
rect 265070 100056 265126 100065
rect 265070 99991 265126 100000
rect 265084 99482 265112 99991
rect 265072 99476 265124 99482
rect 265072 99418 265124 99424
rect 264980 99408 265032 99414
rect 264980 99350 265032 99356
rect 265070 99240 265126 99249
rect 265070 99175 265126 99184
rect 264978 98696 265034 98705
rect 264978 98631 265034 98640
rect 264992 98054 265020 98631
rect 265084 98122 265112 99175
rect 265072 98116 265124 98122
rect 265072 98058 265124 98064
rect 264980 98048 265032 98054
rect 264980 97990 265032 97996
rect 264978 97880 265034 97889
rect 264978 97815 265034 97824
rect 264992 97306 265020 97815
rect 265070 97472 265126 97481
rect 265070 97407 265126 97416
rect 264980 97300 265032 97306
rect 264980 97242 265032 97248
rect 265084 96694 265112 97407
rect 265072 96688 265124 96694
rect 265072 96630 265124 96636
rect 264610 84824 264666 84833
rect 264610 84759 264666 84768
rect 264426 73808 264482 73817
rect 264426 73743 264482 73752
rect 265636 62937 265664 134127
rect 265714 132696 265770 132705
rect 265714 132631 265770 132640
rect 265728 65657 265756 132631
rect 265820 91866 265848 138615
rect 265912 134473 265940 149495
rect 265898 134464 265954 134473
rect 265898 134399 265954 134408
rect 267002 117192 267058 117201
rect 267002 117127 267058 117136
rect 265898 97064 265954 97073
rect 265898 96999 265954 97008
rect 265808 91860 265860 91866
rect 265808 91802 265860 91808
rect 265912 79393 265940 96999
rect 265898 79384 265954 79393
rect 265898 79319 265954 79328
rect 265714 65648 265770 65657
rect 265714 65583 265770 65592
rect 265622 62928 265678 62937
rect 265622 62863 265678 62872
rect 264336 51740 264388 51746
rect 264336 51682 264388 51688
rect 264242 42120 264298 42129
rect 264242 42055 264298 42064
rect 267016 36582 267044 117127
rect 267108 114510 267136 155479
rect 267188 131640 267240 131646
rect 267188 131582 267240 131588
rect 267096 114504 267148 114510
rect 267096 114446 267148 114452
rect 267094 104816 267150 104825
rect 267094 104751 267150 104760
rect 267004 36576 267056 36582
rect 267004 36518 267056 36524
rect 267108 33794 267136 104751
rect 267200 92478 267228 131582
rect 280172 129849 280200 185574
rect 280264 150385 280292 186895
rect 280342 180024 280398 180033
rect 280342 179959 280398 179968
rect 280356 174729 280384 179959
rect 281630 179480 281686 179489
rect 281630 179415 281686 179424
rect 280434 178936 280490 178945
rect 280434 178871 280490 178880
rect 280342 174720 280398 174729
rect 280342 174655 280398 174664
rect 280448 167074 280476 178871
rect 281540 169516 281592 169522
rect 281540 169458 281592 169464
rect 281552 169425 281580 169458
rect 281538 169416 281594 169425
rect 281538 169351 281594 169360
rect 280436 167068 280488 167074
rect 280436 167010 280488 167016
rect 281540 160268 281592 160274
rect 281540 160210 281592 160216
rect 281552 151881 281580 160210
rect 281538 151872 281594 151881
rect 281538 151807 281594 151816
rect 280250 150376 280306 150385
rect 280250 150311 280306 150320
rect 281644 142154 281672 179415
rect 281736 152697 281764 193802
rect 281816 182912 281868 182918
rect 281816 182854 281868 182860
rect 281828 160274 281856 182854
rect 281816 160268 281868 160274
rect 281816 160210 281868 160216
rect 281920 160154 281948 261462
rect 282184 201544 282236 201550
rect 282184 201486 282236 201492
rect 282196 180033 282224 201486
rect 282182 180024 282238 180033
rect 282182 179959 282238 179968
rect 282460 173868 282512 173874
rect 282460 173810 282512 173816
rect 282472 172553 282500 173810
rect 282458 172544 282514 172553
rect 282092 172508 282144 172514
rect 282458 172479 282514 172488
rect 282092 172450 282144 172456
rect 282104 171737 282132 172450
rect 282090 171728 282146 171737
rect 282090 171663 282146 171672
rect 282828 171080 282880 171086
rect 282828 171022 282880 171028
rect 282840 170921 282868 171022
rect 282826 170912 282882 170921
rect 282826 170847 282882 170856
rect 282828 169448 282880 169454
rect 282828 169390 282880 169396
rect 282840 168745 282868 169390
rect 282826 168736 282882 168745
rect 282826 168671 282882 168680
rect 282828 167748 282880 167754
rect 282828 167690 282880 167696
rect 282840 167113 282868 167690
rect 282826 167104 282882 167113
rect 282826 167039 282882 167048
rect 282828 167000 282880 167006
rect 282828 166942 282880 166948
rect 282840 166433 282868 166942
rect 282826 166424 282882 166433
rect 282826 166359 282882 166368
rect 281998 165608 282054 165617
rect 281998 165543 282000 165552
rect 282052 165543 282054 165552
rect 282000 165514 282052 165520
rect 282828 164212 282880 164218
rect 282828 164154 282880 164160
rect 282460 164144 282512 164150
rect 282840 164121 282868 164154
rect 282460 164086 282512 164092
rect 282826 164112 282882 164121
rect 282472 163305 282500 164086
rect 282826 164047 282882 164056
rect 282458 163296 282514 163305
rect 282458 163231 282514 163240
rect 282828 162852 282880 162858
rect 282828 162794 282880 162800
rect 282840 162625 282868 162794
rect 282826 162616 282882 162625
rect 282826 162551 282882 162560
rect 282826 161800 282882 161809
rect 282932 161786 282960 296754
rect 284298 287192 284354 287201
rect 284298 287127 284354 287136
rect 283102 215928 283158 215937
rect 283102 215863 283158 215872
rect 283012 204944 283064 204950
rect 283012 204886 283064 204892
rect 282882 161758 282960 161786
rect 282826 161735 282882 161744
rect 282826 160304 282882 160313
rect 282826 160239 282882 160248
rect 282840 160206 282868 160239
rect 281828 160126 281948 160154
rect 282828 160200 282880 160206
rect 282828 160142 282880 160148
rect 281828 156505 281856 160126
rect 281908 160064 281960 160070
rect 281908 160006 281960 160012
rect 281920 159497 281948 160006
rect 282368 159996 282420 160002
rect 282368 159938 282420 159944
rect 281906 159488 281962 159497
rect 281906 159423 281962 159432
rect 282380 158817 282408 159938
rect 282366 158808 282422 158817
rect 282366 158743 282422 158752
rect 282092 158704 282144 158710
rect 282092 158646 282144 158652
rect 282104 158001 282132 158646
rect 282090 157992 282146 158001
rect 282090 157927 282146 157936
rect 281814 156496 281870 156505
rect 281814 156431 281870 156440
rect 282276 155916 282328 155922
rect 282276 155858 282328 155864
rect 282288 155009 282316 155858
rect 282274 155000 282330 155009
rect 282274 154935 282330 154944
rect 282276 154556 282328 154562
rect 282276 154498 282328 154504
rect 282288 153513 282316 154498
rect 282828 154488 282880 154494
rect 282828 154430 282880 154436
rect 282840 154193 282868 154430
rect 282826 154184 282882 154193
rect 282826 154119 282882 154128
rect 282274 153504 282330 153513
rect 282274 153439 282330 153448
rect 281722 152688 281778 152697
rect 281722 152623 281778 152632
rect 281908 151768 281960 151774
rect 281908 151710 281960 151716
rect 281920 151201 281948 151710
rect 281906 151192 281962 151201
rect 281906 151127 281962 151136
rect 282828 149048 282880 149054
rect 282828 148990 282880 148996
rect 282642 148880 282698 148889
rect 282642 148815 282698 148824
rect 282656 147898 282684 148815
rect 282840 148073 282868 148990
rect 282826 148064 282882 148073
rect 282826 147999 282882 148008
rect 282644 147892 282696 147898
rect 282644 147834 282696 147840
rect 282828 147620 282880 147626
rect 282828 147562 282880 147568
rect 282276 147552 282328 147558
rect 282276 147494 282328 147500
rect 282288 146577 282316 147494
rect 282840 147393 282868 147562
rect 282826 147384 282882 147393
rect 282826 147319 282882 147328
rect 282274 146568 282330 146577
rect 282274 146503 282330 146512
rect 282828 146260 282880 146266
rect 282828 146202 282880 146208
rect 282736 146192 282788 146198
rect 282736 146134 282788 146140
rect 282748 145081 282776 146134
rect 282840 145897 282868 146202
rect 282826 145888 282882 145897
rect 282826 145823 282882 145832
rect 282734 145072 282790 145081
rect 282734 145007 282790 145016
rect 282828 144900 282880 144906
rect 282828 144842 282880 144848
rect 282840 144265 282868 144842
rect 282826 144256 282882 144265
rect 282826 144191 282882 144200
rect 282828 143540 282880 143546
rect 282828 143482 282880 143488
rect 282840 142769 282868 143482
rect 282826 142760 282882 142769
rect 282826 142695 282882 142704
rect 281552 142126 281672 142154
rect 281552 138961 281580 142126
rect 282552 142112 282604 142118
rect 282550 142080 282552 142089
rect 282604 142080 282606 142089
rect 282550 142015 282606 142024
rect 282828 141364 282880 141370
rect 282828 141306 282880 141312
rect 282840 141273 282868 141306
rect 282826 141264 282882 141273
rect 282826 141199 282882 141208
rect 282828 140752 282880 140758
rect 282828 140694 282880 140700
rect 282840 139777 282868 140694
rect 282826 139768 282882 139777
rect 282826 139703 282882 139712
rect 281538 138952 281594 138961
rect 281538 138887 281594 138896
rect 281540 138372 281592 138378
rect 281540 138314 281592 138320
rect 281552 138281 281580 138314
rect 281538 138272 281594 138281
rect 281538 138207 281594 138216
rect 282828 137488 282880 137494
rect 282826 137456 282828 137465
rect 282880 137456 282882 137465
rect 282826 137391 282882 137400
rect 282826 136640 282882 136649
rect 282826 136575 282828 136584
rect 282880 136575 282882 136584
rect 282828 136546 282880 136552
rect 282828 133884 282880 133890
rect 282828 133826 282880 133832
rect 282840 132841 282868 133826
rect 282826 132832 282882 132841
rect 282826 132767 282882 132776
rect 282828 132456 282880 132462
rect 282828 132398 282880 132404
rect 282840 132161 282868 132398
rect 282826 132152 282882 132161
rect 282826 132087 282882 132096
rect 282276 131028 282328 131034
rect 282276 130970 282328 130976
rect 282288 130665 282316 130970
rect 282274 130656 282330 130665
rect 282274 130591 282330 130600
rect 280158 129840 280214 129849
rect 280158 129775 280214 129784
rect 282092 129736 282144 129742
rect 282092 129678 282144 129684
rect 282104 129033 282132 129678
rect 282090 129024 282146 129033
rect 282090 128959 282146 128968
rect 282826 128344 282882 128353
rect 282000 128308 282052 128314
rect 282826 128279 282882 128288
rect 282000 128250 282052 128256
rect 282012 127537 282040 128250
rect 282840 128246 282868 128279
rect 282828 128240 282880 128246
rect 282828 128182 282880 128188
rect 281998 127528 282054 127537
rect 281998 127463 282054 127472
rect 282276 126948 282328 126954
rect 282276 126890 282328 126896
rect 279330 126304 279386 126313
rect 279330 126239 279386 126248
rect 267646 123720 267702 123729
rect 267646 123655 267702 123664
rect 267660 94518 267688 123655
rect 279344 122834 279372 126239
rect 282288 126041 282316 126890
rect 282274 126032 282330 126041
rect 282274 125967 282330 125976
rect 282828 125588 282880 125594
rect 282828 125530 282880 125536
rect 282736 125520 282788 125526
rect 282736 125462 282788 125468
rect 282748 124545 282776 125462
rect 282840 125225 282868 125530
rect 282826 125216 282882 125225
rect 282826 125151 282882 125160
rect 282734 124536 282790 124545
rect 282734 124471 282790 124480
rect 282276 124160 282328 124166
rect 282276 124102 282328 124108
rect 282288 123049 282316 124102
rect 282828 124092 282880 124098
rect 282828 124034 282880 124040
rect 282840 123729 282868 124034
rect 282826 123720 282882 123729
rect 282826 123655 282882 123664
rect 282274 123040 282330 123049
rect 282274 122975 282330 122984
rect 283024 122834 283052 204886
rect 283116 135153 283144 215863
rect 283196 188352 283248 188358
rect 283196 188294 283248 188300
rect 283208 169522 283236 188294
rect 283196 169516 283248 169522
rect 283196 169458 283248 169464
rect 283102 135144 283158 135153
rect 283102 135079 283158 135088
rect 279068 122806 279372 122834
rect 282932 122806 283052 122834
rect 267738 109984 267794 109993
rect 267738 109919 267794 109928
rect 267648 94512 267700 94518
rect 267648 94454 267700 94460
rect 267188 92472 267240 92478
rect 267188 92414 267240 92420
rect 267752 53106 267780 109919
rect 269120 94512 269172 94518
rect 269120 94454 269172 94460
rect 267740 53100 267792 53106
rect 267740 53042 267792 53048
rect 267740 47592 267792 47598
rect 267740 47534 267792 47540
rect 267096 33788 267148 33794
rect 267096 33730 267148 33736
rect 267004 31136 267056 31142
rect 267004 31078 267056 31084
rect 263600 24200 263652 24206
rect 263600 24142 263652 24148
rect 263612 16574 263640 24142
rect 262232 16546 262536 16574
rect 263612 16546 264192 16574
rect 261758 13016 261814 13025
rect 261758 12951 261814 12960
rect 260654 4040 260710 4049
rect 260654 3975 260710 3984
rect 260668 480 260696 3975
rect 261772 480 261800 12951
rect 262508 490 262536 16546
rect 262784 598 262996 626
rect 262784 490 262812 598
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 462 262812 490
rect 262968 480 262996 598
rect 264164 480 264192 16546
rect 265346 4856 265402 4865
rect 265346 4791 265402 4800
rect 265360 480 265388 4791
rect 267016 3466 267044 31078
rect 266544 3460 266596 3466
rect 266544 3402 266596 3408
rect 267004 3460 267056 3466
rect 267004 3402 267056 3408
rect 266556 480 266584 3402
rect 267752 480 267780 47534
rect 269132 43450 269160 94454
rect 274008 93770 274036 96084
rect 278778 95840 278834 95849
rect 278778 95775 278834 95784
rect 278792 95198 278820 95775
rect 278780 95192 278832 95198
rect 278780 95134 278832 95140
rect 273996 93764 274048 93770
rect 273996 93706 274048 93712
rect 270498 93120 270554 93129
rect 270498 93055 270554 93064
rect 269120 43444 269172 43450
rect 269120 43386 269172 43392
rect 270512 16574 270540 93055
rect 279068 86873 279096 122806
rect 282828 122800 282880 122806
rect 282828 122742 282880 122748
rect 282840 122233 282868 122742
rect 282826 122224 282882 122233
rect 282826 122159 282882 122168
rect 282828 121440 282880 121446
rect 282826 121408 282828 121417
rect 282880 121408 282882 121417
rect 282826 121343 282882 121352
rect 282826 120728 282882 120737
rect 282932 120714 282960 122806
rect 282882 120686 282960 120714
rect 282826 120663 282882 120672
rect 282828 120080 282880 120086
rect 282828 120022 282880 120028
rect 282736 120012 282788 120018
rect 282736 119954 282788 119960
rect 282748 119241 282776 119954
rect 282840 119921 282868 120022
rect 282826 119912 282882 119921
rect 282826 119847 282882 119856
rect 282734 119232 282790 119241
rect 282734 119167 282790 119176
rect 282828 118652 282880 118658
rect 282828 118594 282880 118600
rect 282276 118584 282328 118590
rect 282276 118526 282328 118532
rect 282288 117609 282316 118526
rect 282840 118425 282868 118594
rect 282826 118416 282882 118425
rect 282826 118351 282882 118360
rect 282274 117600 282330 117609
rect 282274 117535 282330 117544
rect 282828 117292 282880 117298
rect 282828 117234 282880 117240
rect 282840 116113 282868 117234
rect 282826 116104 282882 116113
rect 282826 116039 282882 116048
rect 282368 115932 282420 115938
rect 282368 115874 282420 115880
rect 282380 114617 282408 115874
rect 282828 115864 282880 115870
rect 282828 115806 282880 115812
rect 282840 115433 282868 115806
rect 282826 115424 282882 115433
rect 282826 115359 282882 115368
rect 282366 114608 282422 114617
rect 282366 114543 282422 114552
rect 282092 114504 282144 114510
rect 282092 114446 282144 114452
rect 282104 113801 282132 114446
rect 282090 113792 282146 113801
rect 282090 113727 282146 113736
rect 282828 113144 282880 113150
rect 282458 113112 282514 113121
rect 282828 113086 282880 113092
rect 282458 113047 282460 113056
rect 282512 113047 282514 113056
rect 282460 113018 282512 113024
rect 282840 112305 282868 113086
rect 282826 112296 282882 112305
rect 282826 112231 282882 112240
rect 282828 111784 282880 111790
rect 282828 111726 282880 111732
rect 281724 111648 281776 111654
rect 281722 111616 281724 111625
rect 281776 111616 281778 111625
rect 281722 111551 281778 111560
rect 282840 110809 282868 111726
rect 284312 111654 284340 287127
rect 285680 249076 285732 249082
rect 285680 249018 285732 249024
rect 284390 196752 284446 196761
rect 284390 196687 284446 196696
rect 284300 111648 284352 111654
rect 284300 111590 284352 111596
rect 282826 110800 282882 110809
rect 282826 110735 282882 110744
rect 282276 110424 282328 110430
rect 282276 110366 282328 110372
rect 282288 109313 282316 110366
rect 282828 110356 282880 110362
rect 282828 110298 282880 110304
rect 282840 109993 282868 110298
rect 282826 109984 282882 109993
rect 282826 109919 282882 109928
rect 282274 109304 282330 109313
rect 282274 109239 282330 109248
rect 282368 108996 282420 109002
rect 282368 108938 282420 108944
rect 282380 107817 282408 108938
rect 282826 108488 282882 108497
rect 282826 108423 282882 108432
rect 282840 107982 282868 108423
rect 282828 107976 282880 107982
rect 282828 107918 282880 107924
rect 282366 107808 282422 107817
rect 282366 107743 282422 107752
rect 282828 106276 282880 106282
rect 282828 106218 282880 106224
rect 282840 105505 282868 106218
rect 282826 105496 282882 105505
rect 282826 105431 282882 105440
rect 282828 104848 282880 104854
rect 282828 104790 282880 104796
rect 281538 104680 281594 104689
rect 281538 104615 281594 104624
rect 279330 98152 279386 98161
rect 279330 98087 279386 98096
rect 279344 95169 279372 98087
rect 279330 95160 279386 95169
rect 279330 95095 279386 95104
rect 281552 92478 281580 104615
rect 282840 104009 282868 104790
rect 282826 104000 282882 104009
rect 282826 103935 282882 103944
rect 282828 103488 282880 103494
rect 282828 103430 282880 103436
rect 282840 103193 282868 103430
rect 282826 103184 282882 103193
rect 282826 103119 282882 103128
rect 284404 102066 284432 196687
rect 284484 182844 284536 182850
rect 284484 182786 284536 182792
rect 284496 138378 284524 182786
rect 284576 176044 284628 176050
rect 284576 175986 284628 175992
rect 284588 165578 284616 175986
rect 284576 165572 284628 165578
rect 284576 165514 284628 165520
rect 284484 138372 284536 138378
rect 284484 138314 284536 138320
rect 285692 131034 285720 249018
rect 285772 200796 285824 200802
rect 285772 200738 285824 200744
rect 285680 131028 285732 131034
rect 285680 130970 285732 130976
rect 285784 113082 285812 200738
rect 286336 186969 286364 307838
rect 295340 305040 295392 305046
rect 295340 304982 295392 304988
rect 298098 305008 298154 305017
rect 289912 291304 289964 291310
rect 289912 291246 289964 291252
rect 288440 256012 288492 256018
rect 288440 255954 288492 255960
rect 287060 250504 287112 250510
rect 287060 250446 287112 250452
rect 286322 186960 286378 186969
rect 286322 186895 286378 186904
rect 285954 184376 286010 184385
rect 285954 184311 286010 184320
rect 285864 177404 285916 177410
rect 285864 177346 285916 177352
rect 285876 142118 285904 177346
rect 285968 164150 285996 184311
rect 285956 164144 286008 164150
rect 285956 164086 286008 164092
rect 285864 142112 285916 142118
rect 285864 142054 285916 142060
rect 287072 137494 287100 250446
rect 287336 192500 287388 192506
rect 287336 192442 287388 192448
rect 287152 178696 287204 178702
rect 287152 178638 287204 178644
rect 287060 137488 287112 137494
rect 287060 137430 287112 137436
rect 285772 113076 285824 113082
rect 285772 113018 285824 113024
rect 287164 107982 287192 178638
rect 287244 177336 287296 177342
rect 287244 177278 287296 177284
rect 287256 147898 287284 177278
rect 287348 169454 287376 192442
rect 287336 169448 287388 169454
rect 287336 169390 287388 169396
rect 287244 147892 287296 147898
rect 287244 147834 287296 147840
rect 288452 141370 288480 255954
rect 289818 229120 289874 229129
rect 289818 229055 289874 229064
rect 288624 187672 288676 187678
rect 288624 187614 288676 187620
rect 288532 180124 288584 180130
rect 288532 180066 288584 180072
rect 288440 141364 288492 141370
rect 288440 141306 288492 141312
rect 288544 120018 288572 180066
rect 288636 160206 288664 187614
rect 288714 177304 288770 177313
rect 288714 177239 288770 177248
rect 288728 167754 288756 177239
rect 288716 167748 288768 167754
rect 288716 167690 288768 167696
rect 288624 160200 288676 160206
rect 288624 160142 288676 160148
rect 288532 120012 288584 120018
rect 288532 119954 288584 119960
rect 289832 111790 289860 229055
rect 289924 173874 289952 291246
rect 294052 267028 294104 267034
rect 294052 266970 294104 266976
rect 291200 259480 291252 259486
rect 291200 259422 291252 259428
rect 290002 213208 290058 213217
rect 290002 213143 290058 213152
rect 289912 173868 289964 173874
rect 289912 173810 289964 173816
rect 289820 111784 289872 111790
rect 289820 111726 289872 111732
rect 287152 107976 287204 107982
rect 287152 107918 287204 107924
rect 290016 103494 290044 213143
rect 290094 180024 290150 180033
rect 290094 179959 290150 179968
rect 290108 160002 290136 179959
rect 290096 159996 290148 160002
rect 290096 159938 290148 159944
rect 291212 113150 291240 259422
rect 292580 234660 292632 234666
rect 292580 234602 292632 234608
rect 291382 214568 291438 214577
rect 291382 214503 291438 214512
rect 291292 200864 291344 200870
rect 291292 200806 291344 200812
rect 291200 113144 291252 113150
rect 291200 113086 291252 113092
rect 291304 106282 291332 200806
rect 291396 167006 291424 214503
rect 291474 178800 291530 178809
rect 291474 178735 291530 178744
rect 291384 167000 291436 167006
rect 291384 166942 291436 166948
rect 291488 140758 291516 178735
rect 291476 140752 291528 140758
rect 291476 140694 291528 140700
rect 291292 106276 291344 106282
rect 291292 106218 291344 106224
rect 292592 104854 292620 234602
rect 292672 231872 292724 231878
rect 292672 231814 292724 231820
rect 292684 118590 292712 231814
rect 292764 191140 292816 191146
rect 292764 191082 292816 191088
rect 292776 162858 292804 191082
rect 293960 186380 294012 186386
rect 293960 186322 294012 186328
rect 292856 180192 292908 180198
rect 292856 180134 292908 180140
rect 292764 162852 292816 162858
rect 292764 162794 292816 162800
rect 292868 154494 292896 180134
rect 292856 154488 292908 154494
rect 292856 154430 292908 154436
rect 292672 118584 292724 118590
rect 292672 118526 292724 118532
rect 292580 104848 292632 104854
rect 292580 104790 292632 104796
rect 290004 103488 290056 103494
rect 290004 103430 290056 103436
rect 281724 102060 281776 102066
rect 281724 102002 281776 102008
rect 284392 102060 284444 102066
rect 284392 102002 284444 102008
rect 281736 101697 281764 102002
rect 281722 101688 281778 101697
rect 281722 101623 281778 101632
rect 281630 100872 281686 100881
rect 281630 100807 281686 100816
rect 281644 93838 281672 100807
rect 281724 100700 281776 100706
rect 281724 100642 281776 100648
rect 281736 100201 281764 100642
rect 281722 100192 281778 100201
rect 281722 100127 281778 100136
rect 282826 99376 282882 99385
rect 282826 99311 282828 99320
rect 282880 99311 282882 99320
rect 282828 99282 282880 99288
rect 282184 97980 282236 97986
rect 282184 97922 282236 97928
rect 282196 97073 282224 97922
rect 282828 97912 282880 97918
rect 282826 97880 282828 97889
rect 282880 97880 282882 97889
rect 282826 97815 282882 97824
rect 282182 97064 282238 97073
rect 282182 96999 282238 97008
rect 281632 93832 281684 93838
rect 281632 93774 281684 93780
rect 281540 92472 281592 92478
rect 281540 92414 281592 92420
rect 280158 89040 280214 89049
rect 280158 88975 280214 88984
rect 279054 86864 279110 86873
rect 279054 86799 279110 86808
rect 273260 77988 273312 77994
rect 273260 77930 273312 77936
rect 270512 16546 270816 16574
rect 269762 15872 269818 15881
rect 269762 15807 269818 15816
rect 269670 14512 269726 14521
rect 269670 14447 269726 14456
rect 268382 11656 268438 11665
rect 268382 11591 268438 11600
rect 268396 490 268424 11591
rect 269684 2938 269712 14447
rect 269776 3126 269804 15807
rect 269764 3120 269816 3126
rect 269764 3062 269816 3068
rect 269684 2910 270080 2938
rect 268672 598 268884 626
rect 268672 490 268700 598
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 462 268700 490
rect 268856 480 268884 598
rect 270052 480 270080 2910
rect 270788 490 270816 16546
rect 272432 3120 272484 3126
rect 272432 3062 272484 3068
rect 271064 598 271276 626
rect 271064 490 271092 598
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270788 462 271092 490
rect 271248 480 271276 598
rect 272444 480 272472 3062
rect 273272 490 273300 77930
rect 278778 72584 278834 72593
rect 278778 72519 278834 72528
rect 276018 67008 276074 67017
rect 276018 66943 276074 66952
rect 276032 3602 276060 66943
rect 276110 39264 276166 39273
rect 276110 39199 276166 39208
rect 276020 3596 276072 3602
rect 276020 3538 276072 3544
rect 276124 3482 276152 39199
rect 278792 16574 278820 72519
rect 280172 16574 280200 88975
rect 281540 84856 281592 84862
rect 281540 84798 281592 84804
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 278318 6216 278374 6225
rect 278318 6151 278374 6160
rect 277124 3596 277176 3602
rect 277124 3538 277176 3544
rect 274824 3460 274876 3466
rect 274824 3402 274876 3408
rect 276032 3454 276152 3482
rect 273456 598 273668 626
rect 273456 490 273484 598
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 462 273484 490
rect 273640 480 273668 598
rect 274836 480 274864 3402
rect 276032 480 276060 3454
rect 277136 480 277164 3538
rect 278332 480 278360 6151
rect 279068 490 279096 16546
rect 279344 598 279556 626
rect 279344 490 279372 598
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 462 279372 490
rect 279528 480 279556 598
rect 280724 480 280752 16546
rect 281446 8936 281502 8945
rect 281446 8871 281502 8880
rect 281460 3534 281488 8871
rect 281448 3528 281500 3534
rect 281448 3470 281500 3476
rect 281552 490 281580 84798
rect 284298 75168 284354 75177
rect 284298 75103 284354 75112
rect 283104 3528 283156 3534
rect 283104 3470 283156 3476
rect 281736 598 281948 626
rect 281736 490 281764 598
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281552 462 281764 490
rect 281920 480 281948 598
rect 283116 480 283144 3470
rect 284312 480 284340 75103
rect 289820 18624 289872 18630
rect 289820 18566 289872 18572
rect 286598 3496 286654 3505
rect 285404 3460 285456 3466
rect 286598 3431 286654 3440
rect 287794 3496 287850 3505
rect 287794 3431 287850 3440
rect 288990 3496 289046 3505
rect 288990 3431 289046 3440
rect 285404 3402 285456 3408
rect 285416 480 285444 3402
rect 286612 480 286640 3431
rect 287808 480 287836 3431
rect 289004 480 289032 3431
rect 289832 490 289860 18566
rect 293972 6914 294000 186322
rect 294064 124098 294092 266970
rect 294144 221468 294196 221474
rect 294144 221410 294196 221416
rect 294156 146198 294184 221410
rect 294236 178764 294288 178770
rect 294236 178706 294288 178712
rect 294248 160070 294276 178706
rect 294236 160064 294288 160070
rect 294236 160006 294288 160012
rect 294144 146192 294196 146198
rect 294144 146134 294196 146140
rect 295352 143546 295380 304982
rect 298098 304943 298154 304952
rect 296720 264240 296772 264246
rect 296720 264182 296772 264188
rect 295432 254584 295484 254590
rect 295432 254526 295484 254532
rect 295340 143540 295392 143546
rect 295340 143482 295392 143488
rect 294052 124092 294104 124098
rect 294052 124034 294104 124040
rect 295444 97918 295472 254526
rect 295524 233300 295576 233306
rect 295524 233242 295576 233248
rect 295536 109002 295564 233242
rect 295616 206304 295668 206310
rect 295616 206246 295668 206252
rect 295628 172514 295656 206246
rect 295616 172508 295668 172514
rect 295616 172450 295668 172456
rect 296732 126954 296760 264182
rect 296812 253224 296864 253230
rect 296812 253166 296864 253172
rect 296720 126948 296772 126954
rect 296720 126890 296772 126896
rect 296824 124166 296852 253166
rect 296902 194032 296958 194041
rect 296902 193967 296958 193976
rect 296916 136610 296944 193967
rect 296904 136604 296956 136610
rect 296904 136546 296956 136552
rect 296812 124160 296864 124166
rect 296812 124102 296864 124108
rect 298112 110362 298140 304943
rect 299570 302424 299626 302433
rect 299570 302359 299626 302368
rect 298192 302320 298244 302326
rect 298192 302262 298244 302268
rect 298204 171086 298232 302262
rect 298284 242208 298336 242214
rect 298284 242150 298336 242156
rect 298192 171080 298244 171086
rect 298192 171022 298244 171028
rect 298296 147558 298324 242150
rect 299478 220144 299534 220153
rect 299478 220079 299534 220088
rect 298376 181484 298428 181490
rect 298376 181426 298428 181432
rect 298284 147552 298336 147558
rect 298284 147494 298336 147500
rect 298100 110356 298152 110362
rect 298100 110298 298152 110304
rect 295524 108996 295576 109002
rect 295524 108938 295576 108944
rect 298388 97986 298416 181426
rect 298376 97980 298428 97986
rect 298376 97922 298428 97928
rect 295432 97912 295484 97918
rect 295432 97854 295484 97860
rect 296720 17264 296772 17270
rect 296720 17206 296772 17212
rect 296732 16574 296760 17206
rect 296732 16546 297312 16574
rect 293696 6886 294000 6914
rect 291382 3496 291438 3505
rect 291382 3431 291438 3440
rect 290016 598 290228 626
rect 290016 490 290044 598
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289832 462 290044 490
rect 290200 480 290228 598
rect 291396 480 291424 3431
rect 292580 2848 292632 2854
rect 292580 2790 292632 2796
rect 292592 480 292620 2790
rect 293696 480 293724 6886
rect 296076 3528 296128 3534
rect 296076 3470 296128 3476
rect 294878 3360 294934 3369
rect 294878 3295 294934 3304
rect 294892 480 294920 3295
rect 296088 480 296116 3470
rect 297284 480 297312 16546
rect 298466 7576 298522 7585
rect 298466 7511 298522 7520
rect 298480 480 298508 7511
rect 299492 3534 299520 220079
rect 299584 110430 299612 302359
rect 300952 258732 301004 258738
rect 300952 258674 301004 258680
rect 299756 228404 299808 228410
rect 299756 228346 299808 228352
rect 299662 192536 299718 192545
rect 299662 192471 299718 192480
rect 299572 110424 299624 110430
rect 299572 110366 299624 110372
rect 299676 16574 299704 192471
rect 299768 144906 299796 228346
rect 300858 207632 300914 207641
rect 300858 207567 300914 207576
rect 299756 144900 299808 144906
rect 299756 144842 299808 144848
rect 300872 16574 300900 207567
rect 300964 158710 300992 258674
rect 301044 191208 301096 191214
rect 301044 191150 301096 191156
rect 300952 158704 301004 158710
rect 300952 158646 301004 158652
rect 301056 129742 301084 191150
rect 301044 129736 301096 129742
rect 301044 129678 301096 129684
rect 302252 120086 302280 314638
rect 304262 300928 304318 300937
rect 304262 300863 304318 300872
rect 302332 240168 302384 240174
rect 302332 240110 302384 240116
rect 302240 120080 302292 120086
rect 302240 120022 302292 120028
rect 302344 100706 302372 240110
rect 303804 236700 303856 236706
rect 303804 236642 303856 236648
rect 302516 213240 302568 213246
rect 302516 213182 302568 213188
rect 302424 210452 302476 210458
rect 302424 210394 302476 210400
rect 302436 121446 302464 210394
rect 302528 154562 302556 213182
rect 303712 203584 303764 203590
rect 303712 203526 303764 203532
rect 303618 188320 303674 188329
rect 303618 188255 303674 188264
rect 302516 154556 302568 154562
rect 302516 154498 302568 154504
rect 302424 121440 302476 121446
rect 302424 121382 302476 121388
rect 302332 100700 302384 100706
rect 302332 100642 302384 100648
rect 303632 16574 303660 188255
rect 303724 117298 303752 203526
rect 303816 164218 303844 236642
rect 304276 188358 304304 300863
rect 304264 188352 304316 188358
rect 304264 188294 304316 188300
rect 303896 184204 303948 184210
rect 303896 184146 303948 184152
rect 303804 164212 303856 164218
rect 303804 164154 303856 164160
rect 303712 117292 303764 117298
rect 303712 117234 303764 117240
rect 303908 115870 303936 184146
rect 303896 115864 303948 115870
rect 303896 115806 303948 115812
rect 299676 16546 299796 16574
rect 300872 16546 301544 16574
rect 303632 16546 303936 16574
rect 299664 14544 299716 14550
rect 299664 14486 299716 14492
rect 299480 3528 299532 3534
rect 299480 3470 299532 3476
rect 299676 480 299704 14486
rect 299768 3369 299796 16546
rect 300766 3496 300822 3505
rect 300766 3431 300822 3440
rect 299754 3360 299810 3369
rect 299754 3295 299810 3304
rect 300780 480 300808 3431
rect 301516 490 301544 16546
rect 303160 6180 303212 6186
rect 303160 6122 303212 6128
rect 301792 598 302004 626
rect 301792 490 301820 598
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 462 301820 490
rect 301976 480 302004 598
rect 303172 480 303200 6122
rect 303908 490 303936 16546
rect 305012 6225 305040 365706
rect 305644 316736 305696 316742
rect 305644 316678 305696 316684
rect 305092 227044 305144 227050
rect 305092 226986 305144 226992
rect 305104 115938 305132 226986
rect 305184 199436 305236 199442
rect 305184 199378 305236 199384
rect 305196 147626 305224 199378
rect 305184 147620 305236 147626
rect 305184 147562 305236 147568
rect 305092 115932 305144 115938
rect 305092 115874 305144 115880
rect 305656 6914 305684 316678
rect 306564 246356 306616 246362
rect 306564 246298 306616 246304
rect 306470 203552 306526 203561
rect 306470 203487 306526 203496
rect 305564 6886 305684 6914
rect 304998 6216 305054 6225
rect 304998 6151 305054 6160
rect 304184 598 304396 626
rect 304184 490 304212 598
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 303908 462 304212 490
rect 304368 480 304396 598
rect 305564 480 305592 6886
rect 306484 3466 306512 203487
rect 306576 149054 306604 246298
rect 306656 220108 306708 220114
rect 306656 220050 306708 220056
rect 306564 149048 306616 149054
rect 306564 148990 306616 148996
rect 306668 128246 306696 220050
rect 306656 128240 306708 128246
rect 306656 128182 306708 128188
rect 306472 3460 306524 3466
rect 306472 3402 306524 3408
rect 306760 480 306788 368494
rect 321558 367160 321614 367169
rect 321558 367095 321614 367104
rect 313922 336832 313978 336841
rect 313922 336767 313978 336776
rect 309138 319424 309194 319433
rect 309138 319359 309194 319368
rect 307758 231160 307814 231169
rect 307758 231095 307814 231104
rect 307772 114510 307800 231095
rect 307852 224256 307904 224262
rect 307852 224198 307904 224204
rect 307864 151774 307892 224198
rect 307944 189780 307996 189786
rect 307944 189722 307996 189728
rect 307852 151768 307904 151774
rect 307852 151710 307904 151716
rect 307956 122806 307984 189722
rect 307944 122800 307996 122806
rect 307944 122742 307996 122748
rect 307760 114504 307812 114510
rect 307760 114446 307812 114452
rect 307758 65512 307814 65521
rect 307758 65447 307814 65456
rect 307772 3534 307800 65447
rect 309152 16574 309180 319359
rect 313280 283892 313332 283898
rect 313280 283834 313332 283840
rect 311900 273964 311952 273970
rect 311900 273906 311952 273912
rect 310612 262880 310664 262886
rect 310612 262822 310664 262828
rect 310520 244928 310572 244934
rect 310520 244870 310572 244876
rect 309232 228472 309284 228478
rect 309232 228414 309284 228420
rect 309244 118658 309272 228414
rect 309324 214600 309376 214606
rect 309324 214542 309376 214548
rect 309336 133890 309364 214542
rect 309324 133884 309376 133890
rect 309324 133826 309376 133832
rect 309232 118652 309284 118658
rect 309232 118594 309284 118600
rect 310532 99346 310560 244870
rect 310624 155922 310652 262822
rect 310612 155916 310664 155922
rect 310612 155858 310664 155864
rect 311912 132462 311940 273906
rect 311992 231124 312044 231130
rect 311992 231066 312044 231072
rect 311900 132456 311952 132462
rect 311900 132398 311952 132404
rect 312004 128314 312032 231066
rect 313292 146266 313320 283834
rect 313280 146260 313332 146266
rect 313280 146202 313332 146208
rect 311992 128308 312044 128314
rect 311992 128250 312044 128256
rect 310520 99340 310572 99346
rect 310520 99282 310572 99288
rect 310520 25560 310572 25566
rect 310520 25502 310572 25508
rect 310532 16574 310560 25502
rect 311898 24168 311954 24177
rect 311898 24103 311954 24112
rect 311912 16574 311940 24103
rect 309152 16546 309824 16574
rect 310532 16546 311480 16574
rect 311912 16546 312216 16574
rect 307944 13116 307996 13122
rect 307944 13058 307996 13064
rect 307760 3528 307812 3534
rect 307760 3470 307812 3476
rect 307956 480 307984 13058
rect 309048 3528 309100 3534
rect 309048 3470 309100 3476
rect 309060 480 309088 3470
rect 309796 490 309824 16546
rect 310072 598 310284 626
rect 310072 490 310100 598
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 462 310100 490
rect 310256 480 310284 598
rect 311452 480 311480 16546
rect 312188 490 312216 16546
rect 313832 4480 313884 4486
rect 313832 4422 313884 4428
rect 312464 598 312676 626
rect 312464 490 312492 598
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 462 312492 490
rect 312648 480 312676 598
rect 313844 480 313872 4422
rect 313936 3534 313964 336767
rect 320180 313948 320232 313954
rect 320180 313890 320232 313896
rect 316038 309224 316094 309233
rect 316038 309159 316094 309168
rect 314658 282976 314714 282985
rect 314658 282911 314714 282920
rect 314014 207768 314070 207777
rect 314014 207703 314070 207712
rect 313924 3528 313976 3534
rect 313924 3470 313976 3476
rect 314028 3126 314056 207703
rect 314672 125526 314700 282911
rect 315302 196616 315358 196625
rect 315302 196551 315358 196560
rect 314660 125520 314712 125526
rect 314660 125462 314712 125468
rect 315028 3528 315080 3534
rect 315028 3470 315080 3476
rect 314016 3120 314068 3126
rect 314016 3062 314068 3068
rect 315040 480 315068 3470
rect 315316 3466 315344 196551
rect 316052 4486 316080 309159
rect 318064 306400 318116 306406
rect 318064 306342 318116 306348
rect 317420 217320 317472 217326
rect 317420 217262 317472 217268
rect 316130 195256 316186 195265
rect 316130 195191 316186 195200
rect 316144 16574 316172 195191
rect 317432 125594 317460 217262
rect 317420 125588 317472 125594
rect 317420 125530 317472 125536
rect 317420 19984 317472 19990
rect 317420 19926 317472 19932
rect 316144 16546 316264 16574
rect 316040 4480 316092 4486
rect 316040 4422 316092 4428
rect 315304 3460 315356 3466
rect 315304 3402 315356 3408
rect 316236 480 316264 16546
rect 317432 6914 317460 19926
rect 318076 15910 318104 306342
rect 318798 191040 318854 191049
rect 318798 190975 318854 190984
rect 318812 16574 318840 190975
rect 320192 16574 320220 313890
rect 321572 16574 321600 367095
rect 582378 365120 582434 365129
rect 582378 365055 582434 365064
rect 582392 349761 582420 365055
rect 582378 349752 582434 349761
rect 582378 349687 582434 349696
rect 357438 345128 357494 345137
rect 357438 345063 357494 345072
rect 336002 340912 336058 340921
rect 336002 340847 336058 340856
rect 324318 332616 324374 332625
rect 324318 332551 324374 332560
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 318064 15904 318116 15910
rect 318064 15846 318116 15852
rect 317432 6886 318104 6914
rect 317328 3120 317380 3126
rect 317328 3062 317380 3068
rect 317340 480 317368 3062
rect 318076 490 318104 6886
rect 318352 598 318564 626
rect 318352 490 318380 598
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 462 318380 490
rect 318536 480 318564 598
rect 319732 480 319760 16546
rect 320468 490 320496 16546
rect 320744 598 320956 626
rect 320744 490 320772 598
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 462 320772 490
rect 320928 480 320956 598
rect 322124 480 322152 16546
rect 324332 3534 324360 332551
rect 331220 327752 331272 327758
rect 331220 327694 331272 327700
rect 327078 313984 327134 313993
rect 327078 313919 327134 313928
rect 325700 188352 325752 188358
rect 325700 188294 325752 188300
rect 324412 40724 324464 40730
rect 324412 40666 324464 40672
rect 324320 3528 324372 3534
rect 324320 3470 324372 3476
rect 323308 3460 323360 3466
rect 323308 3402 323360 3408
rect 323320 480 323348 3402
rect 324424 480 324452 40666
rect 325712 16574 325740 188294
rect 327092 16574 327120 313919
rect 329838 182880 329894 182889
rect 329838 182815 329894 182824
rect 329852 16574 329880 182815
rect 325712 16546 326384 16574
rect 327092 16546 328040 16574
rect 329852 16546 330432 16574
rect 325608 3528 325660 3534
rect 325608 3470 325660 3476
rect 325620 480 325648 3470
rect 326356 490 326384 16546
rect 326632 598 326844 626
rect 326632 490 326660 598
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 462 326660 490
rect 326816 480 326844 598
rect 328012 480 328040 16546
rect 328736 15904 328788 15910
rect 328736 15846 328788 15852
rect 328748 490 328776 15846
rect 329024 598 329236 626
rect 329024 490 329052 598
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 328748 462 329052 490
rect 329208 480 329236 598
rect 330404 480 330432 16546
rect 331232 490 331260 327694
rect 333978 327040 334034 327049
rect 333978 326975 334034 326984
rect 332598 318064 332654 318073
rect 332598 317999 332654 318008
rect 332612 6914 332640 317999
rect 332690 208992 332746 209001
rect 332690 208927 332746 208936
rect 332704 11762 332732 208927
rect 333992 16574 334020 326975
rect 335360 189100 335412 189106
rect 335360 189042 335412 189048
rect 335372 16574 335400 189042
rect 333992 16546 334664 16574
rect 335372 16546 335952 16574
rect 332692 11756 332744 11762
rect 332692 11698 332744 11704
rect 333888 11756 333940 11762
rect 333888 11698 333940 11704
rect 332612 6886 332732 6914
rect 331416 598 331628 626
rect 331416 490 331444 598
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 462 331444 490
rect 331600 480 331628 598
rect 332704 480 332732 6886
rect 333900 480 333928 11698
rect 334636 490 334664 16546
rect 335924 3346 335952 16546
rect 336016 3534 336044 340847
rect 339498 334112 339554 334121
rect 339498 334047 339554 334056
rect 338118 311128 338174 311137
rect 338118 311063 338174 311072
rect 338132 16574 338160 311063
rect 338132 16546 338712 16574
rect 336004 3528 336056 3534
rect 336004 3470 336056 3476
rect 337476 3528 337528 3534
rect 337476 3470 337528 3476
rect 335924 3318 336320 3346
rect 334912 598 335124 626
rect 334912 490 334940 598
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 462 334940 490
rect 335096 480 335124 598
rect 336292 480 336320 3318
rect 337488 480 337516 3470
rect 338684 480 338712 16546
rect 339512 490 339540 334047
rect 349160 323604 349212 323610
rect 349160 323546 349212 323552
rect 345018 210352 345074 210361
rect 345018 210287 345074 210296
rect 340878 204912 340934 204921
rect 340878 204847 340934 204856
rect 340892 3534 340920 204847
rect 342258 184240 342314 184249
rect 342258 184175 342314 184184
rect 342272 16574 342300 184175
rect 345032 16574 345060 210287
rect 347042 57216 347098 57225
rect 347042 57151 347098 57160
rect 342272 16546 342944 16574
rect 345032 16546 345336 16574
rect 340972 6180 341024 6186
rect 340972 6122 341024 6128
rect 340880 3528 340932 3534
rect 340880 3470 340932 3476
rect 339696 598 339908 626
rect 339696 490 339724 598
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 462 339724 490
rect 339880 480 339908 598
rect 340984 480 341012 6122
rect 342168 3528 342220 3534
rect 342168 3470 342220 3476
rect 342180 480 342208 3470
rect 342916 490 342944 16546
rect 344558 3360 344614 3369
rect 344558 3295 344614 3304
rect 343192 598 343404 626
rect 343192 490 343220 598
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 462 343220 490
rect 343376 480 343404 598
rect 344572 480 344600 3295
rect 345308 490 345336 16546
rect 346952 8968 347004 8974
rect 346952 8910 347004 8916
rect 345584 598 345796 626
rect 345584 490 345612 598
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 462 345612 490
rect 345768 480 345796 598
rect 346964 480 346992 8910
rect 347056 3058 347084 57151
rect 349172 6186 349200 323546
rect 356058 222864 356114 222873
rect 356058 222799 356114 222808
rect 353298 199336 353354 199345
rect 353298 199271 353354 199280
rect 349160 6180 349212 6186
rect 349160 6122 349212 6128
rect 348054 3496 348110 3505
rect 348054 3431 348110 3440
rect 351644 3460 351696 3466
rect 347044 3052 347096 3058
rect 347044 2994 347096 3000
rect 348068 480 348096 3431
rect 351644 3402 351696 3408
rect 350448 3188 350500 3194
rect 350448 3130 350500 3136
rect 349252 3052 349304 3058
rect 349252 2994 349304 3000
rect 349264 480 349292 2994
rect 350460 480 350488 3130
rect 351656 480 351684 3402
rect 353312 3194 353340 199271
rect 356072 3369 356100 222799
rect 357452 3505 357480 345063
rect 582378 343768 582434 343777
rect 582378 343703 582434 343712
rect 565084 303680 565136 303686
rect 565084 303622 565136 303628
rect 565096 219434 565124 303622
rect 580262 298752 580318 298761
rect 580262 298687 580318 298696
rect 574744 298172 574796 298178
rect 574744 298114 574796 298120
rect 565084 219428 565136 219434
rect 565084 219370 565136 219376
rect 358818 197976 358874 197985
rect 358818 197911 358874 197920
rect 357438 3496 357494 3505
rect 358832 3466 358860 197911
rect 574756 179382 574784 298114
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 240145 580212 245511
rect 580170 240136 580226 240145
rect 580170 240071 580226 240080
rect 580276 234569 580304 298687
rect 580354 272232 580410 272241
rect 580354 272167 580410 272176
rect 580368 257378 580396 272167
rect 580356 257372 580408 257378
rect 580356 257314 580408 257320
rect 580262 234560 580318 234569
rect 580262 234495 580318 234504
rect 580908 221196 580960 221202
rect 580908 221138 580960 221144
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 574744 179376 574796 179382
rect 574744 179318 574796 179324
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580920 126041 580948 221138
rect 580906 126032 580962 126041
rect 580906 125967 580962 125976
rect 580170 90400 580226 90409
rect 580170 90335 580226 90344
rect 580184 86193 580212 90335
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 582392 16574 582420 343703
rect 582484 291825 582512 418231
rect 582562 404968 582618 404977
rect 582562 404903 582618 404912
rect 582470 291816 582526 291825
rect 582470 291751 582526 291760
rect 582576 291174 582604 404903
rect 582564 291168 582616 291174
rect 582564 291110 582616 291116
rect 582470 284336 582526 284345
rect 582470 284271 582526 284280
rect 582484 258913 582512 284271
rect 582668 276010 582696 471407
rect 582746 378448 582802 378457
rect 582746 378383 582802 378392
rect 582760 282878 582788 378383
rect 583022 351928 583078 351937
rect 583022 351863 583078 351872
rect 582838 325272 582894 325281
rect 582838 325207 582894 325216
rect 582748 282872 582800 282878
rect 582748 282814 582800 282820
rect 582656 276004 582708 276010
rect 582656 275946 582708 275952
rect 582656 268388 582708 268394
rect 582656 268330 582708 268336
rect 582470 258904 582526 258913
rect 582470 258839 582526 258848
rect 582668 232393 582696 268330
rect 582852 247722 582880 325207
rect 582930 295352 582986 295361
rect 582930 295287 582986 295296
rect 582840 247716 582892 247722
rect 582840 247658 582892 247664
rect 582838 237960 582894 237969
rect 582838 237895 582894 237904
rect 582748 235272 582800 235278
rect 582748 235214 582800 235220
rect 582654 232384 582710 232393
rect 582654 232319 582710 232328
rect 582654 225040 582710 225049
rect 582654 224975 582710 224984
rect 582392 16546 582604 16574
rect 582196 3528 582248 3534
rect 582196 3470 582248 3476
rect 357438 3431 357494 3440
rect 358820 3460 358872 3466
rect 358820 3402 358872 3408
rect 356058 3360 356114 3369
rect 356058 3295 356114 3304
rect 353300 3188 353352 3194
rect 353300 3130 353352 3136
rect 581000 3120 581052 3126
rect 581000 3062 581052 3068
rect 581012 480 581040 3062
rect 582208 480 582236 3470
rect 582576 3346 582604 16546
rect 582668 6633 582696 224975
rect 582760 33153 582788 235214
rect 582852 46345 582880 237895
rect 582944 112849 582972 295287
rect 583036 289785 583064 351863
rect 583390 312080 583446 312089
rect 583390 312015 583446 312024
rect 583206 300112 583262 300121
rect 583206 300047 583262 300056
rect 583114 292632 583170 292641
rect 583114 292567 583170 292576
rect 583022 289776 583078 289785
rect 583022 289711 583078 289720
rect 583024 265668 583076 265674
rect 583024 265610 583076 265616
rect 582930 112840 582986 112849
rect 582930 112775 582986 112784
rect 583036 99521 583064 265610
rect 583128 205737 583156 292567
rect 583114 205728 583170 205737
rect 583114 205663 583170 205672
rect 583220 139369 583248 300047
rect 583300 278044 583352 278050
rect 583300 277986 583352 277992
rect 583312 152697 583340 277986
rect 583404 270502 583432 312015
rect 583484 307828 583536 307834
rect 583484 307770 583536 307776
rect 583392 270496 583444 270502
rect 583392 270438 583444 270444
rect 583390 217288 583446 217297
rect 583390 217223 583446 217232
rect 583298 152688 583354 152697
rect 583298 152623 583354 152632
rect 583206 139360 583262 139369
rect 583206 139295 583262 139304
rect 583022 99512 583078 99521
rect 583022 99447 583078 99456
rect 582838 46336 582894 46345
rect 582838 46271 582894 46280
rect 582746 33144 582802 33153
rect 582746 33079 582802 33088
rect 582654 6624 582710 6633
rect 582654 6559 582710 6568
rect 583404 3534 583432 217223
rect 583496 193089 583524 307770
rect 583666 296848 583722 296857
rect 583666 296783 583722 296792
rect 583680 287054 583708 296783
rect 583758 293992 583814 294001
rect 583814 293950 583984 293978
rect 583758 293927 583814 293936
rect 583680 287026 583892 287054
rect 583576 279472 583628 279478
rect 583576 279414 583628 279420
rect 583588 221202 583616 279414
rect 583668 251864 583720 251870
rect 583668 251806 583720 251812
rect 583576 221196 583628 221202
rect 583576 221138 583628 221144
rect 583574 206272 583630 206281
rect 583574 206207 583630 206216
rect 583482 193080 583538 193089
rect 583482 193015 583538 193024
rect 583392 3528 583444 3534
rect 583392 3470 583444 3476
rect 582576 3318 583432 3346
rect 583404 480 583432 3318
rect 583588 3126 583616 206207
rect 583680 166433 583708 251806
rect 583758 220960 583814 220969
rect 583758 220895 583814 220904
rect 583666 166424 583722 166433
rect 583666 166359 583722 166368
rect 583772 80050 583800 220895
rect 583680 80022 583800 80050
rect 583680 70394 583708 80022
rect 583864 72826 583892 287026
rect 583852 72820 583904 72826
rect 583852 72762 583904 72768
rect 583850 72720 583906 72729
rect 583956 72706 583984 293950
rect 583906 72678 583984 72706
rect 583850 72655 583906 72664
rect 583852 72616 583904 72622
rect 583852 72558 583904 72564
rect 583680 70366 583800 70394
rect 583772 60217 583800 70366
rect 583758 60208 583814 60217
rect 583758 60143 583814 60152
rect 583864 20369 583892 72558
rect 583850 20360 583906 20369
rect 583850 20295 583906 20304
rect 583576 3120 583628 3126
rect 583576 3062 583628 3068
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3422 671200 3478 671256
rect 3514 658144 3570 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3422 579944 3478 580000
rect 3422 566888 3478 566944
rect 2778 553852 2834 553888
rect 2778 553832 2780 553852
rect 2780 553832 2832 553852
rect 2832 553832 2834 553852
rect 3422 527856 3478 527912
rect 3330 501744 3386 501800
rect 2778 462596 2834 462632
rect 2778 462576 2780 462596
rect 2780 462576 2832 462596
rect 2832 462576 2834 462596
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 4066 475632 4122 475688
rect 3146 449520 3202 449576
rect 3146 423544 3202 423600
rect 3422 410488 3478 410544
rect 2778 397432 2834 397488
rect 3422 388864 3478 388920
rect 3422 386960 3478 387016
rect 3514 371320 3570 371376
rect 3330 358400 3386 358456
rect 3146 345344 3202 345400
rect 2778 293120 2834 293176
rect 3146 254088 3202 254144
rect 7562 381520 7618 381576
rect 7562 328480 7618 328536
rect 4066 319232 4122 319288
rect 3514 306176 3570 306232
rect 3514 267144 3570 267200
rect 3514 241032 3570 241088
rect 4802 237224 4858 237280
rect 3422 214920 3478 214976
rect 3422 210296 3478 210352
rect 3054 201864 3110 201920
rect 3238 162832 3294 162888
rect 2778 149776 2834 149832
rect 3514 188808 3570 188864
rect 17222 330384 17278 330440
rect 3514 136720 3570 136776
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 12346 80688 12402 80744
rect 5446 79464 5502 79520
rect 3422 71576 3478 71632
rect 4066 68176 4122 68232
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 2870 32408 2926 32464
rect 3974 28192 4030 28248
rect 110 22616 166 22672
rect 18 6704 74 6760
rect 3422 19352 3478 19408
rect 10966 35128 11022 35184
rect 9586 10240 9642 10296
rect 17866 72392 17922 72448
rect 15106 59880 15162 59936
rect 16486 43424 16542 43480
rect 25502 293936 25558 293992
rect 29642 79328 29698 79384
rect 26146 76472 26202 76528
rect 23386 69536 23442 69592
rect 22006 50224 22062 50280
rect 24766 29552 24822 29608
rect 33046 62736 33102 62792
rect 36542 203632 36598 203688
rect 35806 66816 35862 66872
rect 34426 47504 34482 47560
rect 37186 44784 37242 44840
rect 43994 427080 44050 427136
rect 41326 75112 41382 75168
rect 41326 73752 41382 73808
rect 40682 64096 40738 64152
rect 39578 6160 39634 6216
rect 46846 26832 46902 26888
rect 52274 440816 52330 440872
rect 55034 444624 55090 444680
rect 54942 411304 54998 411360
rect 53470 387640 53526 387696
rect 52366 385600 52422 385656
rect 50894 240080 50950 240136
rect 50894 54440 50950 54496
rect 51722 224168 51778 224224
rect 52182 208256 52238 208312
rect 53838 331064 53894 331120
rect 54942 331064 54998 331120
rect 53838 330384 53894 330440
rect 53654 238448 53710 238504
rect 54942 213832 54998 213888
rect 53746 72528 53802 72584
rect 53746 55800 53802 55856
rect 56322 239944 56378 240000
rect 56414 235864 56470 235920
rect 57610 220768 57666 220824
rect 59174 445848 59230 445904
rect 58990 377304 59046 377360
rect 61934 590688 61990 590744
rect 61842 427080 61898 427136
rect 61934 366288 61990 366344
rect 60646 353912 60702 353968
rect 59082 352008 59138 352064
rect 57794 241304 57850 241360
rect 56506 65456 56562 65512
rect 60462 335416 60518 335472
rect 58990 231784 59046 231840
rect 59174 234504 59230 234560
rect 59082 212472 59138 212528
rect 57886 57160 57942 57216
rect 57886 51720 57942 51776
rect 60462 241984 60518 242040
rect 60554 216552 60610 216608
rect 61842 226208 61898 226264
rect 61934 71032 61990 71088
rect 66074 579672 66130 579728
rect 66810 588240 66866 588296
rect 66258 586508 66260 586528
rect 66260 586508 66312 586528
rect 66312 586508 66314 586528
rect 66258 586472 66314 586508
rect 66810 582412 66866 582448
rect 66810 582392 66812 582412
rect 66812 582392 66864 582412
rect 66864 582392 66866 582412
rect 66994 581052 67050 581088
rect 66994 581032 66996 581052
rect 66996 581032 67048 581052
rect 67048 581032 67050 581052
rect 66902 575592 66958 575648
rect 67454 575320 67510 575376
rect 66442 573144 66498 573200
rect 66442 571784 66498 571840
rect 67270 570152 67326 570208
rect 66810 568792 66866 568848
rect 66902 567432 66958 567488
rect 66626 564576 66682 564632
rect 66442 564032 66498 564088
rect 66442 561992 66498 562048
rect 66626 560360 66682 560416
rect 66626 559000 66682 559056
rect 66350 555192 66406 555248
rect 66258 554684 66260 554704
rect 66260 554684 66312 554704
rect 66312 554684 66314 554704
rect 66258 554648 66314 554684
rect 66534 549616 66590 549672
rect 66534 548256 66590 548312
rect 66810 547576 66866 547632
rect 66166 546352 66222 546408
rect 66810 544856 66866 544912
rect 66810 542680 66866 542736
rect 67086 541728 67142 541784
rect 65522 392572 65524 392592
rect 65524 392572 65576 392592
rect 65576 392572 65578 392592
rect 65522 392536 65578 392572
rect 64142 345616 64198 345672
rect 59266 24112 59322 24168
rect 64694 338272 64750 338328
rect 64786 331744 64842 331800
rect 65982 391040 66038 391096
rect 67546 566752 67602 566808
rect 72974 699760 73030 699816
rect 70858 590688 70914 590744
rect 72974 589328 73030 589384
rect 77942 592048 77998 592104
rect 77022 590688 77078 590744
rect 81346 595448 81402 595504
rect 82542 590960 82598 591016
rect 81438 590688 81494 590744
rect 86866 590824 86922 590880
rect 75642 588648 75698 588704
rect 88246 588784 88302 588840
rect 88062 588512 88118 588568
rect 67730 585792 67786 585848
rect 67730 578312 67786 578368
rect 67638 558864 67694 558920
rect 67362 556280 67418 556336
rect 66994 439864 67050 439920
rect 66810 437688 66866 437744
rect 66810 435240 66866 435296
rect 66902 433064 66958 433120
rect 66902 430888 66958 430944
rect 66810 428440 66866 428496
rect 66258 426264 66314 426320
rect 66258 424088 66314 424144
rect 66258 421912 66314 421968
rect 66902 417288 66958 417344
rect 66442 415148 66444 415168
rect 66444 415148 66496 415168
rect 66496 415148 66498 415168
rect 66442 415112 66498 415148
rect 66534 408312 66590 408368
rect 66626 406136 66682 406192
rect 66350 403688 66406 403744
rect 66810 401548 66812 401568
rect 66812 401548 66864 401568
rect 66864 401548 66866 401568
rect 66810 401512 66866 401548
rect 66902 399336 66958 399392
rect 66258 396888 66314 396944
rect 66166 389136 66222 389192
rect 66166 356632 66222 356688
rect 65522 314200 65578 314256
rect 65982 301416 66038 301472
rect 64510 241440 64566 241496
rect 64602 232600 64658 232656
rect 66074 275984 66130 276040
rect 66074 272040 66130 272096
rect 65890 250008 65946 250064
rect 67454 552200 67510 552256
rect 67362 419464 67418 419520
rect 67454 412664 67510 412720
rect 67362 396888 67418 396944
rect 67362 349016 67418 349072
rect 67270 341128 67326 341184
rect 66718 323720 66774 323776
rect 66626 320456 66682 320512
rect 66718 318280 66774 318336
rect 66626 309848 66682 309904
rect 66534 306856 66590 306912
rect 66718 292984 66774 293040
rect 66718 287816 66774 287872
rect 66902 324808 66958 324864
rect 67270 326984 67326 327040
rect 67178 322632 67234 322688
rect 66902 319368 66958 319424
rect 66902 317500 66904 317520
rect 66904 317500 66956 317520
rect 66956 317500 66958 317520
rect 66902 317464 66958 317500
rect 66902 313112 66958 313168
rect 66902 310936 66958 310992
rect 67086 309032 67142 309088
rect 67086 307944 67142 308000
rect 66902 305768 66958 305824
rect 66902 303628 66904 303648
rect 66904 303628 66956 303648
rect 66956 303628 66958 303648
rect 66902 303592 66958 303628
rect 66994 302504 67050 302560
rect 66902 300600 66958 300656
rect 67178 304680 67234 304736
rect 67086 299512 67142 299568
rect 66902 296248 66958 296304
rect 67086 294072 67142 294128
rect 66902 292168 66958 292224
rect 66994 291080 67050 291136
rect 66902 289992 66958 290048
rect 66902 288904 66958 288960
rect 66902 286728 66958 286784
rect 66810 285676 66812 285696
rect 66812 285676 66864 285696
rect 66864 285676 66866 285696
rect 66810 285640 66866 285676
rect 66994 284552 67050 284608
rect 66718 283736 66774 283792
rect 66350 282648 66406 282704
rect 66810 280472 66866 280528
rect 66718 278296 66774 278352
rect 67822 576952 67878 577008
rect 88890 576748 88946 576804
rect 68650 540776 68706 540832
rect 76746 539552 76802 539608
rect 68466 535472 68522 535528
rect 69662 535472 69718 535528
rect 70674 535472 70730 535528
rect 69662 458224 69718 458280
rect 67730 442040 67786 442096
rect 67546 394712 67602 394768
rect 67546 315288 67602 315344
rect 67454 309032 67510 309088
rect 67362 298424 67418 298480
rect 67546 281560 67602 281616
rect 67270 279384 67326 279440
rect 66810 275304 66866 275360
rect 66810 274216 66866 274272
rect 67086 277208 67142 277264
rect 66994 273128 67050 273184
rect 66902 270952 66958 271008
rect 66718 269864 66774 269920
rect 66258 267688 66314 267744
rect 66810 265784 66866 265840
rect 66810 264696 66866 264752
rect 66534 263608 66590 263664
rect 66442 262520 66498 262576
rect 66810 261432 66866 261488
rect 66810 260344 66866 260400
rect 66718 258440 66774 258496
rect 66902 254088 66958 254144
rect 66902 253000 66958 253056
rect 66810 248920 66866 248976
rect 66626 247832 66682 247888
rect 67270 246744 67326 246800
rect 66626 245112 66682 245168
rect 67178 242800 67234 242856
rect 66166 228248 66222 228304
rect 76194 536696 76250 536752
rect 76102 535472 76158 535528
rect 76746 535472 76802 535528
rect 76562 445984 76618 446040
rect 81438 462848 81494 462904
rect 82726 453192 82782 453248
rect 82082 452648 82138 452704
rect 84750 536016 84806 536072
rect 84106 454688 84162 454744
rect 83462 451288 83518 451344
rect 86958 458768 87014 458824
rect 86866 457408 86922 457464
rect 86222 447752 86278 447808
rect 85578 445848 85634 445904
rect 88338 456048 88394 456104
rect 88890 445712 88946 445768
rect 89902 585656 89958 585712
rect 90362 585656 90418 585712
rect 89810 560088 89866 560144
rect 91190 587016 91246 587072
rect 92110 584840 92166 584896
rect 91926 583652 91928 583672
rect 91928 583652 91980 583672
rect 91980 583652 91982 583672
rect 91926 583616 91982 583652
rect 91190 581576 91246 581632
rect 91190 578856 91246 578912
rect 91190 577496 91246 577552
rect 91926 574796 91982 574832
rect 91926 574776 91928 574796
rect 91928 574776 91980 574796
rect 91980 574776 91982 574796
rect 91098 573416 91154 573472
rect 91190 572056 91246 572112
rect 91098 571412 91100 571432
rect 91100 571412 91152 571432
rect 91152 571412 91154 571432
rect 91098 571376 91154 571412
rect 91098 570016 91154 570072
rect 91742 568656 91798 568712
rect 91098 567704 91154 567760
rect 91098 565836 91100 565856
rect 91100 565836 91152 565856
rect 91152 565836 91154 565856
rect 91098 565800 91154 565836
rect 91098 564460 91154 564496
rect 91098 564440 91100 564460
rect 91100 564440 91152 564460
rect 91152 564440 91154 564460
rect 91098 563100 91154 563136
rect 91098 563080 91100 563100
rect 91100 563080 91152 563100
rect 91152 563080 91154 563100
rect 91098 560904 91154 560960
rect 91190 558184 91246 558240
rect 91190 556824 91246 556880
rect 91190 555464 91246 555520
rect 91282 552744 91338 552800
rect 91190 552100 91192 552120
rect 91192 552100 91244 552120
rect 91244 552100 91246 552120
rect 91190 552064 91246 552100
rect 91190 549344 91246 549400
rect 91190 547848 91246 547904
rect 91282 546508 91338 546544
rect 91282 546488 91284 546508
rect 91284 546488 91336 546508
rect 91336 546488 91338 546508
rect 91282 544040 91338 544096
rect 91282 542428 91338 542464
rect 91282 542408 91284 542428
rect 91284 542408 91336 542428
rect 91336 542408 91338 542428
rect 91282 541320 91338 541376
rect 91282 539708 91338 539744
rect 91282 539688 91284 539708
rect 91284 539688 91336 539708
rect 91336 539688 91338 539708
rect 91834 560088 91890 560144
rect 91742 453192 91798 453248
rect 90132 444488 90188 444544
rect 93766 581576 93822 581632
rect 92570 545128 92626 545184
rect 92570 542952 92626 543008
rect 93122 464344 93178 464400
rect 94502 462848 94558 462904
rect 96526 465704 96582 465760
rect 94410 445712 94466 445768
rect 92478 444624 92534 444680
rect 93076 444624 93132 444680
rect 97998 592048 98054 592104
rect 97906 580896 97962 580952
rect 97906 580216 97962 580272
rect 100022 590824 100078 590880
rect 98642 588648 98698 588704
rect 100758 588784 100814 588840
rect 96618 445712 96674 445768
rect 97354 445712 97410 445768
rect 97998 445748 98000 445768
rect 98000 445748 98052 445768
rect 98052 445748 98054 445768
rect 97998 445712 98054 445748
rect 104162 462168 104218 462224
rect 104806 447752 104862 447808
rect 100942 444624 100998 444680
rect 108302 595448 108358 595504
rect 107106 590960 107162 591016
rect 108118 542952 108174 543008
rect 107014 462848 107070 462904
rect 108302 448704 108358 448760
rect 108946 447888 109002 447944
rect 111062 448568 111118 448624
rect 110418 445712 110474 445768
rect 111154 445712 111210 445768
rect 109498 444760 109554 444816
rect 116582 585656 116638 585712
rect 115386 538600 115442 538656
rect 113178 445712 113234 445768
rect 114098 445712 114154 445768
rect 118698 460128 118754 460184
rect 117318 445712 117374 445768
rect 120722 440136 120778 440192
rect 120722 434696 120778 434752
rect 120630 404232 120686 404288
rect 86222 390904 86278 390960
rect 92754 390904 92810 390960
rect 70030 390632 70086 390688
rect 68650 389000 68706 389056
rect 68834 388728 68890 388784
rect 71870 390360 71926 390416
rect 71042 355272 71098 355328
rect 70398 351872 70454 351928
rect 67730 346976 67786 347032
rect 70122 342216 70178 342272
rect 68006 328616 68062 328672
rect 70674 332696 70730 332752
rect 70030 327020 70032 327040
rect 70032 327020 70084 327040
rect 70084 327020 70086 327040
rect 70030 326984 70086 327020
rect 71686 351872 71742 351928
rect 73066 339632 73122 339688
rect 71410 334192 71466 334248
rect 80058 390360 80114 390416
rect 80610 390360 80666 390416
rect 80058 389136 80114 389192
rect 76562 362208 76618 362264
rect 77298 357992 77354 358048
rect 83554 387640 83610 387696
rect 83554 387232 83610 387288
rect 85486 378800 85542 378856
rect 80058 364928 80114 364984
rect 80058 357448 80114 357504
rect 74630 336776 74686 336832
rect 73710 334328 73766 334384
rect 77942 332560 77998 332616
rect 77298 327528 77354 327584
rect 78218 327528 78274 327584
rect 80702 340992 80758 341048
rect 82726 338680 82782 338736
rect 83002 327528 83058 327584
rect 85578 366288 85634 366344
rect 91374 390360 91430 390416
rect 89810 389000 89866 389056
rect 91006 388320 91062 388376
rect 88246 378664 88302 378720
rect 87602 363024 87658 363080
rect 86958 357448 87014 357504
rect 85762 349288 85818 349344
rect 91190 359216 91246 359272
rect 87142 337048 87198 337104
rect 88614 336912 88670 336968
rect 88430 329976 88486 330032
rect 89810 335552 89866 335608
rect 102138 390904 102194 390960
rect 95882 390360 95938 390416
rect 97354 390360 97410 390416
rect 95238 388456 95294 388512
rect 95882 386960 95938 387016
rect 97262 369824 97318 369880
rect 96526 360984 96582 361040
rect 95146 356224 95202 356280
rect 92386 332424 92442 332480
rect 78586 327256 78642 327312
rect 92846 331200 92902 331256
rect 95146 351056 95202 351112
rect 95054 330656 95110 330712
rect 97170 332832 97226 332888
rect 98826 390360 98882 390416
rect 100666 390360 100722 390416
rect 107934 390904 107990 390960
rect 114098 390904 114154 390960
rect 101126 389000 101182 389056
rect 101954 389000 102010 389056
rect 100114 364248 100170 364304
rect 104990 390360 105046 390416
rect 106554 390360 106610 390416
rect 104990 381520 105046 381576
rect 102046 367104 102102 367160
rect 101494 360168 101550 360224
rect 101954 360168 102010 360224
rect 98642 339496 98698 339552
rect 100114 331064 100170 331120
rect 99286 330520 99342 330576
rect 97814 330384 97870 330440
rect 98642 330384 98698 330440
rect 98550 330248 98606 330304
rect 115754 390632 115810 390688
rect 108026 390360 108082 390416
rect 107934 388320 107990 388376
rect 109498 390360 109554 390416
rect 105634 381520 105690 381576
rect 105542 345616 105598 345672
rect 106186 338136 106242 338192
rect 111062 361800 111118 361856
rect 109682 358944 109738 359000
rect 108946 343712 109002 343768
rect 108302 330656 108358 330712
rect 110418 353368 110474 353424
rect 110326 346568 110382 346624
rect 109682 338680 109738 338736
rect 112626 389000 112682 389056
rect 111798 354864 111854 354920
rect 111706 353368 111762 353424
rect 115110 382220 115166 382256
rect 115110 382200 115112 382220
rect 115112 382200 115164 382220
rect 115164 382200 115166 382220
rect 115938 390360 115994 390416
rect 114558 364384 114614 364440
rect 115846 364384 115902 364440
rect 111706 340856 111762 340912
rect 111890 327664 111946 327720
rect 112810 329976 112866 330032
rect 115202 347928 115258 347984
rect 120170 390360 120226 390416
rect 118698 389136 118754 389192
rect 119342 369960 119398 370016
rect 118698 350512 118754 350568
rect 120906 442720 120962 442776
rect 121182 439864 121238 439920
rect 120814 419464 120870 419520
rect 121642 453192 121698 453248
rect 121550 428440 121606 428496
rect 121550 417288 121606 417344
rect 121458 396888 121514 396944
rect 121458 392536 121514 392592
rect 120814 390632 120870 390688
rect 120722 371320 120778 371376
rect 115938 345752 115994 345808
rect 116582 342352 116638 342408
rect 117318 347656 117374 347712
rect 117318 346432 117374 346488
rect 118606 345072 118662 345128
rect 119342 350512 119398 350568
rect 121642 410488 121698 410544
rect 123114 433064 123170 433120
rect 123298 428440 123354 428496
rect 122930 424088 122986 424144
rect 123206 424088 123262 424144
rect 122746 422184 122802 422240
rect 123114 415132 123170 415168
rect 123114 415112 123116 415132
rect 123116 415112 123168 415132
rect 123168 415112 123170 415132
rect 122746 412800 122802 412856
rect 123114 412664 123170 412720
rect 122746 412528 122802 412584
rect 122746 403008 122802 403064
rect 122746 402872 122802 402928
rect 122746 393352 122802 393408
rect 122746 393216 122802 393272
rect 123022 392536 123078 392592
rect 122746 383696 122802 383752
rect 122746 383560 122802 383616
rect 122746 374040 122802 374096
rect 122746 373904 122802 373960
rect 122746 364520 122802 364576
rect 122746 364112 122802 364168
rect 121458 361664 121514 361720
rect 123390 421912 123446 421968
rect 124126 444216 124182 444272
rect 124126 442040 124182 442096
rect 123850 437688 123906 437744
rect 124126 433064 124182 433120
rect 124126 408348 124128 408368
rect 124128 408348 124180 408368
rect 124180 408348 124182 408368
rect 124126 408312 124182 408348
rect 123574 406136 123630 406192
rect 124126 401548 124128 401568
rect 124128 401548 124180 401568
rect 124180 401548 124182 401568
rect 124126 401512 124182 401548
rect 123666 399336 123722 399392
rect 124126 394712 124182 394768
rect 124862 536696 124918 536752
rect 123482 367648 123538 367704
rect 123298 360848 123354 360904
rect 122746 355272 122802 355328
rect 121366 343848 121422 343904
rect 120722 338408 120778 338464
rect 120722 330520 120778 330576
rect 122102 328752 122158 328808
rect 122930 345208 122986 345264
rect 124862 435240 124918 435296
rect 126242 444624 126298 444680
rect 125598 358808 125654 358864
rect 124310 351056 124366 351112
rect 124862 350648 124918 350704
rect 124126 346568 124182 346624
rect 123482 328480 123538 328536
rect 125322 334056 125378 334112
rect 125690 357312 125746 357368
rect 126242 357312 126298 357368
rect 125690 356088 125746 356144
rect 128450 536016 128506 536072
rect 130382 448568 130438 448624
rect 126978 360848 127034 360904
rect 126978 359352 127034 359408
rect 126978 357584 127034 357640
rect 129738 355952 129794 356008
rect 129738 354728 129794 354784
rect 154118 702480 154174 702536
rect 582378 697176 582434 697232
rect 580262 670656 580318 670712
rect 580170 590960 580226 591016
rect 135074 367240 135130 367296
rect 130474 355952 130530 356008
rect 130382 352552 130438 352608
rect 131486 329840 131542 329896
rect 137282 444488 137338 444544
rect 135902 366968 135958 367024
rect 135166 347112 135222 347168
rect 135258 335688 135314 335744
rect 135902 331744 135958 331800
rect 136914 331472 136970 331528
rect 135258 328888 135314 328944
rect 580262 577632 580318 577688
rect 579802 537784 579858 537840
rect 582470 683848 582526 683904
rect 582562 644000 582618 644056
rect 582378 536016 582434 536072
rect 582654 630808 582710 630864
rect 582746 617480 582802 617536
rect 582746 595448 582802 595504
rect 582746 564304 582802 564360
rect 582470 524456 582526 524512
rect 580170 511284 580226 511320
rect 580170 511264 580172 511284
rect 580172 511264 580224 511284
rect 580224 511264 580226 511284
rect 582378 484608 582434 484664
rect 169022 458224 169078 458280
rect 141422 369008 141478 369064
rect 138018 366968 138074 367024
rect 138018 365744 138074 365800
rect 140870 349424 140926 349480
rect 140870 346976 140926 347032
rect 140778 346568 140834 346624
rect 139306 342488 139362 342544
rect 142066 339768 142122 339824
rect 140870 331336 140926 331392
rect 139766 328616 139822 328672
rect 140870 330384 140926 330440
rect 140778 329024 140834 329080
rect 140778 328752 140834 328808
rect 140778 327800 140834 327856
rect 142894 330112 142950 330168
rect 144918 352144 144974 352200
rect 145562 352144 145618 352200
rect 150254 364248 150310 364304
rect 150254 363160 150310 363216
rect 148322 328480 148378 328536
rect 150438 363160 150494 363216
rect 153842 345616 153898 345672
rect 147218 327120 147274 327176
rect 150714 327120 150770 327176
rect 153658 327156 153660 327176
rect 153660 327156 153712 327176
rect 153712 327156 153714 327176
rect 153658 327120 153714 327156
rect 154210 327004 154266 327040
rect 154210 326984 154212 327004
rect 154212 326984 154264 327004
rect 154264 326984 154266 327004
rect 68098 326712 68154 326768
rect 68650 326440 68706 326496
rect 154854 324944 154910 325000
rect 67822 321544 67878 321600
rect 67730 312024 67786 312080
rect 154670 276936 154726 276992
rect 67638 268776 67694 268832
rect 67638 255176 67694 255232
rect 67362 239808 67418 239864
rect 67270 222808 67326 222864
rect 67178 217232 67234 217288
rect 67730 245656 67786 245712
rect 157338 364928 157394 364984
rect 156694 353912 156750 353968
rect 156234 328480 156290 328536
rect 156050 325352 156106 325408
rect 156050 324264 156106 324320
rect 156142 323176 156198 323232
rect 156050 322088 156106 322144
rect 155958 314744 156014 314800
rect 156602 321000 156658 321056
rect 156602 318552 156658 318608
rect 156142 308488 156198 308544
rect 156510 307400 156566 307456
rect 156050 304136 156106 304192
rect 156418 297880 156474 297936
rect 156326 294616 156382 294672
rect 154762 264696 154818 264752
rect 156234 288360 156290 288416
rect 156326 285096 156382 285152
rect 156510 273672 156566 273728
rect 155866 264152 155922 264208
rect 154854 261976 154910 262032
rect 68190 258712 68246 258768
rect 67914 250280 67970 250336
rect 70306 241984 70362 242040
rect 69662 241848 69718 241904
rect 67822 237088 67878 237144
rect 69662 225800 69718 225856
rect 72422 239808 72478 239864
rect 71410 238584 71466 238640
rect 70490 228384 70546 228440
rect 67638 205536 67694 205592
rect 72606 239400 72662 239456
rect 73066 197920 73122 197976
rect 75182 240080 75238 240136
rect 74722 236544 74778 236600
rect 73802 204176 73858 204232
rect 75458 240080 75514 240136
rect 76562 238448 76618 238504
rect 75826 228928 75882 228984
rect 77206 223488 77262 223544
rect 75182 199960 75238 200016
rect 82956 241304 83012 241360
rect 84106 241168 84162 241224
rect 84842 239400 84898 239456
rect 84842 225936 84898 225992
rect 84106 224848 84162 224904
rect 85486 209072 85542 209128
rect 86958 217776 87014 217832
rect 88246 196560 88302 196616
rect 79966 192480 80022 192536
rect 90914 220088 90970 220144
rect 92294 215872 92350 215928
rect 92386 209616 92442 209672
rect 93858 241304 93914 241360
rect 94364 241304 94420 241360
rect 93674 218592 93730 218648
rect 93766 191664 93822 191720
rect 95146 189624 95202 189680
rect 91006 185544 91062 185600
rect 101954 221448 102010 221504
rect 102138 231648 102194 231704
rect 102046 212336 102102 212392
rect 100666 207576 100722 207632
rect 103518 233144 103574 233200
rect 106738 231648 106794 231704
rect 108946 227160 109002 227216
rect 110326 217912 110382 217968
rect 111614 203496 111670 203552
rect 115202 232600 115258 232656
rect 115202 222128 115258 222184
rect 114466 219272 114522 219328
rect 115754 202680 115810 202736
rect 111706 200640 111762 200696
rect 107566 193840 107622 193896
rect 104162 193160 104218 193216
rect 103426 190984 103482 191040
rect 99286 188264 99342 188320
rect 97906 182960 97962 183016
rect 98918 182144 98974 182200
rect 98918 177520 98974 177576
rect 100758 179424 100814 179480
rect 116030 235592 116086 235648
rect 118652 241304 118708 241360
rect 119342 223352 119398 223408
rect 122102 233824 122158 233880
rect 122102 228792 122158 228848
rect 122654 215192 122710 215248
rect 122930 238448 122986 238504
rect 125322 233280 125378 233336
rect 124126 206896 124182 206952
rect 122746 204856 122802 204912
rect 121366 202816 121422 202872
rect 126150 239672 126206 239728
rect 126886 213696 126942 213752
rect 129554 230288 129610 230344
rect 128358 210976 128414 211032
rect 132314 214512 132370 214568
rect 133602 231648 133658 231704
rect 133510 231376 133566 231432
rect 133694 207712 133750 207768
rect 129646 202136 129702 202192
rect 135994 241984 136050 242040
rect 136914 241984 136970 242040
rect 138202 241984 138258 242040
rect 135166 227296 135222 227352
rect 136730 237224 136786 237280
rect 136730 236000 136786 236056
rect 137282 236000 137338 236056
rect 137282 224576 137338 224632
rect 136546 220632 136602 220688
rect 146758 241984 146814 242040
rect 141790 239808 141846 239864
rect 138662 233008 138718 233064
rect 140042 229744 140098 229800
rect 138662 202680 138718 202736
rect 133786 198056 133842 198112
rect 140778 233280 140834 233336
rect 140778 231512 140834 231568
rect 142342 234368 142398 234424
rect 140686 208936 140742 208992
rect 140042 201320 140098 201376
rect 138662 197240 138718 197296
rect 144918 233008 144974 233064
rect 147678 213968 147734 214024
rect 154026 241712 154082 241768
rect 149058 237224 149114 237280
rect 150530 235728 150586 235784
rect 151174 233824 151230 233880
rect 151082 232464 151138 232520
rect 151174 228792 151230 228848
rect 128266 195880 128322 195936
rect 152462 225936 152518 225992
rect 153106 210840 153162 210896
rect 155222 242936 155278 242992
rect 154854 241440 154910 241496
rect 154394 204992 154450 205048
rect 156418 258984 156474 259040
rect 156418 253580 156420 253600
rect 156420 253580 156472 253600
rect 156472 253580 156474 253600
rect 156418 253544 156474 253580
rect 156418 249464 156474 249520
rect 156050 244024 156106 244080
rect 155682 235592 155738 235648
rect 157246 319912 157302 319968
rect 157246 318844 157302 318880
rect 157246 318824 157248 318844
rect 157248 318824 157300 318844
rect 157300 318824 157302 318844
rect 157246 316920 157302 316976
rect 157246 315832 157302 315888
rect 157246 312568 157302 312624
rect 157246 311480 157302 311536
rect 157246 310392 157302 310448
rect 157154 309576 157210 309632
rect 157246 309168 157302 309224
rect 157154 308352 157210 308408
rect 157246 306332 157302 306368
rect 157246 306312 157248 306332
rect 157248 306312 157300 306332
rect 157300 306312 157302 306332
rect 157246 305244 157302 305280
rect 157246 305224 157248 305244
rect 157248 305224 157300 305244
rect 157300 305224 157302 305244
rect 156694 303592 156750 303648
rect 157246 303048 157302 303104
rect 156786 301960 156842 302016
rect 157154 300056 157210 300112
rect 157246 298968 157302 299024
rect 156694 296792 156750 296848
rect 157246 292712 157302 292768
rect 157522 292712 157578 292768
rect 156786 291624 156842 291680
rect 156694 291080 156750 291136
rect 157246 290536 157302 290592
rect 156694 290128 156750 290184
rect 156786 289448 156842 289504
rect 156694 287272 156750 287328
rect 156694 275168 156750 275224
rect 156694 259800 156750 259856
rect 156602 227432 156658 227488
rect 154486 202272 154542 202328
rect 157246 286184 157302 286240
rect 157246 284316 157248 284336
rect 157248 284316 157300 284336
rect 157300 284316 157302 284336
rect 157246 284280 157302 284316
rect 157246 283192 157302 283248
rect 157154 282104 157210 282160
rect 157246 281016 157302 281072
rect 156970 279928 157026 279984
rect 156878 276664 156934 276720
rect 157246 278840 157302 278896
rect 157246 277752 157302 277808
rect 157062 275848 157118 275904
rect 156878 274760 156934 274816
rect 157154 272584 157210 272640
rect 157246 271496 157302 271552
rect 157246 270408 157302 270464
rect 157246 268232 157302 268288
rect 157246 267416 157302 267472
rect 157246 265240 157302 265296
rect 157246 263064 157302 263120
rect 156878 257932 156880 257952
rect 156880 257932 156932 257952
rect 156932 257932 156934 257952
rect 156878 257896 156934 257932
rect 157246 256828 157302 256864
rect 157246 256808 157248 256828
rect 157248 256808 157300 256828
rect 157300 256808 157302 256828
rect 157246 255720 157302 255776
rect 157246 254632 157302 254688
rect 156786 247288 156842 247344
rect 157246 250552 157302 250608
rect 157154 248376 157210 248432
rect 156970 245112 157026 245168
rect 156878 242120 156934 242176
rect 156878 240760 156934 240816
rect 158074 307808 158130 307864
rect 157982 235184 158038 235240
rect 159546 335416 159602 335472
rect 159362 327800 159418 327856
rect 158626 295296 158682 295352
rect 159546 322088 159602 322144
rect 160190 342488 160246 342544
rect 160190 335960 160246 336016
rect 159454 291080 159510 291136
rect 159546 282104 159602 282160
rect 159362 273264 159418 273320
rect 158718 235184 158774 235240
rect 158166 227160 158222 227216
rect 156694 199280 156750 199336
rect 160006 230288 160062 230344
rect 160926 315016 160982 315072
rect 160926 289040 160982 289096
rect 162306 335688 162362 335744
rect 162122 295432 162178 295488
rect 160742 195880 160798 195936
rect 151726 195200 151782 195256
rect 115846 187584 115902 187640
rect 118514 180784 118570 180840
rect 113362 179560 113418 179616
rect 102046 177520 102102 177576
rect 106186 177520 106242 177576
rect 108946 177520 109002 177576
rect 113086 177520 113142 177576
rect 124954 180920 125010 180976
rect 121366 177520 121422 177576
rect 118514 177384 118570 177440
rect 113362 176976 113418 177032
rect 115846 176976 115902 177032
rect 117962 176976 118018 177032
rect 100758 176840 100814 176896
rect 124954 177520 125010 177576
rect 125966 177520 126022 177576
rect 128266 177520 128322 177576
rect 162306 273808 162362 273864
rect 162214 245656 162270 245712
rect 162122 237088 162178 237144
rect 161386 224712 161442 224768
rect 162398 243480 162454 243536
rect 162214 211792 162270 211848
rect 163686 328888 163742 328944
rect 163502 300192 163558 300248
rect 162858 210840 162914 210896
rect 160926 202816 160982 202872
rect 163594 280064 163650 280120
rect 163594 234368 163650 234424
rect 160834 181328 160890 181384
rect 132406 177520 132462 177576
rect 133786 177520 133842 177576
rect 148230 177520 148286 177576
rect 131026 177248 131082 177304
rect 100666 176704 100722 176760
rect 117962 176704 118018 176760
rect 121918 176704 121974 176760
rect 123298 176704 123354 176760
rect 128174 176704 128230 176760
rect 129462 176704 129518 176760
rect 136086 176724 136142 176760
rect 136086 176704 136088 176724
rect 136088 176704 136140 176724
rect 136140 176704 136142 176724
rect 158994 176740 158996 176760
rect 158996 176740 159048 176760
rect 159048 176740 159050 176760
rect 158994 176704 159050 176740
rect 66166 129240 66222 129296
rect 65522 128016 65578 128072
rect 65982 125160 66038 125216
rect 66074 122576 66130 122632
rect 67454 123528 67510 123584
rect 67362 102312 67418 102368
rect 67270 100680 67326 100736
rect 66074 82728 66130 82784
rect 163502 176568 163558 176624
rect 165066 338272 165122 338328
rect 165158 282648 165214 282704
rect 164974 269728 165030 269784
rect 166538 335552 166594 335608
rect 166262 236680 166318 236736
rect 166262 227296 166318 227352
rect 167642 352008 167698 352064
rect 167642 315288 167698 315344
rect 167642 284280 167698 284336
rect 169022 286320 169078 286376
rect 169022 275304 169078 275360
rect 168378 260888 168434 260944
rect 167826 260072 167882 260128
rect 169206 274760 169262 274816
rect 169114 249872 169170 249928
rect 164974 203632 165030 203688
rect 166262 198056 166318 198112
rect 119434 174936 119490 174992
rect 135258 174800 135314 174856
rect 167826 220632 167882 220688
rect 166354 179424 166410 179480
rect 166998 175888 167054 175944
rect 166538 175480 166594 175536
rect 167642 171536 167698 171592
rect 167826 180920 167882 180976
rect 173162 343848 173218 343904
rect 171874 338408 171930 338464
rect 170586 306448 170642 306504
rect 170402 291352 170458 291408
rect 169758 261160 169814 261216
rect 170402 246200 170458 246256
rect 169298 240760 169354 240816
rect 169758 236700 169814 236736
rect 169758 236680 169760 236700
rect 169760 236680 169812 236700
rect 169812 236680 169814 236700
rect 169114 233144 169170 233200
rect 169114 202272 169170 202328
rect 169022 176976 169078 177032
rect 67638 126248 67694 126304
rect 67730 120808 67786 120864
rect 100666 94696 100722 94752
rect 117134 93472 117190 93528
rect 121734 93472 121790 93528
rect 110142 93200 110198 93256
rect 113822 93200 113878 93256
rect 84382 92384 84438 92440
rect 89074 92384 89130 92440
rect 75366 91160 75422 91216
rect 86222 91160 86278 91216
rect 86866 91160 86922 91216
rect 88246 91160 88302 91216
rect 75366 88168 75422 88224
rect 86222 85448 86278 85504
rect 67454 78376 67510 78432
rect 74446 77832 74502 77888
rect 70214 76608 70270 76664
rect 64418 69672 64474 69728
rect 66166 61376 66222 61432
rect 68926 53080 68982 53136
rect 64326 3304 64382 3360
rect 73066 73888 73122 73944
rect 75826 64232 75882 64288
rect 81346 40568 81402 40624
rect 96342 91840 96398 91896
rect 93214 91704 93270 91760
rect 91006 91160 91062 91216
rect 91926 91160 91982 91216
rect 95146 91160 95202 91216
rect 93214 89664 93270 89720
rect 91926 88032 91982 88088
rect 96342 85312 96398 85368
rect 95146 75248 95202 75304
rect 88982 73072 89038 73128
rect 87602 62872 87658 62928
rect 86866 61512 86922 61568
rect 89626 58520 89682 58576
rect 99102 92384 99158 92440
rect 106830 92384 106886 92440
rect 99286 91704 99342 91760
rect 97906 91296 97962 91352
rect 97814 91160 97870 91216
rect 99194 91160 99250 91216
rect 102046 91296 102102 91352
rect 100022 91160 100078 91216
rect 101218 91160 101274 91216
rect 101954 91160 102010 91216
rect 99286 89528 99342 89584
rect 101218 86808 101274 86864
rect 100022 86672 100078 86728
rect 99286 82048 99342 82104
rect 101954 78512 102010 78568
rect 103426 91160 103482 91216
rect 104438 91160 104494 91216
rect 105542 91160 105598 91216
rect 106094 91160 106150 91216
rect 104162 71168 104218 71224
rect 109682 92384 109738 92440
rect 107566 91160 107622 91216
rect 108486 91160 108542 91216
rect 106922 80008 106978 80064
rect 108486 87896 108542 87952
rect 110694 92420 110696 92440
rect 110696 92420 110748 92440
rect 110748 92420 110750 92440
rect 110694 92384 110750 92420
rect 111522 92384 111578 92440
rect 110234 91160 110290 91216
rect 110234 84088 110290 84144
rect 106922 42064 106978 42120
rect 112718 91160 112774 91216
rect 114282 91296 114338 91352
rect 115754 91296 115810 91352
rect 113822 89392 113878 89448
rect 114374 91160 114430 91216
rect 115846 91160 115902 91216
rect 124126 92384 124182 92440
rect 119802 91704 119858 91760
rect 118606 91296 118662 91352
rect 118514 91160 118570 91216
rect 124034 91432 124090 91488
rect 119894 91160 119950 91216
rect 120446 91160 120502 91216
rect 120722 91160 120778 91216
rect 122746 91160 122802 91216
rect 120446 85176 120502 85232
rect 122102 65592 122158 65648
rect 124126 83408 124182 83464
rect 122102 3304 122158 3360
rect 133878 94424 133934 94480
rect 135810 93608 135866 93664
rect 135994 93608 136050 93664
rect 135994 93336 136050 93392
rect 136086 92420 136088 92440
rect 136088 92420 136140 92440
rect 136140 92420 136142 92440
rect 136086 92384 136142 92420
rect 151450 92384 151506 92440
rect 125414 91296 125470 91352
rect 126886 91296 126942 91352
rect 125506 91160 125562 91216
rect 126794 91160 126850 91216
rect 128266 91160 128322 91216
rect 129646 91160 129702 91216
rect 132406 91160 132462 91216
rect 130382 68448 130438 68504
rect 151542 91296 151598 91352
rect 150438 81368 150494 81424
rect 142802 80824 142858 80880
rect 136454 11600 136510 11656
rect 132958 8880 133014 8936
rect 125874 3304 125930 3360
rect 151634 91160 151690 91216
rect 152462 91160 152518 91216
rect 165066 90752 165122 90808
rect 166446 111968 166502 112024
rect 167826 111696 167882 111752
rect 168286 110064 168342 110120
rect 168010 108704 168066 108760
rect 167918 105440 167974 105496
rect 167642 86672 167698 86728
rect 167918 93472 167974 93528
rect 169758 189760 169814 189816
rect 169206 179560 169262 179616
rect 169206 151000 169262 151056
rect 169022 92112 169078 92168
rect 170494 182824 170550 182880
rect 170494 180784 170550 180840
rect 172426 212336 172482 212392
rect 172794 212336 172850 212392
rect 171874 191664 171930 191720
rect 173254 298152 173310 298208
rect 174634 347928 174690 347984
rect 174542 330112 174598 330168
rect 173806 239808 173862 239864
rect 173254 232736 173310 232792
rect 173254 178336 173310 178392
rect 167826 85448 167882 85504
rect 160742 68312 160798 68368
rect 170586 106800 170642 106856
rect 170586 85176 170642 85232
rect 170494 80008 170550 80064
rect 171874 84904 171930 84960
rect 173254 94424 173310 94480
rect 173162 87896 173218 87952
rect 171874 73072 171930 73128
rect 173346 85312 173402 85368
rect 176014 342352 176070 342408
rect 174634 253816 174690 253872
rect 174818 126248 174874 126304
rect 174818 89528 174874 89584
rect 176106 265104 176162 265160
rect 176014 236000 176070 236056
rect 176106 235864 176162 235920
rect 176014 198192 176070 198248
rect 177394 267824 177450 267880
rect 177394 233008 177450 233064
rect 178682 341128 178738 341184
rect 178682 330384 178738 330440
rect 178682 320728 178738 320784
rect 177946 179968 178002 180024
rect 177394 178200 177450 178256
rect 176014 116456 176070 116512
rect 176106 89392 176162 89448
rect 160742 10240 160798 10296
rect 178958 332832 179014 332888
rect 178958 249056 179014 249112
rect 179326 235864 179382 235920
rect 180154 236000 180210 236056
rect 180062 211792 180118 211848
rect 178958 182144 179014 182200
rect 180246 231240 180302 231296
rect 185582 367240 185638 367296
rect 182822 346568 182878 346624
rect 180798 270408 180854 270464
rect 181258 270408 181314 270464
rect 181258 269728 181314 269784
rect 181442 253816 181498 253872
rect 182730 239944 182786 240000
rect 181626 191120 181682 191176
rect 181534 176840 181590 176896
rect 181442 136584 181498 136640
rect 180338 94016 180394 94072
rect 181534 105440 181590 105496
rect 181442 84768 181498 84824
rect 181626 88032 181682 88088
rect 183006 291216 183062 291272
rect 184202 266328 184258 266384
rect 183006 230424 183062 230480
rect 182914 196696 182970 196752
rect 182914 115096 182970 115152
rect 182822 33768 182878 33824
rect 184478 285912 184534 285968
rect 184386 266464 184442 266520
rect 184570 279520 184626 279576
rect 184570 220768 184626 220824
rect 184294 217776 184350 217832
rect 191102 345208 191158 345264
rect 187054 339768 187110 339824
rect 189722 334328 189778 334384
rect 185674 297336 185730 297392
rect 185674 294072 185730 294128
rect 185582 178880 185638 178936
rect 185950 231512 186006 231568
rect 186226 231512 186282 231568
rect 185950 231104 186006 231160
rect 187514 249056 187570 249112
rect 187514 248512 187570 248568
rect 186962 204040 187018 204096
rect 185766 202272 185822 202328
rect 187054 193976 187110 194032
rect 186962 189624 187018 189680
rect 185766 178064 185822 178120
rect 185674 177248 185730 177304
rect 185582 21256 185638 21312
rect 184202 10240 184258 10296
rect 187698 228248 187754 228304
rect 187698 220768 187754 220824
rect 187606 198056 187662 198112
rect 187146 175208 187202 175264
rect 187054 93880 187110 93936
rect 189814 283464 189870 283520
rect 189722 244840 189778 244896
rect 191194 317328 191250 317384
rect 191654 288768 191710 288824
rect 189814 223352 189870 223408
rect 189722 216008 189778 216064
rect 188434 204856 188490 204912
rect 191102 244432 191158 244488
rect 190826 226072 190882 226128
rect 190366 189760 190422 189816
rect 189722 145560 189778 145616
rect 188526 136584 188582 136640
rect 189722 113736 189778 113792
rect 191654 228384 191710 228440
rect 191102 133048 191158 133104
rect 189906 118768 189962 118824
rect 192574 302232 192630 302288
rect 193126 302232 193182 302288
rect 193126 277888 193182 277944
rect 195334 360168 195390 360224
rect 195150 319368 195206 319424
rect 193862 272312 193918 272368
rect 192758 260888 192814 260944
rect 192482 233144 192538 233200
rect 191930 220904 191986 220960
rect 192758 228792 192814 228848
rect 192666 225800 192722 225856
rect 194046 264152 194102 264208
rect 194874 270408 194930 270464
rect 195426 291488 195482 291544
rect 195426 280064 195482 280120
rect 194414 244840 194470 244896
rect 193954 240760 194010 240816
rect 193954 215872 194010 215928
rect 194414 214512 194470 214568
rect 193954 204856 194010 204912
rect 195242 204992 195298 205048
rect 195978 255212 195980 255232
rect 195980 255212 196032 255232
rect 196032 255212 196034 255232
rect 195978 255176 196034 255212
rect 198002 349424 198058 349480
rect 196714 347792 196770 347848
rect 200762 342216 200818 342272
rect 198094 329840 198150 329896
rect 199474 322088 199530 322144
rect 198094 292848 198150 292904
rect 197358 291352 197414 291408
rect 198002 287408 198058 287464
rect 197358 283736 197414 283792
rect 197358 282376 197414 282432
rect 197358 280744 197414 280800
rect 197358 280200 197414 280256
rect 197450 279420 197452 279440
rect 197452 279420 197504 279440
rect 197504 279420 197506 279440
rect 197450 279384 197506 279420
rect 197450 278568 197506 278624
rect 197358 277888 197414 277944
rect 197358 277208 197414 277264
rect 197358 276684 197414 276720
rect 197358 276664 197360 276684
rect 197360 276664 197412 276684
rect 197412 276664 197414 276684
rect 197450 275848 197506 275904
rect 197358 273672 197414 273728
rect 197358 272856 197414 272912
rect 197542 274488 197598 274544
rect 197818 271496 197874 271552
rect 197358 270952 197414 271008
rect 197358 270136 197414 270192
rect 197450 269320 197506 269376
rect 197358 268776 197414 268832
rect 197358 265784 197414 265840
rect 196714 264424 196770 264480
rect 197358 263628 197414 263664
rect 197358 263608 197360 263628
rect 197360 263608 197412 263628
rect 197412 263608 197414 263628
rect 197358 263064 197414 263120
rect 197450 260072 197506 260128
rect 197358 258712 197414 258768
rect 198002 267144 198058 267200
rect 198554 282920 198610 282976
rect 200118 301280 200174 301336
rect 200762 301280 200818 301336
rect 199382 294480 199438 294536
rect 198738 287272 198794 287328
rect 199474 287136 199530 287192
rect 198738 283464 198794 283520
rect 198646 278024 198702 278080
rect 198646 274488 198702 274544
rect 198094 262248 198150 262304
rect 197358 257896 197414 257952
rect 197358 255720 197414 255776
rect 197358 254360 197414 254416
rect 197450 253544 197506 253600
rect 197358 253000 197414 253056
rect 197358 252184 197414 252240
rect 197450 251640 197506 251696
rect 197358 250824 197414 250880
rect 197358 249464 197414 249520
rect 197450 247832 197506 247888
rect 197358 245928 197414 245984
rect 197358 245148 197360 245168
rect 197360 245148 197412 245168
rect 197412 245148 197414 245168
rect 197358 245112 197414 245148
rect 196714 243752 196770 243808
rect 196622 235592 196678 235648
rect 195886 229064 195942 229120
rect 197266 242120 197322 242176
rect 196714 224576 196770 224632
rect 196622 221448 196678 221504
rect 196254 212472 196310 212528
rect 196254 211792 196310 211848
rect 191194 88984 191250 89040
rect 193862 15816 193918 15872
rect 188342 12960 188398 13016
rect 178682 4800 178738 4856
rect 198646 256536 198702 256592
rect 198094 241712 198150 241768
rect 197358 241576 197414 241632
rect 197358 213968 197414 214024
rect 197266 211792 197322 211848
rect 196714 198192 196770 198248
rect 196714 189624 196770 189680
rect 198002 181464 198058 181520
rect 197358 177928 197414 177984
rect 196806 86808 196862 86864
rect 198646 241304 198702 241360
rect 198738 231920 198794 231976
rect 198738 202408 198794 202464
rect 199566 285640 199622 285696
rect 200026 284552 200082 284608
rect 199658 284416 199714 284472
rect 582654 471416 582710 471472
rect 582470 458088 582526 458144
rect 582378 431568 582434 431624
rect 582470 418240 582526 418296
rect 204258 361800 204314 361856
rect 202786 329024 202842 329080
rect 201498 295976 201554 296032
rect 201406 291488 201462 291544
rect 202234 288496 202290 288552
rect 202234 285640 202290 285696
rect 206282 352144 206338 352200
rect 203154 288768 203210 288824
rect 203706 287136 203762 287192
rect 204258 284280 204314 284336
rect 206282 295296 206338 295352
rect 206098 287408 206154 287464
rect 207662 334192 207718 334248
rect 206650 295296 206706 295352
rect 205362 283872 205418 283928
rect 208490 332696 208546 332752
rect 207110 283872 207166 283928
rect 209134 339632 209190 339688
rect 209134 298288 209190 298344
rect 209410 298288 209466 298344
rect 209042 287136 209098 287192
rect 210422 295976 210478 296032
rect 210422 289720 210478 289776
rect 212906 327256 212962 327312
rect 211894 315288 211950 315344
rect 210882 285912 210938 285968
rect 211986 287136 212042 287192
rect 211986 284552 212042 284608
rect 212354 284280 212410 284336
rect 214654 351056 214710 351112
rect 213182 291760 213238 291816
rect 213182 286320 213238 286376
rect 215298 298016 215354 298072
rect 215298 296928 215354 296984
rect 218242 365880 218298 365936
rect 216034 337048 216090 337104
rect 215850 311888 215906 311944
rect 217322 331200 217378 331256
rect 216034 311888 216090 311944
rect 215942 298016 215998 298072
rect 217874 291252 217876 291272
rect 217876 291252 217928 291272
rect 217928 291252 217930 291272
rect 217874 291216 217930 291252
rect 216770 288632 216826 288688
rect 218058 291216 218114 291272
rect 217322 284416 217378 284472
rect 227442 364384 227498 364440
rect 220174 336912 220230 336968
rect 222842 338136 222898 338192
rect 220174 304952 220230 305008
rect 222106 304952 222162 305008
rect 218702 296792 218758 296848
rect 219162 285912 219218 285968
rect 220082 285640 220138 285696
rect 222474 289584 222530 289640
rect 222474 288632 222530 288688
rect 223946 349152 224002 349208
rect 223026 289584 223082 289640
rect 223026 287272 223082 287328
rect 226430 331336 226486 331392
rect 225418 295432 225474 295488
rect 225602 295432 225658 295488
rect 225326 292576 225382 292632
rect 208674 283872 208730 283928
rect 214102 283872 214158 283928
rect 215942 283872 215998 283928
rect 217414 283872 217470 283928
rect 225050 285776 225106 285832
rect 225970 294480 226026 294536
rect 226522 286048 226578 286104
rect 238022 363024 238078 363080
rect 232502 361664 232558 361720
rect 228362 358944 228418 359000
rect 227626 310528 227682 310584
rect 224682 283872 224738 283928
rect 226614 283872 226670 283928
rect 228362 292576 228418 292632
rect 230386 330384 230442 330440
rect 229742 295432 229798 295488
rect 229742 287408 229798 287464
rect 227994 283872 228050 283928
rect 230570 285912 230626 285968
rect 230478 284416 230534 284472
rect 233882 356088 233938 356144
rect 233698 296792 233754 296848
rect 232778 291352 232834 291408
rect 229466 283872 229522 283928
rect 231674 284416 231730 284472
rect 233882 292576 233938 292632
rect 233698 291080 233754 291136
rect 235170 302368 235226 302424
rect 235998 285640 236054 285696
rect 239402 335960 239458 336016
rect 238022 293936 238078 293992
rect 239034 293936 239090 293992
rect 239494 289992 239550 290048
rect 239954 287272 240010 287328
rect 240874 300736 240930 300792
rect 241518 300736 241574 300792
rect 240874 300056 240930 300112
rect 241426 294072 241482 294128
rect 231582 283872 231638 283928
rect 236734 283872 236790 283928
rect 242254 285776 242310 285832
rect 243450 285776 243506 285832
rect 243634 284008 243690 284064
rect 200026 282648 200082 282704
rect 199566 273808 199622 273864
rect 244094 284008 244150 284064
rect 244094 282920 244150 282976
rect 244278 278024 244334 278080
rect 244002 271224 244058 271280
rect 199474 249736 199530 249792
rect 244370 259528 244426 259584
rect 245842 300192 245898 300248
rect 245750 276684 245806 276720
rect 245750 276664 245752 276684
rect 245752 276664 245804 276684
rect 245804 276664 245806 276684
rect 247222 292712 247278 292768
rect 247130 290128 247186 290184
rect 245934 282376 245990 282432
rect 245934 281016 245990 281072
rect 245934 279384 245990 279440
rect 245934 277480 245990 277536
rect 245934 275848 245990 275904
rect 245658 274488 245714 274544
rect 245842 274488 245898 274544
rect 245842 273672 245898 273728
rect 245750 273128 245806 273184
rect 245934 272312 245990 272368
rect 245842 271516 245898 271552
rect 245842 271496 245844 271516
rect 245844 271496 245896 271516
rect 245896 271496 245898 271516
rect 245934 270136 245990 270192
rect 246394 283192 246450 283248
rect 246118 281560 246174 281616
rect 246118 280200 246174 280256
rect 246486 272312 246542 272368
rect 246026 269592 246082 269648
rect 244922 269048 244978 269104
rect 245750 267960 245806 268016
rect 245842 267416 245898 267472
rect 245934 266600 245990 266656
rect 245934 265804 245990 265840
rect 245934 265784 245936 265804
rect 245936 265784 245988 265804
rect 245988 265784 245990 265804
rect 246670 269048 246726 269104
rect 246578 265240 246634 265296
rect 244922 264152 244978 264208
rect 244462 258712 244518 258768
rect 200026 257388 200028 257408
rect 200028 257388 200080 257408
rect 200080 257388 200082 257408
rect 200026 257352 200082 257388
rect 199934 240760 199990 240816
rect 199566 240216 199622 240272
rect 244278 250824 244334 250880
rect 200210 238720 200266 238776
rect 200118 238584 200174 238640
rect 200210 237360 200266 237416
rect 201130 240080 201186 240136
rect 200762 237360 200818 237416
rect 200854 232600 200910 232656
rect 202050 237224 202106 237280
rect 201590 231104 201646 231160
rect 201498 204176 201554 204232
rect 202234 204176 202290 204232
rect 200762 178880 200818 178936
rect 198094 178608 198150 178664
rect 198094 177112 198150 177168
rect 198094 105168 198150 105224
rect 198002 39208 198058 39264
rect 196622 3304 196678 3360
rect 199474 90888 199530 90944
rect 202786 236700 202842 236736
rect 202786 236680 202788 236700
rect 202788 236680 202840 236700
rect 202840 236680 202842 236700
rect 204442 239944 204498 240000
rect 204166 239400 204222 239456
rect 205086 236680 205142 236736
rect 203614 228248 203670 228304
rect 203522 223488 203578 223544
rect 202602 198736 202658 198792
rect 202234 195336 202290 195392
rect 203522 186904 203578 186960
rect 204902 221992 204958 222048
rect 204902 220904 204958 220960
rect 205086 228384 205142 228440
rect 205362 221992 205418 222048
rect 206282 216008 206338 216064
rect 206466 211928 206522 211984
rect 206374 210976 206430 211032
rect 207386 205536 207442 205592
rect 208306 239400 208362 239456
rect 208306 238584 208362 238640
rect 208858 234368 208914 234424
rect 209042 224168 209098 224224
rect 209226 231376 209282 231432
rect 210330 235592 210386 235648
rect 210698 224168 210754 224224
rect 209778 220904 209834 220960
rect 209134 219272 209190 219328
rect 209778 213832 209834 213888
rect 210422 213152 210478 213208
rect 209134 211792 209190 211848
rect 206282 188400 206338 188456
rect 211250 209616 211306 209672
rect 211250 208392 211306 208448
rect 212170 224984 212226 225040
rect 212170 222128 212226 222184
rect 211894 208392 211950 208448
rect 213642 238584 213698 238640
rect 213090 237360 213146 237416
rect 213734 234640 213790 234696
rect 212722 202408 212778 202464
rect 215114 240080 215170 240136
rect 214562 238312 214618 238368
rect 214838 213832 214894 213888
rect 207754 175344 207810 175400
rect 207662 167048 207718 167104
rect 207754 165688 207810 165744
rect 204902 97824 204958 97880
rect 216034 237224 216090 237280
rect 216586 234368 216642 234424
rect 217322 231784 217378 231840
rect 217046 212336 217102 212392
rect 217046 211112 217102 211168
rect 217230 189896 217286 189952
rect 215942 188536 215998 188592
rect 213918 175616 213974 175672
rect 213918 174936 213974 174992
rect 214010 174256 214066 174312
rect 213918 173576 213974 173632
rect 214010 172896 214066 172952
rect 213918 172216 213974 172272
rect 214562 175208 214618 175264
rect 214102 171536 214158 171592
rect 213918 171012 213974 171048
rect 213918 170992 213920 171012
rect 213920 170992 213972 171012
rect 213972 170992 213974 171012
rect 214010 170312 214066 170368
rect 213918 169652 213974 169688
rect 213918 169632 213920 169652
rect 213920 169632 213972 169652
rect 213972 169632 213974 169652
rect 214010 168952 214066 169008
rect 213918 168308 213920 168328
rect 213920 168308 213972 168328
rect 213972 168308 213974 168328
rect 213918 168272 213974 168308
rect 213918 166948 213920 166968
rect 213920 166948 213972 166968
rect 213972 166948 213974 166968
rect 213918 166912 213974 166948
rect 214010 166368 214066 166424
rect 213918 165008 213974 165064
rect 214010 164328 214066 164384
rect 213918 163648 213974 163704
rect 214010 162968 214066 163024
rect 213918 162288 213974 162344
rect 214010 161744 214066 161800
rect 213918 161064 213974 161120
rect 214010 160384 214066 160440
rect 213918 159704 213974 159760
rect 214010 159024 214066 159080
rect 213918 158344 213974 158400
rect 214010 157664 214066 157720
rect 213918 157120 213974 157176
rect 214010 156440 214066 156496
rect 213918 155760 213974 155816
rect 214010 155080 214066 155136
rect 214010 154400 214066 154456
rect 213918 153720 213974 153776
rect 213182 153040 213238 153096
rect 207754 145560 207810 145616
rect 205086 115096 205142 115152
rect 204994 84088 205050 84144
rect 205178 84904 205234 84960
rect 207754 93064 207810 93120
rect 207662 78512 207718 78568
rect 209134 91704 209190 91760
rect 209318 91568 209374 91624
rect 209226 89664 209282 89720
rect 210606 106800 210662 106856
rect 211802 93744 211858 93800
rect 213918 152496 213974 152552
rect 214102 151136 214158 151192
rect 213918 150492 213920 150512
rect 213920 150492 213972 150512
rect 213972 150492 213974 150512
rect 213918 150456 213974 150492
rect 213918 149776 213974 149832
rect 214010 149096 214066 149152
rect 214654 151816 214710 151872
rect 214654 151000 214710 151056
rect 214562 148416 214618 148472
rect 213918 147872 213974 147928
rect 213918 147192 213974 147248
rect 216126 146512 216182 146568
rect 214010 145832 214066 145888
rect 213918 145152 213974 145208
rect 214010 144472 214066 144528
rect 213918 143792 213974 143848
rect 214010 143248 214066 143304
rect 213918 142568 213974 142624
rect 213918 141888 213974 141944
rect 214010 141208 214066 141264
rect 213918 140528 213974 140584
rect 213918 139168 213974 139224
rect 213918 137264 213974 137320
rect 214102 139848 214158 139904
rect 214654 138624 214710 138680
rect 214010 135904 214066 135960
rect 213918 135260 213920 135280
rect 213920 135260 213972 135280
rect 213972 135260 213974 135280
rect 213918 135224 213974 135260
rect 214562 134544 214618 134600
rect 213918 133900 213920 133920
rect 213920 133900 213972 133920
rect 213972 133900 213974 133920
rect 213918 133864 213974 133900
rect 214010 133320 214066 133376
rect 213274 133048 213330 133104
rect 213918 132640 213974 132696
rect 214010 131960 214066 132016
rect 213918 131280 213974 131336
rect 214010 130600 214066 130656
rect 213918 129920 213974 129976
rect 213918 129240 213974 129296
rect 214010 128696 214066 128752
rect 214010 128016 214066 128072
rect 213918 127336 213974 127392
rect 214010 126248 214066 126304
rect 213918 125976 213974 126032
rect 214562 125296 214618 125352
rect 213918 124616 213974 124672
rect 214010 124072 214066 124128
rect 213918 123392 213974 123448
rect 213918 122712 213974 122768
rect 213366 122032 213422 122088
rect 214010 121352 214066 121408
rect 213918 120672 213974 120728
rect 214010 119992 214066 120048
rect 213918 119448 213974 119504
rect 214010 118088 214066 118144
rect 213918 117428 213974 117464
rect 213918 117408 213920 117428
rect 213920 117408 213972 117428
rect 213972 117408 213974 117428
rect 214010 116728 214066 116784
rect 213918 116068 213974 116104
rect 213918 116048 213920 116068
rect 213920 116048 213972 116068
rect 213972 116048 213974 116068
rect 214562 116456 214618 116512
rect 214010 115368 214066 115424
rect 213918 114824 213974 114880
rect 213918 114144 213974 114200
rect 214286 113464 214342 113520
rect 213918 112784 213974 112840
rect 214010 111424 214066 111480
rect 213918 110744 213974 110800
rect 214010 110200 214066 110256
rect 213918 109520 213974 109576
rect 214010 108840 214066 108896
rect 213918 108160 213974 108216
rect 214010 107480 214066 107536
rect 213918 106800 213974 106856
rect 214010 106120 214066 106176
rect 213918 104932 213920 104952
rect 213920 104932 213972 104952
rect 213972 104932 213974 104952
rect 213918 104896 213974 104932
rect 214010 104216 214066 104272
rect 213918 103556 213974 103592
rect 213918 103536 213920 103556
rect 213920 103536 213972 103556
rect 213972 103536 213974 103556
rect 213458 102176 213514 102232
rect 211986 91024 212042 91080
rect 213274 87488 213330 87544
rect 214194 101496 214250 101552
rect 213918 100952 213974 101008
rect 214010 100272 214066 100328
rect 213918 99592 213974 99648
rect 214102 98912 214158 98968
rect 213918 98232 213974 98288
rect 213918 97552 213974 97608
rect 214010 96328 214066 96384
rect 214470 97824 214526 97880
rect 214194 95784 214250 95840
rect 214010 88168 214066 88224
rect 213458 82728 213514 82784
rect 213274 71168 213330 71224
rect 216034 137944 216090 138000
rect 215942 136584 215998 136640
rect 214746 126656 214802 126712
rect 215942 113736 215998 113792
rect 214746 96872 214802 96928
rect 211802 6160 211858 6216
rect 215942 93200 215998 93256
rect 216218 94424 216274 94480
rect 216126 93608 216182 93664
rect 216034 92248 216090 92304
rect 217506 212336 217562 212392
rect 219530 238584 219586 238640
rect 219530 217912 219586 217968
rect 218794 216552 218850 216608
rect 218058 208256 218114 208312
rect 218058 207032 218114 207088
rect 218702 207032 218758 207088
rect 218702 181600 218758 181656
rect 217322 177384 217378 177440
rect 221094 240080 221150 240136
rect 221922 232736 221978 232792
rect 221370 232600 221426 232656
rect 221554 232464 221610 232520
rect 220266 213696 220322 213752
rect 220266 211112 220322 211168
rect 222106 231104 222162 231160
rect 221554 197240 221610 197296
rect 222106 187584 222162 187640
rect 220726 187040 220782 187096
rect 220266 179424 220322 179480
rect 224958 240116 224960 240136
rect 224960 240116 225012 240136
rect 225012 240116 225014 240136
rect 224958 240080 225014 240116
rect 225234 237088 225290 237144
rect 226706 238448 226762 238504
rect 225694 227432 225750 227488
rect 225602 226072 225658 226128
rect 224958 215192 225014 215248
rect 224958 214784 225014 214840
rect 225694 214784 225750 214840
rect 225602 202272 225658 202328
rect 224406 199960 224462 200016
rect 228730 239672 228786 239728
rect 229006 239672 229062 239728
rect 228178 233144 228234 233200
rect 229742 240080 229798 240136
rect 226982 211792 227038 211848
rect 225878 204992 225934 205048
rect 226338 196016 226394 196072
rect 225694 193976 225750 194032
rect 225878 193976 225934 194032
rect 225602 184320 225658 184376
rect 225694 180104 225750 180160
rect 228454 196016 228510 196072
rect 228362 189760 228418 189816
rect 227718 177384 227774 177440
rect 224958 177248 225014 177304
rect 226982 177248 227038 177304
rect 220266 176568 220322 176624
rect 222934 176568 222990 176624
rect 227718 176160 227774 176216
rect 228454 176024 228510 176080
rect 229098 175072 229154 175128
rect 229098 173712 229154 173768
rect 229282 174936 229338 174992
rect 230570 240080 230626 240136
rect 230570 237360 230626 237416
rect 231766 237904 231822 237960
rect 231674 237360 231730 237416
rect 231490 231240 231546 231296
rect 230202 219136 230258 219192
rect 229742 176704 229798 176760
rect 229374 167592 229430 167648
rect 229190 164328 229246 164384
rect 232594 224712 232650 224768
rect 231766 196016 231822 196072
rect 231766 175888 231822 175944
rect 231766 175208 231822 175264
rect 231122 174664 231178 174720
rect 231766 173168 231822 173224
rect 231582 172760 231638 172816
rect 231766 171808 231822 171864
rect 231582 171400 231638 171456
rect 230110 162152 230166 162208
rect 229742 148144 229798 148200
rect 229098 146784 229154 146840
rect 229742 138352 229798 138408
rect 219254 95920 219310 95976
rect 219162 95784 219218 95840
rect 216218 51720 216274 51776
rect 226982 95920 227038 95976
rect 224222 91840 224278 91896
rect 220174 86128 220230 86184
rect 221462 50360 221518 50416
rect 220082 6160 220138 6216
rect 224406 79464 224462 79520
rect 225602 26832 225658 26888
rect 227718 95260 227774 95296
rect 227718 95240 227720 95260
rect 227720 95240 227772 95260
rect 227772 95240 227774 95260
rect 227074 50224 227130 50280
rect 229834 120400 229890 120456
rect 230478 151544 230534 151600
rect 230294 149232 230350 149288
rect 230570 149096 230626 149152
rect 230386 148008 230442 148064
rect 230294 138760 230350 138816
rect 230110 138216 230166 138272
rect 231122 170856 231178 170912
rect 230754 166096 230810 166152
rect 230754 162016 230810 162072
rect 230754 159024 230810 159080
rect 231490 164736 231546 164792
rect 231766 168952 231822 169008
rect 233514 233824 233570 233880
rect 235906 238584 235962 238640
rect 235354 238312 235410 238368
rect 236458 235728 236514 235784
rect 234986 226208 235042 226264
rect 237930 240080 237986 240136
rect 238022 239400 238078 239456
rect 237378 228792 237434 228848
rect 237378 227704 237434 227760
rect 232962 193160 233018 193216
rect 232042 175072 232098 175128
rect 231950 170448 232006 170504
rect 231766 168000 231822 168056
rect 231766 166676 231768 166696
rect 231768 166676 231820 166696
rect 231820 166676 231822 166696
rect 231766 166640 231822 166676
rect 231766 163784 231822 163840
rect 231674 162832 231730 162888
rect 231122 162424 231178 162480
rect 231306 161880 231362 161936
rect 231766 160928 231822 160984
rect 230938 160520 230994 160576
rect 231766 159568 231822 159624
rect 231766 158616 231822 158672
rect 231214 158072 231270 158128
rect 231490 157936 231546 157992
rect 230846 157664 230902 157720
rect 230938 156168 230994 156224
rect 230846 155216 230902 155272
rect 231306 153856 231362 153912
rect 230846 153720 230902 153776
rect 230662 147736 230718 147792
rect 231674 157392 231730 157448
rect 231674 154264 231730 154320
rect 231490 152904 231546 152960
rect 232594 162832 232650 162888
rect 231766 150592 231822 150648
rect 231582 150048 231638 150104
rect 231674 149640 231730 149696
rect 230846 145832 230902 145888
rect 230570 142024 230626 142080
rect 230938 135360 230994 135416
rect 230478 131144 230534 131200
rect 230938 132096 230994 132152
rect 231766 148688 231822 148744
rect 231674 144880 231730 144936
rect 231766 143928 231822 143984
rect 231766 143384 231822 143440
rect 231766 143248 231822 143304
rect 231766 142432 231822 142488
rect 231766 140700 231768 140720
rect 231768 140700 231820 140720
rect 231820 140700 231822 140720
rect 231766 140664 231822 140700
rect 231766 137844 231768 137864
rect 231768 137844 231820 137864
rect 231820 137844 231822 137864
rect 231766 137808 231822 137844
rect 231490 136856 231546 136912
rect 231766 136312 231822 136368
rect 231674 135904 231730 135960
rect 231766 134952 231822 135008
rect 231674 134408 231730 134464
rect 231306 134000 231362 134056
rect 231490 133048 231546 133104
rect 231214 132504 231270 132560
rect 231306 130328 231362 130384
rect 231122 130192 231178 130248
rect 230754 128968 230810 129024
rect 230662 127336 230718 127392
rect 230754 126928 230810 126984
rect 231214 126248 231270 126304
rect 230754 122168 230810 122224
rect 230662 118904 230718 118960
rect 230938 123120 230994 123176
rect 230846 116048 230902 116104
rect 231766 130600 231822 130656
rect 231490 129784 231546 129840
rect 231766 129240 231822 129296
rect 231490 128832 231546 128888
rect 231766 128308 231822 128344
rect 231766 128288 231768 128308
rect 231768 128288 231820 128308
rect 231820 128288 231822 128308
rect 231674 127880 231730 127936
rect 231766 125976 231822 126032
rect 232502 125976 232558 126032
rect 231306 125024 231362 125080
rect 231766 123528 231822 123584
rect 231582 121624 231638 121680
rect 231766 121216 231822 121272
rect 231214 120672 231270 120728
rect 231674 120264 231730 120320
rect 231766 119312 231822 119368
rect 231122 114552 231178 114608
rect 230846 113736 230902 113792
rect 230570 113600 230626 113656
rect 230754 110744 230810 110800
rect 231398 117952 231454 118008
rect 231490 117408 231546 117464
rect 231766 117000 231822 117056
rect 231674 116456 231730 116512
rect 231490 115096 231546 115152
rect 231766 114144 231822 114200
rect 231490 113192 231546 113248
rect 231766 112648 231822 112704
rect 231398 112240 231454 112296
rect 231214 111288 231270 111344
rect 231490 111016 231546 111072
rect 231490 109792 231546 109848
rect 230846 109384 230902 109440
rect 231306 107072 231362 107128
rect 231766 110372 231768 110392
rect 231768 110372 231820 110392
rect 231820 110372 231822 110392
rect 231766 110336 231822 110372
rect 230478 106120 230534 106176
rect 231214 105440 231270 105496
rect 231122 103672 231178 103728
rect 230570 101768 230626 101824
rect 230570 100408 230626 100464
rect 230478 97008 230534 97064
rect 230570 96192 230626 96248
rect 231122 99456 231178 99512
rect 231122 98504 231178 98560
rect 231398 105576 231454 105632
rect 231766 108432 231822 108488
rect 231582 107888 231638 107944
rect 231766 106528 231822 106584
rect 231766 105168 231822 105224
rect 231766 104216 231822 104272
rect 231766 102720 231822 102776
rect 231398 102312 231454 102368
rect 231766 102040 231822 102096
rect 231766 101360 231822 101416
rect 231674 100816 231730 100872
rect 231306 99864 231362 99920
rect 231766 97552 231822 97608
rect 231674 96600 231730 96656
rect 227074 7520 227130 7576
rect 232686 154944 232742 155000
rect 233422 180104 233478 180160
rect 233514 176024 233570 176080
rect 233330 155896 233386 155952
rect 232778 126384 232834 126440
rect 232870 124480 232926 124536
rect 232778 121760 232834 121816
rect 232686 109656 232742 109712
rect 232502 35128 232558 35184
rect 233882 118360 233938 118416
rect 233882 116184 233938 116240
rect 234802 177248 234858 177304
rect 234710 165688 234766 165744
rect 234894 168680 234950 168736
rect 234802 157392 234858 157448
rect 234158 125432 234214 125488
rect 234158 117816 234214 117872
rect 233974 103944 234030 104000
rect 235262 114824 235318 114880
rect 235446 124616 235502 124672
rect 235354 98640 235410 98696
rect 236182 178744 236238 178800
rect 236090 169496 236146 169552
rect 237378 210840 237434 210896
rect 236734 198736 236790 198792
rect 236642 176024 236698 176080
rect 236182 163376 236238 163432
rect 238114 227704 238170 227760
rect 239218 239944 239274 240000
rect 238942 236544 238998 236600
rect 238114 187176 238170 187232
rect 237470 169904 237526 169960
rect 236918 150048 236974 150104
rect 238022 119040 238078 119096
rect 236918 100000 236974 100056
rect 238298 146376 238354 146432
rect 238850 153720 238906 153776
rect 238758 153312 238814 153368
rect 240874 239808 240930 239864
rect 239770 224848 239826 224904
rect 240138 213288 240194 213344
rect 239034 173848 239090 173904
rect 238942 141072 238998 141128
rect 239402 137128 239458 137184
rect 240230 204176 240286 204232
rect 242162 238584 242218 238640
rect 241610 237360 241666 237416
rect 242162 237360 242218 237416
rect 240874 206896 240930 206952
rect 240966 204176 241022 204232
rect 241426 187720 241482 187776
rect 240874 172760 240930 172816
rect 239586 153176 239642 153232
rect 239494 112104 239550 112160
rect 239586 111696 239642 111752
rect 241426 172352 241482 172408
rect 240874 155216 240930 155272
rect 240782 126248 240838 126304
rect 239586 106800 239642 106856
rect 239494 68312 239550 68368
rect 239310 6160 239366 6216
rect 200854 1944 200910 2000
rect 242806 238448 242862 238504
rect 242714 235864 242770 235920
rect 244002 243208 244058 243264
rect 244002 241304 244058 241360
rect 244002 239808 244058 239864
rect 243726 228248 243782 228304
rect 242438 187720 242494 187776
rect 242162 101088 242218 101144
rect 241058 93200 241114 93256
rect 244462 247288 244518 247344
rect 244370 240760 244426 240816
rect 244462 230288 244518 230344
rect 244278 205128 244334 205184
rect 243726 175888 243782 175944
rect 245842 263064 245898 263120
rect 245014 258712 245070 258768
rect 245658 256536 245714 256592
rect 245658 253000 245714 253056
rect 245658 250280 245714 250336
rect 245750 248648 245806 248704
rect 245658 245112 245714 245168
rect 244462 176024 244518 176080
rect 244278 172216 244334 172272
rect 244922 171536 244978 171592
rect 243634 111152 243690 111208
rect 245106 167048 245162 167104
rect 245014 131416 245070 131472
rect 243818 123120 243874 123176
rect 243818 82048 243874 82104
rect 243726 80824 243782 80880
rect 245106 128968 245162 129024
rect 245106 102176 245162 102232
rect 245014 55800 245070 55856
rect 244922 44784 244978 44840
rect 244278 33768 244334 33824
rect 245934 262268 245990 262304
rect 245934 262248 245936 262268
rect 245936 262248 245988 262268
rect 245988 262248 245990 262268
rect 246394 260888 246450 260944
rect 245934 260072 245990 260128
rect 245934 258168 245990 258224
rect 246946 255992 247002 256048
rect 247130 257352 247186 257408
rect 246946 255176 247002 255232
rect 245934 253852 245936 253872
rect 245936 253852 245988 253872
rect 245988 253852 245990 253872
rect 245934 253816 245990 253852
rect 245934 252184 245990 252240
rect 246026 251640 246082 251696
rect 245934 248104 245990 248160
rect 245934 245928 245990 245984
rect 245934 243752 245990 243808
rect 246394 242392 246450 242448
rect 245842 222944 245898 223000
rect 247130 244568 247186 244624
rect 245658 141616 245714 141672
rect 245842 179424 245898 179480
rect 245842 157936 245898 157992
rect 247222 175888 247278 175944
rect 247130 167184 247186 167240
rect 246394 139712 246450 139768
rect 246486 127336 246542 127392
rect 245198 94424 245254 94480
rect 259458 360848 259514 360904
rect 252558 353368 252614 353424
rect 249890 307808 249946 307864
rect 248602 283736 248658 283792
rect 248510 261704 248566 261760
rect 249798 287408 249854 287464
rect 248602 236544 248658 236600
rect 247682 135360 247738 135416
rect 246486 87488 246542 87544
rect 246578 76472 246634 76528
rect 247682 61512 247738 61568
rect 248694 220768 248750 220824
rect 249154 173984 249210 174040
rect 249982 265648 250038 265704
rect 251270 296928 251326 296984
rect 249982 162016 250038 162072
rect 249798 157120 249854 157176
rect 250442 156440 250498 156496
rect 246394 47504 246450 47560
rect 249338 142432 249394 142488
rect 249246 109792 249302 109848
rect 253938 303592 253994 303648
rect 251362 173168 251418 173224
rect 251178 144744 251234 144800
rect 250442 115776 250498 115832
rect 250442 113192 250498 113248
rect 249154 66816 249210 66872
rect 244094 10240 244150 10296
rect 242898 4936 242954 4992
rect 247590 3440 247646 3496
rect 246394 3304 246450 3360
rect 250626 111968 250682 112024
rect 251914 157936 251970 157992
rect 251822 124072 251878 124128
rect 252098 144064 252154 144120
rect 251914 107888 251970 107944
rect 254030 292848 254086 292904
rect 253294 168408 253350 168464
rect 253202 160384 253258 160440
rect 252834 142976 252890 143032
rect 254122 291216 254178 291272
rect 253938 159976 253994 160032
rect 256698 316104 256754 316160
rect 255502 254088 255558 254144
rect 255410 238312 255466 238368
rect 255410 237904 255466 237960
rect 256146 174256 256202 174312
rect 255318 168544 255374 168600
rect 255962 161744 256018 161800
rect 253202 119992 253258 120048
rect 252098 108976 252154 109032
rect 253202 92520 253258 92576
rect 253386 109656 253442 109712
rect 253294 83408 253350 83464
rect 253386 64096 253442 64152
rect 254674 110336 254730 110392
rect 254858 129920 254914 129976
rect 254858 92520 254914 92576
rect 256882 298152 256938 298208
rect 257342 209072 257398 209128
rect 256054 106256 256110 106312
rect 255962 76608 256018 76664
rect 256330 107752 256386 107808
rect 256238 105440 256294 105496
rect 256054 73888 256110 73944
rect 255318 71032 255374 71088
rect 252374 3440 252430 3496
rect 254674 1944 254730 2000
rect 262218 358808 262274 358864
rect 260102 301008 260158 301064
rect 258722 160248 258778 160304
rect 257618 130328 257674 130384
rect 258814 139984 258870 140040
rect 258814 122984 258870 123040
rect 258078 114688 258134 114744
rect 258078 110336 258134 110392
rect 257526 100000 257582 100056
rect 257434 64232 257490 64288
rect 258814 75248 258870 75304
rect 263598 351872 263654 351928
rect 262862 302232 262918 302288
rect 262218 240080 262274 240136
rect 260194 237224 260250 237280
rect 267738 346432 267794 346488
rect 267002 310528 267058 310584
rect 262862 181464 262918 181520
rect 260286 170176 260342 170232
rect 260194 151272 260250 151328
rect 260194 111016 260250 111072
rect 260194 105168 260250 105224
rect 259090 80688 259146 80744
rect 262862 147736 262918 147792
rect 261482 113736 261538 113792
rect 260286 77832 260342 77888
rect 262770 133184 262826 133240
rect 262770 132776 262826 132832
rect 262770 127608 262826 127664
rect 262770 127200 262826 127256
rect 261758 109792 261814 109848
rect 263230 161472 263286 161528
rect 262862 99592 262918 99648
rect 262862 95920 262918 95976
rect 262218 69672 262274 69728
rect 261666 69536 261722 69592
rect 261574 62736 261630 62792
rect 259458 21256 259514 21312
rect 269762 298288 269818 298344
rect 266358 179424 266414 179480
rect 267094 179424 267150 179480
rect 266358 177928 266414 177984
rect 269854 286048 269910 286104
rect 269762 185544 269818 185600
rect 276662 211792 276718 211848
rect 276018 201320 276074 201376
rect 274546 178880 274602 178936
rect 273902 178744 273958 178800
rect 276754 201320 276810 201376
rect 278134 198056 278190 198112
rect 276754 177384 276810 177440
rect 278134 177248 278190 177304
rect 278870 176976 278926 177032
rect 273350 175888 273406 175944
rect 278778 175924 278780 175944
rect 278780 175924 278832 175944
rect 278832 175924 278834 175944
rect 278778 175888 278834 175924
rect 264978 175616 265034 175672
rect 265070 175208 265126 175264
rect 264978 174800 265034 174856
rect 265070 173576 265126 173632
rect 264978 172644 265034 172680
rect 264978 172624 264980 172644
rect 264980 172624 265032 172644
rect 265032 172624 265034 172644
rect 265070 172216 265126 172272
rect 264978 171400 265034 171456
rect 265070 170992 265126 171048
rect 264978 170040 265034 170096
rect 265070 169632 265126 169688
rect 264978 169224 265034 169280
rect 265162 168816 265218 168872
rect 264978 167864 265034 167920
rect 265070 167456 265126 167512
rect 264978 166640 265034 166696
rect 265070 165280 265126 165336
rect 264978 164464 265034 164520
rect 265070 164056 265126 164112
rect 264978 163648 265034 163704
rect 264518 163240 264574 163296
rect 264334 156304 264390 156360
rect 264242 128424 264298 128480
rect 263138 72392 263194 72448
rect 262954 61376 263010 61432
rect 264426 146920 264482 146976
rect 264334 110744 264390 110800
rect 264978 162288 265034 162344
rect 265346 166232 265402 166288
rect 265714 165824 265770 165880
rect 265622 164872 265678 164928
rect 264978 161064 265034 161120
rect 265070 159704 265126 159760
rect 264978 159296 265034 159352
rect 265162 158888 265218 158944
rect 265070 158072 265126 158128
rect 264978 157664 265034 157720
rect 265254 158480 265310 158536
rect 265162 157936 265218 157992
rect 264978 157120 265034 157176
rect 265070 155896 265126 155952
rect 264978 154572 264980 154592
rect 264980 154572 265032 154592
rect 265032 154572 265034 154592
rect 264978 154536 265034 154572
rect 265346 154128 265402 154184
rect 265162 153720 265218 153776
rect 265070 152904 265126 152960
rect 264978 151952 265034 152008
rect 264978 151136 265034 151192
rect 264978 149912 265034 149968
rect 265254 152496 265310 152552
rect 264978 148960 265034 149016
rect 265070 148552 265126 148608
rect 264978 147328 265034 147384
rect 280250 186904 280306 186960
rect 279330 185680 279386 185736
rect 279422 174392 279478 174448
rect 279330 170584 279386 170640
rect 280066 164872 280122 164928
rect 279330 161336 279386 161392
rect 279330 155896 279386 155952
rect 267094 155488 267150 155544
rect 265346 150728 265402 150784
rect 265070 145968 265126 146024
rect 264978 145152 265034 145208
rect 265070 144744 265126 144800
rect 264978 144336 265034 144392
rect 265898 149504 265954 149560
rect 265346 144064 265402 144120
rect 265162 143792 265218 143848
rect 265070 143384 265126 143440
rect 264978 142180 265034 142216
rect 264978 142160 264980 142180
rect 264980 142160 265032 142180
rect 265032 142160 265034 142180
rect 264978 141752 265034 141808
rect 265254 142976 265310 143032
rect 265162 141344 265218 141400
rect 265070 141208 265126 141264
rect 264978 139576 265034 139632
rect 265162 140800 265218 140856
rect 265070 138896 265126 138952
rect 265806 138624 265862 138680
rect 264978 138216 265034 138272
rect 265070 137808 265126 137864
rect 264978 136992 265034 137048
rect 264978 136176 265034 136232
rect 265070 134816 265126 134872
rect 264978 134000 265034 134056
rect 265622 134136 265678 134192
rect 265070 132232 265126 132288
rect 264978 131824 265034 131880
rect 264978 130464 265034 130520
rect 264978 129240 265034 129296
rect 265162 128832 265218 128888
rect 265070 126248 265126 126304
rect 264978 125840 265034 125896
rect 265070 125296 265126 125352
rect 264978 124480 265034 124536
rect 264978 124072 265034 124128
rect 264518 122712 264574 122768
rect 264978 122304 265034 122360
rect 264610 121488 264666 121544
rect 264426 104760 264482 104816
rect 264426 102584 264482 102640
rect 264978 120264 265034 120320
rect 264978 119720 265034 119776
rect 265438 118904 265494 118960
rect 265070 118088 265126 118144
rect 264978 117680 265034 117736
rect 265070 116728 265126 116784
rect 264978 115948 264980 115968
rect 264980 115948 265032 115968
rect 265032 115948 265034 115968
rect 264978 115912 265034 115948
rect 264978 115504 265034 115560
rect 264978 114144 265034 114200
rect 264978 112512 265034 112568
rect 264978 111560 265034 111616
rect 265070 111152 265126 111208
rect 265070 110336 265126 110392
rect 264978 109520 265034 109576
rect 265070 108976 265126 109032
rect 264978 108568 265034 108624
rect 264978 107344 265034 107400
rect 265070 106936 265126 106992
rect 264978 105984 265034 106040
rect 265070 105576 265126 105632
rect 264978 103808 265034 103864
rect 264978 103400 265034 103456
rect 265162 102992 265218 103048
rect 264978 101768 265034 101824
rect 264978 100408 265034 100464
rect 265070 100000 265126 100056
rect 265070 99184 265126 99240
rect 264978 98640 265034 98696
rect 264978 97824 265034 97880
rect 265070 97416 265126 97472
rect 264610 84768 264666 84824
rect 264426 73752 264482 73808
rect 265714 132640 265770 132696
rect 265898 134408 265954 134464
rect 267002 117136 267058 117192
rect 265898 97008 265954 97064
rect 265898 79328 265954 79384
rect 265714 65592 265770 65648
rect 265622 62872 265678 62928
rect 264242 42064 264298 42120
rect 267094 104760 267150 104816
rect 280342 179968 280398 180024
rect 281630 179424 281686 179480
rect 280434 178880 280490 178936
rect 280342 174664 280398 174720
rect 281538 169360 281594 169416
rect 281538 151816 281594 151872
rect 280250 150320 280306 150376
rect 282182 179968 282238 180024
rect 282458 172488 282514 172544
rect 282090 171672 282146 171728
rect 282826 170856 282882 170912
rect 282826 168680 282882 168736
rect 282826 167048 282882 167104
rect 282826 166368 282882 166424
rect 281998 165572 282054 165608
rect 281998 165552 282000 165572
rect 282000 165552 282052 165572
rect 282052 165552 282054 165572
rect 282826 164056 282882 164112
rect 282458 163240 282514 163296
rect 282826 162560 282882 162616
rect 282826 161744 282882 161800
rect 284298 287136 284354 287192
rect 283102 215872 283158 215928
rect 282826 160248 282882 160304
rect 281906 159432 281962 159488
rect 282366 158752 282422 158808
rect 282090 157936 282146 157992
rect 281814 156440 281870 156496
rect 282274 154944 282330 155000
rect 282826 154128 282882 154184
rect 282274 153448 282330 153504
rect 281722 152632 281778 152688
rect 281906 151136 281962 151192
rect 282642 148824 282698 148880
rect 282826 148008 282882 148064
rect 282826 147328 282882 147384
rect 282274 146512 282330 146568
rect 282826 145832 282882 145888
rect 282734 145016 282790 145072
rect 282826 144200 282882 144256
rect 282826 142704 282882 142760
rect 282550 142060 282552 142080
rect 282552 142060 282604 142080
rect 282604 142060 282606 142080
rect 282550 142024 282606 142060
rect 282826 141208 282882 141264
rect 282826 139712 282882 139768
rect 281538 138896 281594 138952
rect 281538 138216 281594 138272
rect 282826 137436 282828 137456
rect 282828 137436 282880 137456
rect 282880 137436 282882 137456
rect 282826 137400 282882 137436
rect 282826 136604 282882 136640
rect 282826 136584 282828 136604
rect 282828 136584 282880 136604
rect 282880 136584 282882 136604
rect 282826 132776 282882 132832
rect 282826 132096 282882 132152
rect 282274 130600 282330 130656
rect 280158 129784 280214 129840
rect 282090 128968 282146 129024
rect 282826 128288 282882 128344
rect 281998 127472 282054 127528
rect 279330 126248 279386 126304
rect 267646 123664 267702 123720
rect 282274 125976 282330 126032
rect 282826 125160 282882 125216
rect 282734 124480 282790 124536
rect 282826 123664 282882 123720
rect 282274 122984 282330 123040
rect 283102 135088 283158 135144
rect 267738 109928 267794 109984
rect 261758 12960 261814 13016
rect 260654 3984 260710 4040
rect 265346 4800 265402 4856
rect 278778 95784 278834 95840
rect 270498 93064 270554 93120
rect 282826 122168 282882 122224
rect 282826 121388 282828 121408
rect 282828 121388 282880 121408
rect 282880 121388 282882 121408
rect 282826 121352 282882 121388
rect 282826 120672 282882 120728
rect 282826 119856 282882 119912
rect 282734 119176 282790 119232
rect 282826 118360 282882 118416
rect 282274 117544 282330 117600
rect 282826 116048 282882 116104
rect 282826 115368 282882 115424
rect 282366 114552 282422 114608
rect 282090 113736 282146 113792
rect 282458 113076 282514 113112
rect 282458 113056 282460 113076
rect 282460 113056 282512 113076
rect 282512 113056 282514 113076
rect 282826 112240 282882 112296
rect 281722 111596 281724 111616
rect 281724 111596 281776 111616
rect 281776 111596 281778 111616
rect 281722 111560 281778 111596
rect 284390 196696 284446 196752
rect 282826 110744 282882 110800
rect 282826 109928 282882 109984
rect 282274 109248 282330 109304
rect 282826 108432 282882 108488
rect 282366 107752 282422 107808
rect 282826 105440 282882 105496
rect 281538 104624 281594 104680
rect 279330 98096 279386 98152
rect 279330 95104 279386 95160
rect 282826 103944 282882 104000
rect 282826 103128 282882 103184
rect 286322 186904 286378 186960
rect 285954 184320 286010 184376
rect 289818 229064 289874 229120
rect 288714 177248 288770 177304
rect 290002 213152 290058 213208
rect 290094 179968 290150 180024
rect 291382 214512 291438 214568
rect 291474 178744 291530 178800
rect 281722 101632 281778 101688
rect 281630 100816 281686 100872
rect 281722 100136 281778 100192
rect 282826 99340 282882 99376
rect 282826 99320 282828 99340
rect 282828 99320 282880 99340
rect 282880 99320 282882 99340
rect 282826 97860 282828 97880
rect 282828 97860 282880 97880
rect 282880 97860 282882 97880
rect 282826 97824 282882 97860
rect 282182 97008 282238 97064
rect 280158 88984 280214 89040
rect 279054 86808 279110 86864
rect 269762 15816 269818 15872
rect 269670 14456 269726 14512
rect 268382 11600 268438 11656
rect 278778 72528 278834 72584
rect 276018 66952 276074 67008
rect 276110 39208 276166 39264
rect 278318 6160 278374 6216
rect 281446 8880 281502 8936
rect 284298 75112 284354 75168
rect 286598 3440 286654 3496
rect 287794 3440 287850 3496
rect 288990 3440 289046 3496
rect 298098 304952 298154 305008
rect 296902 193976 296958 194032
rect 299570 302368 299626 302424
rect 299478 220088 299534 220144
rect 291382 3440 291438 3496
rect 294878 3304 294934 3360
rect 298466 7520 298522 7576
rect 299662 192480 299718 192536
rect 300858 207576 300914 207632
rect 304262 300872 304318 300928
rect 303618 188264 303674 188320
rect 300766 3440 300822 3496
rect 299754 3304 299810 3360
rect 306470 203496 306526 203552
rect 304998 6160 305054 6216
rect 321558 367104 321614 367160
rect 313922 336776 313978 336832
rect 309138 319368 309194 319424
rect 307758 231104 307814 231160
rect 307758 65456 307814 65512
rect 311898 24112 311954 24168
rect 316038 309168 316094 309224
rect 314658 282920 314714 282976
rect 314014 207712 314070 207768
rect 315302 196560 315358 196616
rect 316130 195200 316186 195256
rect 318798 190984 318854 191040
rect 582378 365064 582434 365120
rect 582378 349696 582434 349752
rect 357438 345072 357494 345128
rect 336002 340856 336058 340912
rect 324318 332560 324374 332616
rect 327078 313928 327134 313984
rect 329838 182824 329894 182880
rect 333978 326984 334034 327040
rect 332598 318008 332654 318064
rect 332690 208936 332746 208992
rect 339498 334056 339554 334112
rect 338118 311072 338174 311128
rect 345018 210296 345074 210352
rect 340878 204856 340934 204912
rect 342258 184184 342314 184240
rect 347042 57160 347098 57216
rect 344558 3304 344614 3360
rect 356058 222808 356114 222864
rect 353298 199280 353354 199336
rect 348054 3440 348110 3496
rect 582378 343712 582434 343768
rect 580262 298696 580318 298752
rect 358818 197920 358874 197976
rect 357438 3440 357494 3496
rect 580170 245520 580226 245576
rect 580170 240080 580226 240136
rect 580354 272176 580410 272232
rect 580262 234504 580318 234560
rect 580170 219000 580226 219056
rect 580170 179152 580226 179208
rect 580906 125976 580962 126032
rect 580170 90344 580226 90400
rect 580170 86128 580226 86184
rect 582562 404912 582618 404968
rect 582470 291760 582526 291816
rect 582470 284280 582526 284336
rect 582746 378392 582802 378448
rect 583022 351872 583078 351928
rect 582838 325216 582894 325272
rect 582470 258848 582526 258904
rect 582930 295296 582986 295352
rect 582838 237904 582894 237960
rect 582654 232328 582710 232384
rect 582654 224984 582710 225040
rect 356058 3304 356114 3360
rect 583390 312024 583446 312080
rect 583206 300056 583262 300112
rect 583114 292576 583170 292632
rect 583022 289720 583078 289776
rect 582930 112784 582986 112840
rect 583114 205672 583170 205728
rect 583390 217232 583446 217288
rect 583298 152632 583354 152688
rect 583206 139304 583262 139360
rect 583022 99456 583078 99512
rect 582838 46280 582894 46336
rect 582746 33088 582802 33144
rect 582654 6568 582710 6624
rect 583666 296792 583722 296848
rect 583758 293936 583814 293992
rect 583574 206216 583630 206272
rect 583482 193024 583538 193080
rect 583758 220904 583814 220960
rect 583666 166368 583722 166424
rect 583850 72664 583906 72720
rect 583758 60152 583814 60208
rect 583850 20304 583906 20360
<< metal3 >>
rect 69606 702476 69612 702540
rect 69676 702538 69682 702540
rect 154113 702538 154179 702541
rect 69676 702536 154179 702538
rect 69676 702480 154118 702536
rect 154174 702480 154179 702536
rect 69676 702478 154179 702480
rect 69676 702476 69682 702478
rect 154113 702475 154179 702478
rect 72969 699818 73035 699821
rect 76046 699818 76052 699820
rect 72969 699816 76052 699818
rect 72969 699760 72974 699816
rect 73030 699760 76052 699816
rect 72969 699758 76052 699760
rect 72969 699755 73035 699758
rect 76046 699756 76052 699758
rect 76116 699756 76122 699820
rect -960 697220 480 697460
rect 582373 697234 582439 697237
rect 583520 697234 584960 697324
rect 582373 697232 584960 697234
rect 582373 697176 582378 697232
rect 582434 697176 584960 697232
rect 582373 697174 584960 697176
rect 582373 697171 582439 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 582465 683906 582531 683909
rect 583520 683906 584960 683996
rect 582465 683904 584960 683906
rect 582465 683848 582470 683904
rect 582526 683848 584960 683904
rect 582465 683846 584960 683848
rect 582465 683843 582531 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3417 671258 3483 671261
rect -960 671256 3483 671258
rect -960 671200 3422 671256
rect 3478 671200 3483 671256
rect -960 671198 3483 671200
rect -960 671108 480 671198
rect 3417 671195 3483 671198
rect 580257 670714 580323 670717
rect 583520 670714 584960 670804
rect 580257 670712 584960 670714
rect 580257 670656 580262 670712
rect 580318 670656 584960 670712
rect 580257 670654 584960 670656
rect 580257 670651 580323 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3509 658202 3575 658205
rect -960 658200 3575 658202
rect -960 658144 3514 658200
rect 3570 658144 3575 658200
rect -960 658142 3575 658144
rect -960 658052 480 658142
rect 3509 658139 3575 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 582557 644058 582623 644061
rect 583520 644058 584960 644148
rect 582557 644056 584960 644058
rect 582557 644000 582562 644056
rect 582618 644000 584960 644056
rect 582557 643998 584960 644000
rect 582557 643995 582623 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 582649 630866 582715 630869
rect 583520 630866 584960 630956
rect 582649 630864 584960 630866
rect 582649 630808 582654 630864
rect 582710 630808 584960 630864
rect 582649 630806 584960 630808
rect 582649 630803 582715 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 582741 617538 582807 617541
rect 583520 617538 584960 617628
rect 582741 617536 584960 617538
rect 582741 617480 582746 617536
rect 582802 617480 584960 617536
rect 582741 617478 584960 617480
rect 582741 617475 582807 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect 81341 595506 81407 595509
rect 108297 595506 108363 595509
rect 582741 595506 582807 595509
rect 81341 595504 582807 595506
rect 81341 595448 81346 595504
rect 81402 595448 108302 595504
rect 108358 595448 582746 595504
rect 582802 595448 582807 595504
rect 81341 595446 582807 595448
rect 81341 595443 81407 595446
rect 108297 595443 108363 595446
rect 582741 595443 582807 595446
rect -960 592908 480 593148
rect 77937 592106 78003 592109
rect 97993 592106 98059 592109
rect 77937 592104 98059 592106
rect 77937 592048 77942 592104
rect 77998 592048 97998 592104
rect 98054 592048 98059 592104
rect 77937 592046 98059 592048
rect 77937 592043 78003 592046
rect 97993 592043 98059 592046
rect 82537 591018 82603 591021
rect 107101 591018 107167 591021
rect 82537 591016 107167 591018
rect 82537 590960 82542 591016
rect 82598 590960 107106 591016
rect 107162 590960 107167 591016
rect 82537 590958 107167 590960
rect 82537 590955 82603 590958
rect 107101 590955 107167 590958
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 86861 590882 86927 590885
rect 100017 590882 100083 590885
rect 86861 590880 100083 590882
rect 86861 590824 86866 590880
rect 86922 590824 100022 590880
rect 100078 590824 100083 590880
rect 583520 590868 584960 590958
rect 86861 590822 100083 590824
rect 86861 590819 86927 590822
rect 100017 590819 100083 590822
rect 61929 590746 61995 590749
rect 70853 590746 70919 590749
rect 61929 590744 70919 590746
rect 61929 590688 61934 590744
rect 61990 590688 70858 590744
rect 70914 590688 70919 590744
rect 61929 590686 70919 590688
rect 61929 590683 61995 590686
rect 70853 590683 70919 590686
rect 77017 590746 77083 590749
rect 81433 590746 81499 590749
rect 77017 590744 81499 590746
rect 77017 590688 77022 590744
rect 77078 590688 81438 590744
rect 81494 590688 81499 590744
rect 77017 590686 81499 590688
rect 77017 590683 77083 590686
rect 81433 590683 81499 590686
rect 93894 589522 93900 589524
rect 80010 589462 93900 589522
rect 72969 589386 73035 589389
rect 80010 589386 80070 589462
rect 93894 589460 93900 589462
rect 93964 589460 93970 589524
rect 72969 589384 80070 589386
rect 72969 589328 72974 589384
rect 73030 589328 80070 589384
rect 72969 589326 80070 589328
rect 72969 589323 73035 589326
rect 88241 588842 88307 588845
rect 100753 588842 100819 588845
rect 88241 588840 100819 588842
rect 88241 588784 88246 588840
rect 88302 588784 100758 588840
rect 100814 588784 100819 588840
rect 88241 588782 100819 588784
rect 88241 588779 88307 588782
rect 100753 588779 100819 588782
rect 75637 588706 75703 588709
rect 98637 588706 98703 588709
rect 75637 588704 98703 588706
rect 75637 588648 75642 588704
rect 75698 588648 98642 588704
rect 98698 588648 98703 588704
rect 75637 588646 98703 588648
rect 75637 588643 75703 588646
rect 98637 588643 98703 588646
rect 88057 588570 88123 588573
rect 88190 588570 88196 588572
rect 88057 588568 88196 588570
rect 88057 588512 88062 588568
rect 88118 588512 88196 588568
rect 88057 588510 88196 588512
rect 88057 588507 88123 588510
rect 88190 588508 88196 588510
rect 88260 588508 88266 588572
rect 66805 588298 66871 588301
rect 68878 588298 68938 588472
rect 66805 588296 68938 588298
rect 66805 588240 66810 588296
rect 66866 588240 68938 588296
rect 66805 588238 68938 588240
rect 66805 588235 66871 588238
rect 66253 586530 66319 586533
rect 66253 586528 66362 586530
rect 66253 586472 66258 586528
rect 66314 586472 66362 586528
rect 66253 586467 66362 586472
rect 66302 586394 66362 586467
rect 68878 586394 68938 587112
rect 88566 587074 88626 587656
rect 91185 587074 91251 587077
rect 88566 587072 91251 587074
rect 88566 587016 91190 587072
rect 91246 587016 91251 587072
rect 88566 587014 91251 587016
rect 91185 587011 91251 587014
rect 66302 586334 68938 586394
rect 67725 585850 67791 585853
rect 67725 585848 68938 585850
rect 67725 585792 67730 585848
rect 67786 585792 68938 585848
rect 67725 585790 68938 585792
rect 67725 585787 67791 585790
rect 68878 585752 68938 585790
rect 88566 585714 88626 586296
rect 89897 585714 89963 585717
rect 88566 585712 89963 585714
rect 88566 585656 89902 585712
rect 89958 585656 89963 585712
rect 88566 585654 89963 585656
rect 89897 585651 89963 585654
rect 90357 585714 90423 585717
rect 116577 585714 116643 585717
rect 90357 585712 116643 585714
rect 90357 585656 90362 585712
rect 90418 585656 116582 585712
rect 116638 585656 116643 585712
rect 90357 585654 116643 585656
rect 90357 585651 90423 585654
rect 116577 585651 116643 585654
rect 88566 584898 88626 584936
rect 92105 584898 92171 584901
rect 88566 584896 92171 584898
rect 88566 584840 92110 584896
rect 92166 584840 92171 584896
rect 88566 584838 92171 584840
rect 92105 584835 92171 584838
rect 67766 583748 67772 583812
rect 67836 583810 67842 583812
rect 68878 583810 68938 584392
rect 67836 583750 68938 583810
rect 67836 583748 67842 583750
rect 91921 583674 91987 583677
rect 88566 583672 91987 583674
rect 88566 583616 91926 583672
rect 91982 583616 91987 583672
rect 88566 583614 91987 583616
rect 88566 583576 88626 583614
rect 91921 583611 91987 583614
rect 66805 582450 66871 582453
rect 68878 582450 68938 583032
rect 66805 582448 68938 582450
rect 66805 582392 66810 582448
rect 66866 582392 68938 582448
rect 66805 582390 68938 582392
rect 66805 582387 66871 582390
rect 69422 582252 69428 582316
rect 69492 582252 69498 582316
rect 66989 581090 67055 581093
rect 69430 581090 69490 582252
rect 88566 581634 88626 582216
rect 91185 581634 91251 581637
rect 88566 581632 91251 581634
rect 88566 581576 91190 581632
rect 91246 581576 91251 581632
rect 88566 581574 91251 581576
rect 91185 581571 91251 581574
rect 93761 581634 93827 581637
rect 122966 581634 122972 581636
rect 93761 581632 122972 581634
rect 93761 581576 93766 581632
rect 93822 581576 122972 581632
rect 93761 581574 122972 581576
rect 93761 581571 93827 581574
rect 122966 581572 122972 581574
rect 123036 581572 123042 581636
rect 66989 581088 69490 581090
rect 66989 581032 66994 581088
rect 67050 581032 69490 581088
rect 66989 581030 69490 581032
rect 66989 581027 67055 581030
rect 97901 580954 97967 580957
rect 88566 580952 97967 580954
rect 88566 580896 97906 580952
rect 97962 580896 97967 580952
rect 88566 580894 97967 580896
rect 88566 580856 88626 580894
rect 97901 580891 97967 580894
rect -960 580002 480 580092
rect 3417 580002 3483 580005
rect -960 580000 3483 580002
rect -960 579944 3422 580000
rect 3478 579944 3483 580000
rect -960 579942 3483 579944
rect -960 579852 480 579942
rect 3417 579939 3483 579942
rect 66069 579730 66135 579733
rect 68878 579730 68938 580312
rect 97901 580274 97967 580277
rect 119470 580274 119476 580276
rect 97901 580272 119476 580274
rect 97901 580216 97906 580272
rect 97962 580216 119476 580272
rect 97901 580214 119476 580216
rect 97901 580211 97967 580214
rect 119470 580212 119476 580214
rect 119540 580212 119546 580276
rect 66069 579728 68938 579730
rect 66069 579672 66074 579728
rect 66130 579672 68938 579728
rect 66069 579670 68938 579672
rect 66069 579667 66135 579670
rect 67725 578370 67791 578373
rect 68878 578370 68938 578952
rect 88566 578914 88626 579496
rect 91185 578914 91251 578917
rect 88566 578912 91251 578914
rect 88566 578856 91190 578912
rect 91246 578856 91251 578912
rect 88566 578854 91251 578856
rect 91185 578851 91251 578854
rect 67725 578368 68938 578370
rect 67725 578312 67730 578368
rect 67786 578312 68938 578368
rect 67725 578310 68938 578312
rect 67725 578307 67791 578310
rect 67817 577010 67883 577013
rect 68878 577010 68938 577592
rect 88566 577554 88626 578136
rect 580257 577690 580323 577693
rect 583520 577690 584960 577780
rect 580257 577688 584960 577690
rect 580257 577632 580262 577688
rect 580318 577632 584960 577688
rect 580257 577630 584960 577632
rect 580257 577627 580323 577630
rect 91185 577554 91251 577557
rect 88566 577552 91251 577554
rect 88566 577496 91190 577552
rect 91246 577496 91251 577552
rect 583520 577540 584960 577630
rect 88566 577494 91251 577496
rect 91185 577491 91251 577494
rect 67817 577008 68938 577010
rect 67817 576952 67822 577008
rect 67878 576952 68938 577008
rect 67817 576950 68938 576952
rect 67817 576947 67883 576950
rect 88885 576806 88951 576809
rect 88596 576804 88951 576806
rect 88596 576748 88890 576804
rect 88946 576748 88951 576804
rect 88596 576746 88951 576748
rect 88885 576743 88951 576746
rect 66897 575650 66963 575653
rect 68878 575650 68938 576232
rect 66897 575648 68938 575650
rect 66897 575592 66902 575648
rect 66958 575592 68938 575648
rect 66897 575590 68938 575592
rect 66897 575587 66963 575590
rect 67449 575378 67515 575381
rect 67449 575376 68938 575378
rect 67449 575320 67454 575376
rect 67510 575320 68938 575376
rect 67449 575318 68938 575320
rect 67449 575315 67515 575318
rect 68878 574872 68938 575318
rect 88566 574834 88626 575416
rect 91921 574834 91987 574837
rect 88566 574832 91987 574834
rect 88566 574776 91926 574832
rect 91982 574776 91987 574832
rect 88566 574774 91987 574776
rect 91921 574771 91987 574774
rect 66437 573202 66503 573205
rect 68878 573202 68938 573512
rect 88566 573474 88626 574056
rect 91093 573474 91159 573477
rect 88566 573472 91159 573474
rect 88566 573416 91098 573472
rect 91154 573416 91159 573472
rect 88566 573414 91159 573416
rect 91093 573411 91159 573414
rect 66437 573200 68938 573202
rect 66437 573144 66442 573200
rect 66498 573144 68938 573200
rect 66437 573142 68938 573144
rect 66437 573139 66503 573142
rect 66437 571842 66503 571845
rect 68878 571842 68938 572152
rect 88566 572114 88626 572696
rect 91185 572114 91251 572117
rect 88566 572112 91251 572114
rect 88566 572056 91190 572112
rect 91246 572056 91251 572112
rect 88566 572054 91251 572056
rect 91185 572051 91251 572054
rect 66437 571840 68938 571842
rect 66437 571784 66442 571840
rect 66498 571784 68938 571840
rect 66437 571782 68938 571784
rect 66437 571779 66503 571782
rect 91093 571434 91159 571437
rect 88566 571432 91159 571434
rect 88566 571376 91098 571432
rect 91154 571376 91159 571432
rect 88566 571374 91159 571376
rect 88566 571336 88626 571374
rect 91093 571371 91159 571374
rect 67265 570210 67331 570213
rect 68878 570210 68938 570792
rect 67265 570208 68938 570210
rect 67265 570152 67270 570208
rect 67326 570152 68938 570208
rect 67265 570150 68938 570152
rect 67265 570147 67331 570150
rect 91093 570074 91159 570077
rect 88566 570072 91159 570074
rect 88566 570016 91098 570072
rect 91154 570016 91159 570072
rect 88566 570014 91159 570016
rect 88566 569976 88626 570014
rect 91093 570011 91159 570014
rect 66805 568850 66871 568853
rect 68878 568850 68938 569432
rect 66805 568848 68938 568850
rect 66805 568792 66810 568848
rect 66866 568792 68938 568848
rect 66805 568790 68938 568792
rect 66805 568787 66871 568790
rect 91737 568714 91803 568717
rect 88566 568712 91803 568714
rect 88566 568656 91742 568712
rect 91798 568656 91803 568712
rect 88566 568654 91803 568656
rect 88566 568616 88626 568654
rect 91737 568651 91803 568654
rect 66897 567490 66963 567493
rect 68878 567490 68938 568072
rect 91093 567762 91159 567765
rect 66897 567488 68938 567490
rect 66897 567432 66902 567488
rect 66958 567432 68938 567488
rect 66897 567430 68938 567432
rect 88566 567760 91159 567762
rect 88566 567704 91098 567760
rect 91154 567704 91159 567760
rect 88566 567702 91159 567704
rect 66897 567427 66963 567430
rect 88566 567256 88626 567702
rect 91093 567699 91159 567702
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 67541 566810 67607 566813
rect 67541 566808 68938 566810
rect 67541 566752 67546 566808
rect 67602 566752 68938 566808
rect 67541 566750 68938 566752
rect 67541 566747 67607 566750
rect 68878 566712 68938 566750
rect 88566 565858 88626 565896
rect 91093 565858 91159 565861
rect 88566 565856 91159 565858
rect 88566 565800 91098 565856
rect 91154 565800 91159 565856
rect 88566 565798 91159 565800
rect 91093 565795 91159 565798
rect 66621 564634 66687 564637
rect 68878 564634 68938 565080
rect 66621 564632 68938 564634
rect 66621 564576 66626 564632
rect 66682 564576 68938 564632
rect 66621 564574 68938 564576
rect 66621 564571 66687 564574
rect 88566 564498 88626 564536
rect 91093 564498 91159 564501
rect 88566 564496 91159 564498
rect 88566 564440 91098 564496
rect 91154 564440 91159 564496
rect 88566 564438 91159 564440
rect 91093 564435 91159 564438
rect 582741 564362 582807 564365
rect 583520 564362 584960 564452
rect 582741 564360 584960 564362
rect 582741 564304 582746 564360
rect 582802 564304 584960 564360
rect 582741 564302 584960 564304
rect 582741 564299 582807 564302
rect 583520 564212 584960 564302
rect 66437 564090 66503 564093
rect 66437 564088 68938 564090
rect 66437 564032 66442 564088
rect 66498 564032 68938 564088
rect 66437 564030 68938 564032
rect 66437 564027 66503 564030
rect 68878 563720 68938 564030
rect 88566 563138 88626 563176
rect 91093 563138 91159 563141
rect 88566 563136 91159 563138
rect 88566 563080 91098 563136
rect 91154 563080 91159 563136
rect 88566 563078 91159 563080
rect 91093 563075 91159 563078
rect 66437 562050 66503 562053
rect 68878 562050 68938 562360
rect 66437 562048 68938 562050
rect 66437 561992 66442 562048
rect 66498 561992 68938 562048
rect 66437 561990 68938 561992
rect 66437 561987 66503 561990
rect 66621 560418 66687 560421
rect 68878 560418 68938 561000
rect 88566 560962 88626 561544
rect 91093 560962 91159 560965
rect 88566 560960 91159 560962
rect 88566 560904 91098 560960
rect 91154 560904 91159 560960
rect 88566 560902 91159 560904
rect 91093 560899 91159 560902
rect 66621 560416 68938 560418
rect 66621 560360 66626 560416
rect 66682 560360 68938 560416
rect 66621 560358 68938 560360
rect 66621 560355 66687 560358
rect 88566 560146 88626 560184
rect 89805 560146 89871 560149
rect 91829 560146 91895 560149
rect 88566 560144 91895 560146
rect 88566 560088 89810 560144
rect 89866 560088 91834 560144
rect 91890 560088 91895 560144
rect 88566 560086 91895 560088
rect 89805 560083 89871 560086
rect 91829 560083 91895 560086
rect 66621 559058 66687 559061
rect 68878 559058 68938 559640
rect 66621 559056 68938 559058
rect 66621 559000 66626 559056
rect 66682 559000 68938 559056
rect 66621 558998 68938 559000
rect 66621 558995 66687 558998
rect 67633 558922 67699 558925
rect 67633 558920 68938 558922
rect 67633 558864 67638 558920
rect 67694 558864 68938 558920
rect 67633 558862 68938 558864
rect 67633 558859 67699 558862
rect 68878 558280 68938 558862
rect 88566 558242 88626 558824
rect 91185 558242 91251 558245
rect 88566 558240 91251 558242
rect 88566 558184 91190 558240
rect 91246 558184 91251 558240
rect 88566 558182 91251 558184
rect 91185 558179 91251 558182
rect 67357 556338 67423 556341
rect 68878 556338 68938 556920
rect 88566 556882 88626 557464
rect 91185 556882 91251 556885
rect 88566 556880 91251 556882
rect 88566 556824 91190 556880
rect 91246 556824 91251 556880
rect 88566 556822 91251 556824
rect 91185 556819 91251 556822
rect 67357 556336 68938 556338
rect 67357 556280 67362 556336
rect 67418 556280 68938 556336
rect 67357 556278 68938 556280
rect 67357 556275 67423 556278
rect 66345 555250 66411 555253
rect 68878 555250 68938 555560
rect 88566 555522 88626 556104
rect 91185 555522 91251 555525
rect 88566 555520 91251 555522
rect 88566 555464 91190 555520
rect 91246 555464 91251 555520
rect 88566 555462 91251 555464
rect 91185 555459 91251 555462
rect 66345 555248 68938 555250
rect 66345 555192 66350 555248
rect 66406 555192 68938 555248
rect 66345 555190 68938 555192
rect 66345 555187 66411 555190
rect 66253 554706 66319 554709
rect 66253 554704 68938 554706
rect 66253 554648 66258 554704
rect 66314 554648 68938 554704
rect 66253 554646 68938 554648
rect 66253 554643 66319 554646
rect 68878 554200 68938 554646
rect 88566 554026 88626 554744
rect -960 553890 480 553980
rect 88566 553966 93870 554026
rect 2773 553890 2839 553893
rect -960 553888 2839 553890
rect -960 553832 2778 553888
rect 2834 553832 2839 553888
rect -960 553830 2839 553832
rect -960 553740 480 553830
rect 2773 553827 2839 553830
rect 93810 553482 93870 553966
rect 111006 553482 111012 553484
rect 93810 553422 111012 553482
rect 111006 553420 111012 553422
rect 111076 553420 111082 553484
rect 67449 552258 67515 552261
rect 68878 552258 68938 552840
rect 88566 552802 88626 553384
rect 91277 552802 91343 552805
rect 88566 552800 91343 552802
rect 88566 552744 91282 552800
rect 91338 552744 91343 552800
rect 88566 552742 91343 552744
rect 91277 552739 91343 552742
rect 67449 552256 68938 552258
rect 67449 552200 67454 552256
rect 67510 552200 68938 552256
rect 67449 552198 68938 552200
rect 67449 552195 67515 552198
rect 91185 552122 91251 552125
rect 88566 552120 91251 552122
rect 88566 552064 91190 552120
rect 91246 552064 91251 552120
rect 88566 552062 91251 552064
rect 88566 552024 88626 552062
rect 91185 552059 91251 552062
rect 66662 550836 66668 550900
rect 66732 550898 66738 550900
rect 68878 550898 68938 551480
rect 583520 551020 584960 551260
rect 66732 550838 68938 550898
rect 66732 550836 66738 550838
rect 99966 550762 99972 550764
rect 88566 550702 99972 550762
rect 88566 550664 88626 550702
rect 99966 550700 99972 550702
rect 100036 550700 100042 550764
rect 66529 549674 66595 549677
rect 68878 549674 68938 550120
rect 66529 549672 68938 549674
rect 66529 549616 66534 549672
rect 66590 549616 68938 549672
rect 66529 549614 68938 549616
rect 66529 549611 66595 549614
rect 91185 549402 91251 549405
rect 88566 549400 91251 549402
rect 88566 549344 91190 549400
rect 91246 549344 91251 549400
rect 88566 549342 91251 549344
rect 88566 549304 88626 549342
rect 91185 549339 91251 549342
rect 66529 548314 66595 548317
rect 68878 548314 68938 548760
rect 66529 548312 68938 548314
rect 66529 548256 66534 548312
rect 66590 548256 68938 548312
rect 66529 548254 68938 548256
rect 66529 548251 66595 548254
rect 88566 547906 88626 547944
rect 91185 547906 91251 547909
rect 88566 547904 91251 547906
rect 88566 547848 91190 547904
rect 91246 547848 91251 547904
rect 88566 547846 91251 547848
rect 91185 547843 91251 547846
rect 66805 547634 66871 547637
rect 66805 547632 68938 547634
rect 66805 547576 66810 547632
rect 66866 547576 68938 547632
rect 66805 547574 68938 547576
rect 66805 547571 66871 547574
rect 68878 547400 68938 547574
rect 88566 546546 88626 546584
rect 91277 546546 91343 546549
rect 88566 546544 91343 546546
rect 88566 546488 91282 546544
rect 91338 546488 91343 546544
rect 88566 546486 91343 546488
rect 91277 546483 91343 546486
rect 66161 546410 66227 546413
rect 66161 546408 68938 546410
rect 66161 546352 66166 546408
rect 66222 546352 68938 546408
rect 66161 546350 68938 546352
rect 66161 546347 66227 546350
rect 68878 546040 68938 546350
rect 88566 545186 88626 545224
rect 92565 545186 92631 545189
rect 88566 545184 92631 545186
rect 88566 545128 92570 545184
rect 92626 545128 92631 545184
rect 88566 545126 92631 545128
rect 92565 545123 92631 545126
rect 66805 544914 66871 544917
rect 66805 544912 68938 544914
rect 66805 544856 66810 544912
rect 66866 544856 68938 544912
rect 66805 544854 68938 544856
rect 66805 544851 66871 544854
rect 68878 544680 68938 544854
rect 91277 544098 91343 544101
rect 88566 544096 91343 544098
rect 88566 544040 91282 544096
rect 91338 544040 91343 544096
rect 88566 544038 91343 544040
rect 88566 543864 88626 544038
rect 91277 544035 91343 544038
rect 66805 542738 66871 542741
rect 68878 542738 68938 543320
rect 92565 543010 92631 543013
rect 107694 543010 107700 543012
rect 92565 543008 107700 543010
rect 92565 542952 92570 543008
rect 92626 542952 107700 543008
rect 92565 542950 107700 542952
rect 92565 542947 92631 542950
rect 107694 542948 107700 542950
rect 107764 543010 107770 543012
rect 108113 543010 108179 543013
rect 107764 543008 108179 543010
rect 107764 542952 108118 543008
rect 108174 542952 108179 543008
rect 107764 542950 108179 542952
rect 107764 542948 107770 542950
rect 108113 542947 108179 542950
rect 66805 542736 68938 542738
rect 66805 542680 66810 542736
rect 66866 542680 68938 542736
rect 66805 542678 68938 542680
rect 66805 542675 66871 542678
rect 88566 542466 88626 542504
rect 91277 542466 91343 542469
rect 88566 542464 91343 542466
rect 88566 542408 91282 542464
rect 91338 542408 91343 542464
rect 88566 542406 91343 542408
rect 91277 542403 91343 542406
rect 67081 541786 67147 541789
rect 68878 541786 68938 541960
rect 67081 541784 68938 541786
rect 67081 541728 67086 541784
rect 67142 541728 68938 541784
rect 67081 541726 68938 541728
rect 67081 541723 67147 541726
rect 91277 541378 91343 541381
rect 88566 541376 91343 541378
rect 88566 541320 91282 541376
rect 91338 541320 91343 541376
rect 88566 541318 91343 541320
rect 88566 541144 88626 541318
rect 91277 541315 91343 541318
rect -960 540684 480 540924
rect 68645 540834 68711 540837
rect 68645 540832 68938 540834
rect 68645 540776 68650 540832
rect 68706 540776 68938 540832
rect 68645 540774 68938 540776
rect 68645 540771 68711 540774
rect 68878 540600 68938 540774
rect 88566 539746 88626 539784
rect 91277 539746 91343 539749
rect 88566 539744 91343 539746
rect 88566 539688 91282 539744
rect 91338 539688 91343 539744
rect 88566 539686 91343 539688
rect 91277 539683 91343 539686
rect 76046 539548 76052 539612
rect 76116 539610 76122 539612
rect 76741 539610 76807 539613
rect 76116 539608 76807 539610
rect 76116 539552 76746 539608
rect 76802 539552 76807 539608
rect 76116 539550 76807 539552
rect 76116 539548 76122 539550
rect 76741 539547 76807 539550
rect 115054 538596 115060 538660
rect 115124 538658 115130 538660
rect 115381 538658 115447 538661
rect 115124 538656 115447 538658
rect 115124 538600 115386 538656
rect 115442 538600 115447 538656
rect 115124 538598 115447 538600
rect 115124 538596 115130 538598
rect 115381 538595 115447 538598
rect 579797 537842 579863 537845
rect 583520 537842 584960 537932
rect 579797 537840 584960 537842
rect 579797 537784 579802 537840
rect 579858 537784 584960 537840
rect 579797 537782 584960 537784
rect 579797 537779 579863 537782
rect 583520 537692 584960 537782
rect 76189 536754 76255 536757
rect 124857 536754 124923 536757
rect 76189 536752 124923 536754
rect 76189 536696 76194 536752
rect 76250 536696 124862 536752
rect 124918 536696 124923 536752
rect 76189 536694 124923 536696
rect 76189 536691 76255 536694
rect 124857 536691 124923 536694
rect 84745 536074 84811 536077
rect 128445 536074 128511 536077
rect 582373 536074 582439 536077
rect 84745 536072 582439 536074
rect 84745 536016 84750 536072
rect 84806 536016 128450 536072
rect 128506 536016 582378 536072
rect 582434 536016 582439 536072
rect 84745 536014 582439 536016
rect 84745 536011 84811 536014
rect 128445 536011 128511 536014
rect 582373 536011 582439 536014
rect 68134 535468 68140 535532
rect 68204 535530 68210 535532
rect 68461 535530 68527 535533
rect 69657 535532 69723 535533
rect 69606 535530 69612 535532
rect 68204 535528 68527 535530
rect 68204 535472 68466 535528
rect 68522 535472 68527 535528
rect 68204 535470 68527 535472
rect 69566 535470 69612 535530
rect 69676 535528 69723 535532
rect 69718 535472 69723 535528
rect 68204 535468 68210 535470
rect 68461 535467 68527 535470
rect 69606 535468 69612 535470
rect 69676 535468 69723 535472
rect 69657 535467 69723 535468
rect 70669 535530 70735 535533
rect 71814 535530 71820 535532
rect 70669 535528 71820 535530
rect 70669 535472 70674 535528
rect 70730 535472 71820 535528
rect 70669 535470 71820 535472
rect 70669 535467 70735 535470
rect 71814 535468 71820 535470
rect 71884 535468 71890 535532
rect 76097 535530 76163 535533
rect 76741 535530 76807 535533
rect 76097 535528 76807 535530
rect 76097 535472 76102 535528
rect 76158 535472 76746 535528
rect 76802 535472 76807 535528
rect 76097 535470 76807 535472
rect 76097 535467 76163 535470
rect 76741 535467 76807 535470
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 582465 524514 582531 524517
rect 583520 524514 584960 524604
rect 582465 524512 584960 524514
rect 582465 524456 582470 524512
rect 582526 524456 584960 524512
rect 582465 524454 584960 524456
rect 582465 524451 582531 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3325 501802 3391 501805
rect -960 501800 3391 501802
rect -960 501744 3330 501800
rect 3386 501744 3391 501800
rect -960 501742 3391 501744
rect -960 501652 480 501742
rect 3325 501739 3391 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 582373 484666 582439 484669
rect 583520 484666 584960 484756
rect 582373 484664 584960 484666
rect 582373 484608 582378 484664
rect 582434 484608 584960 484664
rect 582373 484606 584960 484608
rect 582373 484603 582439 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 4061 475690 4127 475693
rect -960 475688 4127 475690
rect -960 475632 4066 475688
rect 4122 475632 4127 475688
rect -960 475630 4127 475632
rect -960 475540 480 475630
rect 4061 475627 4127 475630
rect 582649 471474 582715 471477
rect 583520 471474 584960 471564
rect 582649 471472 584960 471474
rect 582649 471416 582654 471472
rect 582710 471416 584960 471472
rect 582649 471414 584960 471416
rect 582649 471411 582715 471414
rect 583520 471324 584960 471414
rect 96521 465762 96587 465765
rect 106406 465762 106412 465764
rect 96521 465760 106412 465762
rect 96521 465704 96526 465760
rect 96582 465704 106412 465760
rect 96521 465702 106412 465704
rect 96521 465699 96587 465702
rect 106406 465700 106412 465702
rect 106476 465700 106482 465764
rect 93117 464402 93183 464405
rect 102174 464402 102180 464404
rect 93117 464400 102180 464402
rect 93117 464344 93122 464400
rect 93178 464344 102180 464400
rect 93117 464342 102180 464344
rect 93117 464339 93183 464342
rect 102174 464340 102180 464342
rect 102244 464340 102250 464404
rect 81433 462906 81499 462909
rect 89662 462906 89668 462908
rect 81433 462904 89668 462906
rect 81433 462848 81438 462904
rect 81494 462848 89668 462904
rect 81433 462846 89668 462848
rect 81433 462843 81499 462846
rect 89662 462844 89668 462846
rect 89732 462844 89738 462908
rect 94497 462906 94563 462909
rect 104934 462906 104940 462908
rect 94497 462904 104940 462906
rect 94497 462848 94502 462904
rect 94558 462848 104940 462904
rect 94497 462846 104940 462848
rect 94497 462843 94563 462846
rect 104934 462844 104940 462846
rect 105004 462844 105010 462908
rect 107009 462906 107075 462909
rect 115974 462906 115980 462908
rect 107009 462904 115980 462906
rect 107009 462848 107014 462904
rect 107070 462848 115980 462904
rect 107009 462846 115980 462848
rect 107009 462843 107075 462846
rect 115974 462844 115980 462846
rect 116044 462844 116050 462908
rect -960 462634 480 462724
rect 2773 462634 2839 462637
rect -960 462632 2839 462634
rect -960 462576 2778 462632
rect 2834 462576 2839 462632
rect -960 462574 2839 462576
rect -960 462484 480 462574
rect 2773 462571 2839 462574
rect 104157 462226 104223 462229
rect 109166 462226 109172 462228
rect 104157 462224 109172 462226
rect 104157 462168 104162 462224
rect 104218 462168 109172 462224
rect 104157 462166 109172 462168
rect 104157 462163 104223 462166
rect 109166 462164 109172 462166
rect 109236 462164 109242 462228
rect 88190 460124 88196 460188
rect 88260 460186 88266 460188
rect 118693 460186 118759 460189
rect 88260 460184 118759 460186
rect 88260 460128 118698 460184
rect 118754 460128 118759 460184
rect 88260 460126 118759 460128
rect 88260 460124 88266 460126
rect 118693 460123 118759 460126
rect 86953 458826 87019 458829
rect 98126 458826 98132 458828
rect 86953 458824 98132 458826
rect 86953 458768 86958 458824
rect 87014 458768 98132 458824
rect 86953 458766 98132 458768
rect 86953 458763 87019 458766
rect 98126 458764 98132 458766
rect 98196 458764 98202 458828
rect 69657 458282 69723 458285
rect 169017 458282 169083 458285
rect 69657 458280 169083 458282
rect 69657 458224 69662 458280
rect 69718 458224 169022 458280
rect 169078 458224 169083 458280
rect 69657 458222 169083 458224
rect 69657 458219 69723 458222
rect 169017 458219 169083 458222
rect 582465 458146 582531 458149
rect 583520 458146 584960 458236
rect 582465 458144 584960 458146
rect 582465 458088 582470 458144
rect 582526 458088 584960 458144
rect 582465 458086 584960 458088
rect 582465 458083 582531 458086
rect 583520 457996 584960 458086
rect 86861 457466 86927 457469
rect 96654 457466 96660 457468
rect 86861 457464 96660 457466
rect 86861 457408 86866 457464
rect 86922 457408 96660 457464
rect 86861 457406 96660 457408
rect 86861 457403 86927 457406
rect 96654 457404 96660 457406
rect 96724 457404 96730 457468
rect 88333 456106 88399 456109
rect 100702 456106 100708 456108
rect 88333 456104 100708 456106
rect 88333 456048 88338 456104
rect 88394 456048 100708 456104
rect 88333 456046 100708 456048
rect 88333 456043 88399 456046
rect 100702 456044 100708 456046
rect 100772 456044 100778 456108
rect 84101 454746 84167 454749
rect 92606 454746 92612 454748
rect 84101 454744 92612 454746
rect 84101 454688 84106 454744
rect 84162 454688 92612 454744
rect 84101 454686 92612 454688
rect 84101 454683 84167 454686
rect 92606 454684 92612 454686
rect 92676 454684 92682 454748
rect 67766 453868 67772 453932
rect 67836 453930 67842 453932
rect 68318 453930 68324 453932
rect 67836 453870 68324 453930
rect 67836 453868 67842 453870
rect 68318 453868 68324 453870
rect 68388 453868 68394 453932
rect 82721 453250 82787 453253
rect 91318 453250 91324 453252
rect 82721 453248 91324 453250
rect 82721 453192 82726 453248
rect 82782 453192 91324 453248
rect 82721 453190 91324 453192
rect 82721 453187 82787 453190
rect 91318 453188 91324 453190
rect 91388 453188 91394 453252
rect 91737 453250 91803 453253
rect 121637 453250 121703 453253
rect 91737 453248 121703 453250
rect 91737 453192 91742 453248
rect 91798 453192 121642 453248
rect 121698 453192 121703 453248
rect 91737 453190 121703 453192
rect 91737 453187 91803 453190
rect 121637 453187 121703 453190
rect 68318 452644 68324 452708
rect 68388 452706 68394 452708
rect 82077 452706 82143 452709
rect 68388 452704 82143 452706
rect 68388 452648 82082 452704
rect 82138 452648 82143 452704
rect 68388 452646 82143 452648
rect 68388 452644 68394 452646
rect 82077 452643 82143 452646
rect 83457 451346 83523 451349
rect 158662 451346 158668 451348
rect 83457 451344 158668 451346
rect 83457 451288 83462 451344
rect 83518 451288 158668 451344
rect 83457 451286 158668 451288
rect 83457 451283 83523 451286
rect 158662 451284 158668 451286
rect 158732 451284 158738 451348
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 108297 448762 108363 448765
rect 108297 448760 113190 448762
rect 108297 448704 108302 448760
rect 108358 448704 113190 448760
rect 108297 448702 113190 448704
rect 108297 448699 108363 448702
rect 111057 448626 111123 448629
rect 111742 448626 111748 448628
rect 111057 448624 111748 448626
rect 111057 448568 111062 448624
rect 111118 448568 111748 448624
rect 111057 448566 111748 448568
rect 111057 448563 111123 448566
rect 111742 448564 111748 448566
rect 111812 448564 111818 448628
rect 113130 448626 113190 448702
rect 130377 448626 130443 448629
rect 113130 448624 130443 448626
rect 113130 448568 130382 448624
rect 130438 448568 130443 448624
rect 113130 448566 130443 448568
rect 130377 448563 130443 448566
rect 108941 447946 109007 447949
rect 120022 447946 120028 447948
rect 108941 447944 120028 447946
rect 108941 447888 108946 447944
rect 109002 447888 120028 447944
rect 108941 447886 120028 447888
rect 108941 447883 109007 447886
rect 120022 447884 120028 447886
rect 120092 447884 120098 447948
rect 86217 447810 86283 447813
rect 95182 447810 95188 447812
rect 86217 447808 95188 447810
rect 86217 447752 86222 447808
rect 86278 447752 95188 447808
rect 86217 447750 95188 447752
rect 86217 447747 86283 447750
rect 95182 447748 95188 447750
rect 95252 447748 95258 447812
rect 104801 447810 104867 447813
rect 122598 447810 122604 447812
rect 104801 447808 122604 447810
rect 104801 447752 104806 447808
rect 104862 447752 122604 447808
rect 104801 447750 122604 447752
rect 104801 447747 104867 447750
rect 122598 447748 122604 447750
rect 122668 447748 122674 447812
rect 76557 446042 76623 446045
rect 155166 446042 155172 446044
rect 76557 446040 155172 446042
rect 76557 445984 76562 446040
rect 76618 445984 155172 446040
rect 76557 445982 155172 445984
rect 76557 445979 76623 445982
rect 155166 445980 155172 445982
rect 155236 445980 155242 446044
rect 59169 445906 59235 445909
rect 85573 445906 85639 445909
rect 59169 445904 85639 445906
rect 59169 445848 59174 445904
rect 59230 445848 85578 445904
rect 85634 445848 85639 445904
rect 59169 445846 85639 445848
rect 59169 445843 59235 445846
rect 85573 445843 85639 445846
rect 88885 445770 88951 445773
rect 91134 445770 91140 445772
rect 88885 445768 91140 445770
rect 88885 445712 88890 445768
rect 88946 445712 91140 445768
rect 88885 445710 91140 445712
rect 88885 445707 88951 445710
rect 91134 445708 91140 445710
rect 91204 445708 91210 445772
rect 93894 445708 93900 445772
rect 93964 445770 93970 445772
rect 94405 445770 94471 445773
rect 93964 445768 94471 445770
rect 93964 445712 94410 445768
rect 94466 445712 94471 445768
rect 93964 445710 94471 445712
rect 93964 445708 93970 445710
rect 94405 445707 94471 445710
rect 96470 445708 96476 445772
rect 96540 445770 96546 445772
rect 96613 445770 96679 445773
rect 97349 445770 97415 445773
rect 96540 445768 97415 445770
rect 96540 445712 96618 445768
rect 96674 445712 97354 445768
rect 97410 445712 97415 445768
rect 96540 445710 97415 445712
rect 96540 445708 96546 445710
rect 96613 445707 96679 445710
rect 97349 445707 97415 445710
rect 97758 445708 97764 445772
rect 97828 445770 97834 445772
rect 97993 445770 98059 445773
rect 97828 445768 98059 445770
rect 97828 445712 97998 445768
rect 98054 445712 98059 445768
rect 97828 445710 98059 445712
rect 97828 445708 97834 445710
rect 97993 445707 98059 445710
rect 110413 445770 110479 445773
rect 111149 445770 111215 445773
rect 111558 445770 111564 445772
rect 110413 445768 111564 445770
rect 110413 445712 110418 445768
rect 110474 445712 111154 445768
rect 111210 445712 111564 445768
rect 110413 445710 111564 445712
rect 110413 445707 110479 445710
rect 111149 445707 111215 445710
rect 111558 445708 111564 445710
rect 111628 445708 111634 445772
rect 113173 445770 113239 445773
rect 114093 445770 114159 445773
rect 114318 445770 114324 445772
rect 113173 445768 114324 445770
rect 113173 445712 113178 445768
rect 113234 445712 114098 445768
rect 114154 445712 114324 445768
rect 113173 445710 114324 445712
rect 113173 445707 113239 445710
rect 114093 445707 114159 445710
rect 114318 445708 114324 445710
rect 114388 445708 114394 445772
rect 117313 445770 117379 445773
rect 118550 445770 118556 445772
rect 117313 445768 118556 445770
rect 117313 445712 117318 445768
rect 117374 445712 118556 445768
rect 117313 445710 118556 445712
rect 117313 445707 117379 445710
rect 118550 445708 118556 445710
rect 118620 445708 118626 445772
rect 109493 444820 109559 444821
rect 109493 444816 109540 444820
rect 109604 444818 109610 444820
rect 109493 444760 109498 444816
rect 109493 444756 109540 444760
rect 109604 444758 109650 444818
rect 109604 444756 109610 444758
rect 109493 444755 109559 444756
rect 55029 444682 55095 444685
rect 92473 444682 92539 444685
rect 93071 444682 93137 444685
rect 55029 444680 93137 444682
rect 55029 444624 55034 444680
rect 55090 444624 92478 444680
rect 92534 444624 93076 444680
rect 93132 444624 93137 444680
rect 55029 444622 93137 444624
rect 55029 444619 55095 444622
rect 92473 444619 92539 444622
rect 93071 444619 93137 444622
rect 100937 444682 101003 444685
rect 126237 444682 126303 444685
rect 100937 444680 126303 444682
rect 100937 444624 100942 444680
rect 100998 444624 126242 444680
rect 126298 444624 126303 444680
rect 583520 444668 584960 444908
rect 100937 444622 126303 444624
rect 100937 444619 101003 444622
rect 126237 444619 126303 444622
rect 90127 444546 90193 444549
rect 137277 444546 137343 444549
rect 90127 444544 137343 444546
rect 90127 444488 90132 444544
rect 90188 444488 137282 444544
rect 137338 444488 137343 444544
rect 90127 444486 137343 444488
rect 90127 444483 90193 444486
rect 137277 444483 137343 444486
rect 124121 444274 124187 444277
rect 120612 444272 124187 444274
rect 120612 444216 124126 444272
rect 124182 444216 124187 444272
rect 120612 444214 124187 444216
rect 124121 444211 124187 444214
rect 120901 442778 120967 442781
rect 120901 442776 122850 442778
rect 120901 442720 120906 442776
rect 120962 442720 122850 442776
rect 120901 442718 122850 442720
rect 120901 442715 120967 442718
rect 122790 442370 122850 442718
rect 133086 442370 133092 442372
rect 122790 442310 133092 442370
rect 133086 442308 133092 442310
rect 133156 442308 133162 442372
rect 67725 442098 67791 442101
rect 124121 442098 124187 442101
rect 67725 442096 68908 442098
rect 67725 442040 67730 442096
rect 67786 442040 68908 442096
rect 67725 442038 68908 442040
rect 120612 442096 124187 442098
rect 120612 442040 124126 442096
rect 124182 442040 124187 442096
rect 120612 442038 124187 442040
rect 67725 442035 67791 442038
rect 124121 442035 124187 442038
rect 52269 440874 52335 440877
rect 68318 440874 68324 440876
rect 52269 440872 68324 440874
rect 52269 440816 52274 440872
rect 52330 440816 68324 440872
rect 52269 440814 68324 440816
rect 52269 440811 52335 440814
rect 68318 440812 68324 440814
rect 68388 440812 68394 440876
rect 120717 440194 120783 440197
rect 120582 440192 120783 440194
rect 120582 440136 120722 440192
rect 120778 440136 120783 440192
rect 120582 440134 120783 440136
rect 66989 439922 67055 439925
rect 120582 439922 120642 440134
rect 120717 440131 120783 440134
rect 121177 439922 121243 439925
rect 66989 439920 68908 439922
rect 66989 439864 66994 439920
rect 67050 439864 68908 439920
rect 120582 439920 121243 439922
rect 120582 439892 121182 439920
rect 66989 439862 68908 439864
rect 120612 439864 121182 439892
rect 121238 439864 121243 439920
rect 120612 439862 121243 439864
rect 66989 439859 67055 439862
rect 121177 439859 121243 439862
rect 66805 437746 66871 437749
rect 123845 437746 123911 437749
rect 66805 437744 68908 437746
rect 66805 437688 66810 437744
rect 66866 437688 68908 437744
rect 66805 437686 68908 437688
rect 120612 437744 123911 437746
rect 120612 437688 123850 437744
rect 123906 437688 123911 437744
rect 120612 437686 123911 437688
rect 66805 437683 66871 437686
rect 123845 437683 123911 437686
rect -960 436508 480 436748
rect 66805 435298 66871 435301
rect 122966 435298 122972 435300
rect 66805 435296 68908 435298
rect 66805 435240 66810 435296
rect 66866 435240 68908 435296
rect 120612 435268 122972 435298
rect 66805 435238 68908 435240
rect 120582 435238 122972 435268
rect 66805 435235 66871 435238
rect 120582 434754 120642 435238
rect 122966 435236 122972 435238
rect 123036 435236 123042 435300
rect 124857 435298 124923 435301
rect 146886 435298 146892 435300
rect 124857 435296 146892 435298
rect 124857 435240 124862 435296
rect 124918 435240 146892 435296
rect 124857 435238 146892 435240
rect 124857 435235 124923 435238
rect 146886 435236 146892 435238
rect 146956 435236 146962 435300
rect 120717 434754 120783 434757
rect 120582 434752 120783 434754
rect 120582 434696 120722 434752
rect 120778 434696 120783 434752
rect 120582 434694 120783 434696
rect 120717 434691 120783 434694
rect 66897 433122 66963 433125
rect 123109 433122 123175 433125
rect 124121 433122 124187 433125
rect 66897 433120 68908 433122
rect 66897 433064 66902 433120
rect 66958 433064 68908 433120
rect 66897 433062 68908 433064
rect 120612 433120 124187 433122
rect 120612 433064 123114 433120
rect 123170 433064 124126 433120
rect 124182 433064 124187 433120
rect 120612 433062 124187 433064
rect 66897 433059 66963 433062
rect 123109 433059 123175 433062
rect 124121 433059 124187 433062
rect 582373 431626 582439 431629
rect 583520 431626 584960 431716
rect 582373 431624 584960 431626
rect 582373 431568 582378 431624
rect 582434 431568 584960 431624
rect 582373 431566 584960 431568
rect 582373 431563 582439 431566
rect 120022 431428 120028 431492
rect 120092 431428 120098 431492
rect 583520 431476 584960 431566
rect 66897 430946 66963 430949
rect 120030 430946 120090 431428
rect 122598 430946 122604 430948
rect 66897 430944 68908 430946
rect 66897 430888 66902 430944
rect 66958 430888 68908 430944
rect 120030 430916 122604 430946
rect 66897 430886 68908 430888
rect 120060 430886 122604 430916
rect 66897 430883 66963 430886
rect 122598 430884 122604 430886
rect 122668 430884 122674 430948
rect 66805 428498 66871 428501
rect 121545 428498 121611 428501
rect 123293 428498 123359 428501
rect 66805 428496 68908 428498
rect 66805 428440 66810 428496
rect 66866 428440 68908 428496
rect 66805 428438 68908 428440
rect 120612 428496 123359 428498
rect 120612 428440 121550 428496
rect 121606 428440 123298 428496
rect 123354 428440 123359 428496
rect 120612 428438 123359 428440
rect 66805 428435 66871 428438
rect 121545 428435 121611 428438
rect 123293 428435 123359 428438
rect 43989 427138 44055 427141
rect 61837 427138 61903 427141
rect 43989 427136 61903 427138
rect 43989 427080 43994 427136
rect 44050 427080 61842 427136
rect 61898 427080 61903 427136
rect 43989 427078 61903 427080
rect 43989 427075 44055 427078
rect 61837 427075 61903 427078
rect 66253 426322 66319 426325
rect 122414 426322 122420 426324
rect 66253 426320 68908 426322
rect 66253 426264 66258 426320
rect 66314 426264 68908 426320
rect 66253 426262 68908 426264
rect 120612 426262 122420 426322
rect 66253 426259 66319 426262
rect 122414 426260 122420 426262
rect 122484 426260 122490 426324
rect 66110 424084 66116 424148
rect 66180 424146 66186 424148
rect 66253 424146 66319 424149
rect 122925 424146 122991 424149
rect 123201 424146 123267 424149
rect 66180 424144 68908 424146
rect 66180 424088 66258 424144
rect 66314 424088 68908 424144
rect 66180 424086 68908 424088
rect 120612 424144 123267 424146
rect 120612 424088 122930 424144
rect 122986 424088 123206 424144
rect 123262 424088 123267 424144
rect 120612 424086 123267 424088
rect 66180 424084 66186 424086
rect 66253 424083 66319 424086
rect 122925 424083 122991 424086
rect 123201 424083 123267 424086
rect -960 423602 480 423692
rect 3141 423602 3207 423605
rect -960 423600 3207 423602
rect -960 423544 3146 423600
rect 3202 423544 3207 423600
rect -960 423542 3207 423544
rect -960 423452 480 423542
rect 3141 423539 3207 423542
rect 122414 422316 122420 422380
rect 122484 422378 122490 422380
rect 122782 422378 122788 422380
rect 122484 422318 122788 422378
rect 122484 422316 122490 422318
rect 122782 422316 122788 422318
rect 122852 422316 122858 422380
rect 122741 422242 122807 422245
rect 122696 422240 122850 422242
rect 122696 422184 122746 422240
rect 122802 422184 122850 422240
rect 122696 422182 122850 422184
rect 122741 422179 122850 422182
rect 122790 422108 122850 422179
rect 122782 422044 122788 422108
rect 122852 422044 122858 422108
rect 66253 421970 66319 421973
rect 123385 421970 123451 421973
rect 66253 421968 68908 421970
rect 66253 421912 66258 421968
rect 66314 421912 68908 421968
rect 66253 421910 68908 421912
rect 120612 421968 123451 421970
rect 120612 421912 123390 421968
rect 123446 421912 123451 421968
rect 120612 421910 123451 421912
rect 66253 421907 66319 421910
rect 123385 421907 123451 421910
rect 67357 419522 67423 419525
rect 120809 419522 120875 419525
rect 67357 419520 69276 419522
rect 67357 419464 67362 419520
rect 67418 419492 69276 419520
rect 120612 419520 120875 419522
rect 67418 419464 69306 419492
rect 67357 419462 69306 419464
rect 120612 419464 120814 419520
rect 120870 419464 120875 419520
rect 120612 419462 120875 419464
rect 67357 419459 67423 419462
rect 69246 419388 69306 419462
rect 120809 419459 120875 419462
rect 69238 419324 69244 419388
rect 69308 419324 69314 419388
rect 582465 418298 582531 418301
rect 583520 418298 584960 418388
rect 582465 418296 584960 418298
rect 582465 418240 582470 418296
rect 582526 418240 584960 418296
rect 582465 418238 584960 418240
rect 582465 418235 582531 418238
rect 583520 418148 584960 418238
rect 66897 417346 66963 417349
rect 121545 417346 121611 417349
rect 66897 417344 68908 417346
rect 66897 417288 66902 417344
rect 66958 417288 68908 417344
rect 66897 417286 68908 417288
rect 120612 417344 121611 417346
rect 120612 417288 121550 417344
rect 121606 417288 121611 417344
rect 120612 417286 121611 417288
rect 66897 417283 66963 417286
rect 121545 417283 121611 417286
rect 66437 415170 66503 415173
rect 123109 415170 123175 415173
rect 66437 415168 68908 415170
rect 66437 415112 66442 415168
rect 66498 415112 68908 415168
rect 66437 415110 68908 415112
rect 120612 415168 123175 415170
rect 120612 415112 123114 415168
rect 123170 415112 123175 415168
rect 120612 415110 123175 415112
rect 66437 415107 66503 415110
rect 123109 415107 123175 415110
rect 122741 412860 122807 412861
rect 122741 412858 122788 412860
rect 122696 412856 122788 412858
rect 122852 412858 122858 412860
rect 122696 412800 122746 412856
rect 122696 412798 122788 412800
rect 122741 412796 122788 412798
rect 122852 412798 122934 412858
rect 122852 412796 122858 412798
rect 122741 412795 122807 412796
rect 67449 412722 67515 412725
rect 123109 412722 123175 412725
rect 67449 412720 68908 412722
rect 67449 412664 67454 412720
rect 67510 412664 68908 412720
rect 67449 412662 68908 412664
rect 120612 412720 123175 412722
rect 120612 412664 123114 412720
rect 123170 412664 123175 412720
rect 120612 412662 123175 412664
rect 67449 412659 67515 412662
rect 123109 412659 123175 412662
rect 122741 412586 122807 412589
rect 122696 412584 122850 412586
rect 122696 412528 122746 412584
rect 122802 412528 122850 412584
rect 122696 412526 122850 412528
rect 122741 412523 122850 412526
rect 122790 412452 122850 412523
rect 122782 412388 122788 412452
rect 122852 412388 122858 412452
rect 54937 411362 55003 411365
rect 66662 411362 66668 411364
rect 54937 411360 66668 411362
rect 54937 411304 54942 411360
rect 54998 411304 66668 411360
rect 54937 411302 66668 411304
rect 54937 411299 55003 411302
rect 66662 411300 66668 411302
rect 66732 411362 66738 411364
rect 66732 411302 66914 411362
rect 66732 411300 66738 411302
rect 66854 411226 66914 411302
rect 66854 411166 68938 411226
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect 68878 410516 68938 411166
rect 121637 410546 121703 410549
rect 120612 410544 121703 410546
rect -960 410486 3483 410488
rect 120612 410488 121642 410544
rect 121698 410488 121703 410544
rect 120612 410486 121703 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 121637 410483 121703 410486
rect 66529 408370 66595 408373
rect 124121 408370 124187 408373
rect 66529 408368 68908 408370
rect 66529 408312 66534 408368
rect 66590 408312 68908 408368
rect 66529 408310 68908 408312
rect 120612 408368 124187 408370
rect 120612 408312 124126 408368
rect 124182 408312 124187 408368
rect 120612 408310 124187 408312
rect 66529 408307 66595 408310
rect 124121 408307 124187 408310
rect 66621 406194 66687 406197
rect 123569 406194 123635 406197
rect 66621 406192 68908 406194
rect 66621 406136 66626 406192
rect 66682 406136 68908 406192
rect 66621 406134 68908 406136
rect 120612 406192 123635 406194
rect 120612 406136 123574 406192
rect 123630 406136 123635 406192
rect 120612 406134 123635 406136
rect 66621 406131 66687 406134
rect 123569 406131 123635 406134
rect 582557 404970 582623 404973
rect 583520 404970 584960 405060
rect 582557 404968 584960 404970
rect 582557 404912 582562 404968
rect 582618 404912 584960 404968
rect 582557 404910 584960 404912
rect 582557 404907 582623 404910
rect 583520 404820 584960 404910
rect 120625 404290 120691 404293
rect 120582 404288 120691 404290
rect 120582 404232 120630 404288
rect 120686 404232 120691 404288
rect 120582 404227 120691 404232
rect 66345 403746 66411 403749
rect 66345 403744 68908 403746
rect 66345 403688 66350 403744
rect 66406 403688 68908 403744
rect 120582 403716 120642 404227
rect 66345 403686 68908 403688
rect 66345 403683 66411 403686
rect 122741 403068 122807 403069
rect 122741 403066 122788 403068
rect 122696 403064 122788 403066
rect 122852 403066 122858 403068
rect 122696 403008 122746 403064
rect 122696 403006 122788 403008
rect 122741 403004 122788 403006
rect 122852 403006 122934 403066
rect 122852 403004 122858 403006
rect 122741 403003 122807 403004
rect 122741 402930 122807 402933
rect 122966 402930 122972 402932
rect 122696 402928 122972 402930
rect 122696 402872 122746 402928
rect 122802 402872 122972 402928
rect 122696 402870 122972 402872
rect 122741 402867 122807 402870
rect 122966 402868 122972 402870
rect 123036 402868 123042 402932
rect 66805 401570 66871 401573
rect 124121 401570 124187 401573
rect 66805 401568 68908 401570
rect 66805 401512 66810 401568
rect 66866 401512 68908 401568
rect 66805 401510 68908 401512
rect 120612 401568 124187 401570
rect 120612 401512 124126 401568
rect 124182 401512 124187 401568
rect 120612 401510 124187 401512
rect 66805 401507 66871 401510
rect 124121 401507 124187 401510
rect 66897 399394 66963 399397
rect 123661 399394 123727 399397
rect 66897 399392 68908 399394
rect 66897 399336 66902 399392
rect 66958 399336 68908 399392
rect 66897 399334 68908 399336
rect 120612 399392 123727 399394
rect 120612 399336 123666 399392
rect 123722 399336 123727 399392
rect 120612 399334 123727 399336
rect 66897 399331 66963 399334
rect 123661 399331 123727 399334
rect -960 397490 480 397580
rect 2773 397490 2839 397493
rect -960 397488 2839 397490
rect -960 397432 2778 397488
rect 2834 397432 2839 397488
rect -960 397430 2839 397432
rect -960 397340 480 397430
rect 2773 397427 2839 397430
rect 66253 396946 66319 396949
rect 67357 396946 67423 396949
rect 121453 396946 121519 396949
rect 66253 396944 68908 396946
rect 66253 396888 66258 396944
rect 66314 396888 67362 396944
rect 67418 396888 68908 396944
rect 66253 396886 68908 396888
rect 120612 396944 121519 396946
rect 120612 396888 121458 396944
rect 121514 396888 121519 396944
rect 120612 396886 121519 396888
rect 66253 396883 66319 396886
rect 67357 396883 67423 396886
rect 121453 396883 121519 396886
rect 67541 394770 67607 394773
rect 122966 394770 122972 394772
rect 67541 394768 68908 394770
rect 67541 394712 67546 394768
rect 67602 394712 68908 394768
rect 67541 394710 68908 394712
rect 120612 394710 122972 394770
rect 67541 394707 67607 394710
rect 122966 394708 122972 394710
rect 123036 394770 123042 394772
rect 124121 394770 124187 394773
rect 123036 394768 124187 394770
rect 123036 394712 124126 394768
rect 124182 394712 124187 394768
rect 123036 394710 124187 394712
rect 123036 394708 123042 394710
rect 124121 394707 124187 394710
rect 122741 393412 122807 393413
rect 122741 393410 122788 393412
rect 122696 393408 122788 393410
rect 122852 393410 122858 393412
rect 122696 393352 122746 393408
rect 122696 393350 122788 393352
rect 122741 393348 122788 393350
rect 122852 393350 122934 393410
rect 122852 393348 122858 393350
rect 122741 393347 122807 393348
rect 122741 393276 122807 393277
rect 122741 393274 122788 393276
rect 122696 393272 122788 393274
rect 122852 393274 122858 393276
rect 122696 393216 122746 393272
rect 122696 393214 122788 393216
rect 122741 393212 122788 393214
rect 122852 393214 122934 393274
rect 122852 393212 122858 393214
rect 122741 393211 122807 393212
rect 65517 392594 65583 392597
rect 121453 392594 121519 392597
rect 123017 392594 123083 392597
rect 65517 392592 68908 392594
rect 65517 392536 65522 392592
rect 65578 392536 68908 392592
rect 65517 392534 68908 392536
rect 120612 392592 123083 392594
rect 120612 392536 121458 392592
rect 121514 392536 123022 392592
rect 123078 392536 123083 392592
rect 120612 392534 123083 392536
rect 65517 392531 65583 392534
rect 121453 392531 121519 392534
rect 123017 392531 123083 392534
rect 583520 391628 584960 391868
rect 65977 391098 66043 391101
rect 65977 391096 70410 391098
rect 65977 391040 65982 391096
rect 66038 391040 70410 391096
rect 65977 391038 70410 391040
rect 65977 391035 66043 391038
rect 70350 390962 70410 391038
rect 86217 390962 86283 390965
rect 70350 390960 86283 390962
rect 70350 390904 86222 390960
rect 86278 390904 86283 390960
rect 70350 390902 86283 390904
rect 86217 390899 86283 390902
rect 92606 390900 92612 390964
rect 92676 390962 92682 390964
rect 92749 390962 92815 390965
rect 102133 390964 102199 390965
rect 102133 390962 102180 390964
rect 92676 390960 92815 390962
rect 92676 390904 92754 390960
rect 92810 390904 92815 390960
rect 92676 390902 92815 390904
rect 102088 390960 102180 390962
rect 102088 390904 102138 390960
rect 102088 390902 102180 390904
rect 92676 390900 92682 390902
rect 92749 390899 92815 390902
rect 102133 390900 102180 390902
rect 102244 390900 102250 390964
rect 107929 390962 107995 390965
rect 114093 390962 114159 390965
rect 107929 390960 114159 390962
rect 107929 390904 107934 390960
rect 107990 390904 114098 390960
rect 114154 390904 114159 390960
rect 107929 390902 114159 390904
rect 102133 390899 102199 390900
rect 107929 390899 107995 390902
rect 114093 390899 114159 390902
rect 69606 390628 69612 390692
rect 69676 390690 69682 390692
rect 70025 390690 70091 390693
rect 69676 390688 70091 390690
rect 69676 390632 70030 390688
rect 70086 390632 70091 390688
rect 69676 390630 70091 390632
rect 69676 390628 69682 390630
rect 70025 390627 70091 390630
rect 115749 390690 115815 390693
rect 120809 390690 120875 390693
rect 115749 390688 120875 390690
rect 115749 390632 115754 390688
rect 115810 390632 120814 390688
rect 120870 390632 120875 390688
rect 115749 390630 120875 390632
rect 115749 390627 115815 390630
rect 120809 390627 120875 390630
rect 71865 390420 71931 390421
rect 71814 390418 71820 390420
rect 71774 390358 71820 390418
rect 71884 390416 71931 390420
rect 71926 390360 71931 390416
rect 71814 390356 71820 390358
rect 71884 390356 71931 390360
rect 71865 390355 71931 390356
rect 80053 390418 80119 390421
rect 80605 390418 80671 390421
rect 91369 390420 91435 390421
rect 91318 390418 91324 390420
rect 80053 390416 80671 390418
rect 80053 390360 80058 390416
rect 80114 390360 80610 390416
rect 80666 390360 80671 390416
rect 80053 390358 80671 390360
rect 91278 390358 91324 390418
rect 91388 390416 91435 390420
rect 91430 390360 91435 390416
rect 80053 390355 80119 390358
rect 80605 390355 80671 390358
rect 91318 390356 91324 390358
rect 91388 390356 91435 390360
rect 95182 390356 95188 390420
rect 95252 390418 95258 390420
rect 95877 390418 95943 390421
rect 95252 390416 95943 390418
rect 95252 390360 95882 390416
rect 95938 390360 95943 390416
rect 95252 390358 95943 390360
rect 95252 390356 95258 390358
rect 91369 390355 91435 390356
rect 95877 390355 95943 390358
rect 96654 390356 96660 390420
rect 96724 390418 96730 390420
rect 97349 390418 97415 390421
rect 96724 390416 97415 390418
rect 96724 390360 97354 390416
rect 97410 390360 97415 390416
rect 96724 390358 97415 390360
rect 96724 390356 96730 390358
rect 97349 390355 97415 390358
rect 98126 390356 98132 390420
rect 98196 390418 98202 390420
rect 98821 390418 98887 390421
rect 98196 390416 98887 390418
rect 98196 390360 98826 390416
rect 98882 390360 98887 390416
rect 98196 390358 98887 390360
rect 98196 390356 98202 390358
rect 98821 390355 98887 390358
rect 100661 390420 100727 390421
rect 104985 390420 105051 390421
rect 100661 390416 100708 390420
rect 100772 390418 100778 390420
rect 104934 390418 104940 390420
rect 100661 390360 100666 390416
rect 100661 390356 100708 390360
rect 100772 390358 100818 390418
rect 104894 390358 104940 390418
rect 105004 390416 105051 390420
rect 105046 390360 105051 390416
rect 100772 390356 100778 390358
rect 104934 390356 104940 390358
rect 105004 390356 105051 390360
rect 106406 390356 106412 390420
rect 106476 390418 106482 390420
rect 106549 390418 106615 390421
rect 106476 390416 106615 390418
rect 106476 390360 106554 390416
rect 106610 390360 106615 390416
rect 106476 390358 106615 390360
rect 106476 390356 106482 390358
rect 100661 390355 100727 390356
rect 104985 390355 105051 390356
rect 106549 390355 106615 390358
rect 107694 390356 107700 390420
rect 107764 390418 107770 390420
rect 108021 390418 108087 390421
rect 107764 390416 108087 390418
rect 107764 390360 108026 390416
rect 108082 390360 108087 390416
rect 107764 390358 108087 390360
rect 107764 390356 107770 390358
rect 108021 390355 108087 390358
rect 109166 390356 109172 390420
rect 109236 390418 109242 390420
rect 109493 390418 109559 390421
rect 109236 390416 109559 390418
rect 109236 390360 109498 390416
rect 109554 390360 109559 390416
rect 109236 390358 109559 390360
rect 109236 390356 109242 390358
rect 109493 390355 109559 390358
rect 115933 390420 115999 390421
rect 115933 390416 115980 390420
rect 116044 390418 116050 390420
rect 115933 390360 115938 390416
rect 115933 390356 115980 390360
rect 116044 390358 116090 390418
rect 116044 390356 116050 390358
rect 120022 390356 120028 390420
rect 120092 390418 120098 390420
rect 120165 390418 120231 390421
rect 120092 390416 120231 390418
rect 120092 390360 120170 390416
rect 120226 390360 120231 390416
rect 120092 390358 120231 390360
rect 120092 390356 120098 390358
rect 115933 390355 115999 390356
rect 120165 390355 120231 390358
rect 66161 389194 66227 389197
rect 80053 389194 80119 389197
rect 66161 389192 80119 389194
rect 66161 389136 66166 389192
rect 66222 389136 80058 389192
rect 80114 389136 80119 389192
rect 66161 389134 80119 389136
rect 66161 389131 66227 389134
rect 80053 389131 80119 389134
rect 111006 389132 111012 389196
rect 111076 389194 111082 389196
rect 118693 389194 118759 389197
rect 111076 389192 118759 389194
rect 111076 389136 118698 389192
rect 118754 389136 118759 389192
rect 111076 389134 118759 389136
rect 111076 389132 111082 389134
rect 118693 389131 118759 389134
rect 68645 389058 68711 389061
rect 76414 389058 76420 389060
rect 68645 389056 76420 389058
rect 68645 389000 68650 389056
rect 68706 389000 76420 389056
rect 68645 388998 76420 389000
rect 68645 388995 68711 388998
rect 76414 388996 76420 388998
rect 76484 388996 76490 389060
rect 89662 389058 89668 389060
rect 84150 388998 89668 389058
rect 3417 388922 3483 388925
rect 84150 388922 84210 388998
rect 89662 388996 89668 388998
rect 89732 389058 89738 389060
rect 89805 389058 89871 389061
rect 89732 389056 89871 389058
rect 89732 389000 89810 389056
rect 89866 389000 89871 389056
rect 89732 388998 89871 389000
rect 89732 388996 89738 388998
rect 89805 388995 89871 388998
rect 101121 389058 101187 389061
rect 101949 389058 102015 389061
rect 101121 389056 102015 389058
rect 101121 389000 101126 389056
rect 101182 389000 101954 389056
rect 102010 389000 102015 389056
rect 101121 388998 102015 389000
rect 101121 388995 101187 388998
rect 101949 388995 102015 388998
rect 111742 388996 111748 389060
rect 111812 389058 111818 389060
rect 112621 389058 112687 389061
rect 111812 389056 112687 389058
rect 111812 389000 112626 389056
rect 112682 389000 112687 389056
rect 111812 388998 112687 389000
rect 111812 388996 111818 388998
rect 112621 388995 112687 388998
rect 3417 388920 84210 388922
rect 3417 388864 3422 388920
rect 3478 388864 84210 388920
rect 3417 388862 84210 388864
rect 3417 388859 3483 388862
rect 67766 388724 67772 388788
rect 67836 388786 67842 388788
rect 68134 388786 68140 388788
rect 67836 388726 68140 388786
rect 67836 388724 67842 388726
rect 68134 388724 68140 388726
rect 68204 388786 68210 388788
rect 68829 388786 68895 388789
rect 68204 388784 68895 388786
rect 68204 388728 68834 388784
rect 68890 388728 68895 388784
rect 68204 388726 68895 388728
rect 68204 388724 68210 388726
rect 68829 388723 68895 388726
rect 95233 388514 95299 388517
rect 96470 388514 96476 388516
rect 95233 388512 96476 388514
rect 95233 388456 95238 388512
rect 95294 388456 96476 388512
rect 95233 388454 96476 388456
rect 95233 388451 95299 388454
rect 96470 388452 96476 388454
rect 96540 388452 96546 388516
rect 91001 388378 91067 388381
rect 99966 388378 99972 388380
rect 91001 388376 99972 388378
rect 91001 388320 91006 388376
rect 91062 388320 99972 388376
rect 91001 388318 99972 388320
rect 91001 388315 91067 388318
rect 99966 388316 99972 388318
rect 100036 388378 100042 388380
rect 107929 388378 107995 388381
rect 100036 388376 107995 388378
rect 100036 388320 107934 388376
rect 107990 388320 107995 388376
rect 100036 388318 107995 388320
rect 100036 388316 100042 388318
rect 107929 388315 107995 388318
rect 53465 387698 53531 387701
rect 83549 387698 83615 387701
rect 53465 387696 83615 387698
rect 53465 387640 53470 387696
rect 53526 387640 83554 387696
rect 83610 387640 83615 387696
rect 53465 387638 83615 387640
rect 53465 387635 53531 387638
rect 83549 387635 83615 387638
rect 83406 387228 83412 387292
rect 83476 387290 83482 387292
rect 83549 387290 83615 387293
rect 83476 387288 83615 387290
rect 83476 387232 83554 387288
rect 83610 387232 83615 387288
rect 83476 387230 83615 387232
rect 83476 387228 83482 387230
rect 83549 387227 83615 387230
rect 3417 387018 3483 387021
rect 95877 387018 95943 387021
rect 3417 387016 95943 387018
rect 3417 386960 3422 387016
rect 3478 386960 95882 387016
rect 95938 386960 95943 387016
rect 3417 386958 95943 386960
rect 3417 386955 3483 386958
rect 95877 386955 95943 386958
rect 52361 385658 52427 385661
rect 122966 385658 122972 385660
rect 52361 385656 122972 385658
rect 52361 385600 52366 385656
rect 52422 385600 122972 385656
rect 52361 385598 122972 385600
rect 52361 385595 52427 385598
rect 122966 385596 122972 385598
rect 123036 385596 123042 385660
rect -960 384284 480 384524
rect 122782 383828 122788 383892
rect 122852 383828 122858 383892
rect 122790 383757 122850 383828
rect 122741 383754 122850 383757
rect 122696 383752 122850 383754
rect 122696 383696 122746 383752
rect 122802 383696 122850 383752
rect 122696 383694 122850 383696
rect 122741 383691 122807 383694
rect 122741 383620 122807 383621
rect 122741 383618 122788 383620
rect 122696 383616 122788 383618
rect 122852 383618 122858 383620
rect 122696 383560 122746 383616
rect 122696 383558 122788 383560
rect 122741 383556 122788 383558
rect 122852 383558 122934 383618
rect 122852 383556 122858 383558
rect 122741 383555 122807 383556
rect 115105 382260 115171 382261
rect 115054 382258 115060 382260
rect 115014 382198 115060 382258
rect 115124 382256 115171 382260
rect 115166 382200 115171 382256
rect 115054 382196 115060 382198
rect 115124 382196 115171 382200
rect 115105 382195 115171 382196
rect 7557 381578 7623 381581
rect 104985 381578 105051 381581
rect 105629 381578 105695 381581
rect 7557 381576 105695 381578
rect 7557 381520 7562 381576
rect 7618 381520 104990 381576
rect 105046 381520 105634 381576
rect 105690 381520 105695 381576
rect 7557 381518 105695 381520
rect 7557 381515 7623 381518
rect 104985 381515 105051 381518
rect 105629 381515 105695 381518
rect 85481 378858 85547 378861
rect 89662 378858 89668 378860
rect 85481 378856 89668 378858
rect 85481 378800 85486 378856
rect 85542 378800 89668 378856
rect 85481 378798 89668 378800
rect 85481 378795 85547 378798
rect 89662 378796 89668 378798
rect 89732 378796 89738 378860
rect 88241 378722 88307 378725
rect 136582 378722 136588 378724
rect 88241 378720 136588 378722
rect 88241 378664 88246 378720
rect 88302 378664 136588 378720
rect 88241 378662 136588 378664
rect 88241 378659 88307 378662
rect 136582 378660 136588 378662
rect 136652 378660 136658 378724
rect 582741 378450 582807 378453
rect 583520 378450 584960 378540
rect 582741 378448 584960 378450
rect 582741 378392 582746 378448
rect 582802 378392 584960 378448
rect 582741 378390 584960 378392
rect 582741 378387 582807 378390
rect 583520 378300 584960 378390
rect 58985 377362 59051 377365
rect 163446 377362 163452 377364
rect 58985 377360 163452 377362
rect 58985 377304 58990 377360
rect 59046 377304 163452 377360
rect 58985 377302 163452 377304
rect 58985 377299 59051 377302
rect 163446 377300 163452 377302
rect 163516 377300 163522 377364
rect 122782 374172 122788 374236
rect 122852 374172 122858 374236
rect 122790 374101 122850 374172
rect 122741 374098 122850 374101
rect 122696 374096 122850 374098
rect 122696 374040 122746 374096
rect 122802 374040 122850 374096
rect 122696 374038 122850 374040
rect 122741 374035 122807 374038
rect 122741 373964 122807 373965
rect 122741 373962 122788 373964
rect 122696 373960 122788 373962
rect 122852 373962 122858 373964
rect 122696 373904 122746 373960
rect 122696 373902 122788 373904
rect 122741 373900 122788 373902
rect 122852 373902 122934 373962
rect 122852 373900 122858 373902
rect 122741 373899 122807 373900
rect -960 371378 480 371468
rect 3509 371378 3575 371381
rect -960 371376 3575 371378
rect -960 371320 3514 371376
rect 3570 371320 3575 371376
rect -960 371318 3575 371320
rect -960 371228 480 371318
rect 3509 371315 3575 371318
rect 120717 371378 120783 371381
rect 244222 371378 244228 371380
rect 120717 371376 244228 371378
rect 120717 371320 120722 371376
rect 120778 371320 244228 371376
rect 120717 371318 244228 371320
rect 120717 371315 120783 371318
rect 244222 371316 244228 371318
rect 244292 371316 244298 371380
rect 114318 369956 114324 370020
rect 114388 370018 114394 370020
rect 119337 370018 119403 370021
rect 114388 370016 119403 370018
rect 114388 369960 119342 370016
rect 119398 369960 119403 370016
rect 114388 369958 119403 369960
rect 114388 369956 114394 369958
rect 119337 369955 119403 369958
rect 97257 369882 97323 369885
rect 97758 369882 97764 369884
rect 97257 369880 97764 369882
rect 97257 369824 97262 369880
rect 97318 369824 97764 369880
rect 97257 369822 97764 369824
rect 97257 369819 97323 369822
rect 97758 369820 97764 369822
rect 97828 369882 97834 369884
rect 252502 369882 252508 369884
rect 97828 369822 252508 369882
rect 97828 369820 97834 369822
rect 252502 369820 252508 369822
rect 252572 369820 252578 369884
rect 141417 369066 141483 369069
rect 169702 369066 169708 369068
rect 141417 369064 169708 369066
rect 141417 369008 141422 369064
rect 141478 369008 169708 369064
rect 141417 369006 169708 369008
rect 141417 369003 141483 369006
rect 169702 369004 169708 369006
rect 169772 369004 169778 369068
rect 69790 367644 69796 367708
rect 69860 367706 69866 367708
rect 123477 367706 123543 367709
rect 69860 367704 123543 367706
rect 69860 367648 123482 367704
rect 123538 367648 123543 367704
rect 69860 367646 123543 367648
rect 69860 367644 69866 367646
rect 123477 367643 123543 367646
rect 135069 367298 135135 367301
rect 185577 367298 185643 367301
rect 135069 367296 185643 367298
rect 135069 367240 135074 367296
rect 135130 367240 185582 367296
rect 185638 367240 185643 367296
rect 135069 367238 185643 367240
rect 135069 367235 135135 367238
rect 185577 367235 185643 367238
rect 102041 367162 102107 367165
rect 321553 367162 321619 367165
rect 102041 367160 321619 367162
rect 102041 367104 102046 367160
rect 102102 367104 321558 367160
rect 321614 367104 321619 367160
rect 102041 367102 321619 367104
rect 102041 367099 102107 367102
rect 321553 367099 321619 367102
rect 135897 367026 135963 367029
rect 138013 367026 138079 367029
rect 135897 367024 138079 367026
rect 135897 366968 135902 367024
rect 135958 366968 138018 367024
rect 138074 366968 138079 367024
rect 135897 366966 138079 366968
rect 135897 366963 135963 366966
rect 138013 366963 138079 366966
rect 61929 366346 61995 366349
rect 69054 366346 69060 366348
rect 61929 366344 69060 366346
rect 61929 366288 61934 366344
rect 61990 366288 69060 366344
rect 61929 366286 69060 366288
rect 61929 366283 61995 366286
rect 69054 366284 69060 366286
rect 69124 366346 69130 366348
rect 85573 366346 85639 366349
rect 69124 366344 85639 366346
rect 69124 366288 85578 366344
rect 85634 366288 85639 366344
rect 69124 366286 85639 366288
rect 69124 366284 69130 366286
rect 85573 366283 85639 366286
rect 146886 365876 146892 365940
rect 146956 365938 146962 365940
rect 218237 365938 218303 365941
rect 146956 365936 218303 365938
rect 146956 365880 218242 365936
rect 218298 365880 218303 365936
rect 146956 365878 218303 365880
rect 146956 365876 146962 365878
rect 218237 365875 218303 365878
rect 138013 365802 138079 365805
rect 222326 365802 222332 365804
rect 138013 365800 222332 365802
rect 138013 365744 138018 365800
rect 138074 365744 222332 365800
rect 138013 365742 222332 365744
rect 138013 365739 138079 365742
rect 222326 365740 222332 365742
rect 222396 365740 222402 365804
rect 582373 365122 582439 365125
rect 583520 365122 584960 365212
rect 582373 365120 584960 365122
rect 582373 365064 582378 365120
rect 582434 365064 584960 365120
rect 582373 365062 584960 365064
rect 582373 365059 582439 365062
rect 80053 364986 80119 364989
rect 157333 364986 157399 364989
rect 80053 364984 157399 364986
rect 80053 364928 80058 364984
rect 80114 364928 157338 364984
rect 157394 364928 157399 364984
rect 583520 364972 584960 365062
rect 80053 364926 157399 364928
rect 80053 364923 80119 364926
rect 157333 364923 157399 364926
rect 122741 364578 122807 364581
rect 122966 364578 122972 364580
rect 122696 364576 122972 364578
rect 122696 364520 122746 364576
rect 122802 364520 122972 364576
rect 122696 364518 122972 364520
rect 122741 364515 122807 364518
rect 122966 364516 122972 364518
rect 123036 364516 123042 364580
rect 114553 364442 114619 364445
rect 115841 364442 115907 364445
rect 227437 364442 227503 364445
rect 114553 364440 227503 364442
rect 114553 364384 114558 364440
rect 114614 364384 115846 364440
rect 115902 364384 227442 364440
rect 227498 364384 227503 364440
rect 114553 364382 227503 364384
rect 114553 364379 114619 364382
rect 115841 364379 115907 364382
rect 227437 364379 227503 364382
rect 100109 364306 100175 364309
rect 150249 364306 150315 364309
rect 100109 364304 150315 364306
rect 100109 364248 100114 364304
rect 100170 364248 150254 364304
rect 150310 364248 150315 364304
rect 100109 364246 150315 364248
rect 100109 364243 100175 364246
rect 150249 364243 150315 364246
rect 122741 364170 122807 364173
rect 122966 364170 122972 364172
rect 122696 364168 122972 364170
rect 122696 364112 122746 364168
rect 122802 364112 122972 364168
rect 122696 364110 122972 364112
rect 122741 364107 122807 364110
rect 122966 364108 122972 364110
rect 123036 364108 123042 364172
rect 150249 363218 150315 363221
rect 150433 363218 150499 363221
rect 150249 363216 150499 363218
rect 150249 363160 150254 363216
rect 150310 363160 150438 363216
rect 150494 363160 150499 363216
rect 150249 363158 150499 363160
rect 150249 363155 150315 363158
rect 150433 363155 150499 363158
rect 87597 363082 87663 363085
rect 238017 363082 238083 363085
rect 87597 363080 238083 363082
rect 87597 363024 87602 363080
rect 87658 363024 238022 363080
rect 238078 363024 238083 363080
rect 87597 363022 238083 363024
rect 87597 363019 87663 363022
rect 238017 363019 238083 363022
rect 76557 362266 76623 362269
rect 138054 362266 138060 362268
rect 76557 362264 138060 362266
rect 76557 362208 76562 362264
rect 76618 362208 138060 362264
rect 76557 362206 138060 362208
rect 76557 362203 76623 362206
rect 138054 362204 138060 362206
rect 138124 362204 138130 362268
rect 111057 361858 111123 361861
rect 111558 361858 111564 361860
rect 111057 361856 111564 361858
rect 111057 361800 111062 361856
rect 111118 361800 111564 361856
rect 111057 361798 111564 361800
rect 111057 361795 111123 361798
rect 111558 361796 111564 361798
rect 111628 361858 111634 361860
rect 204253 361858 204319 361861
rect 111628 361856 204319 361858
rect 111628 361800 204258 361856
rect 204314 361800 204319 361856
rect 111628 361798 204319 361800
rect 111628 361796 111634 361798
rect 204253 361795 204319 361798
rect 121453 361722 121519 361725
rect 122598 361722 122604 361724
rect 121453 361720 122604 361722
rect 121453 361664 121458 361720
rect 121514 361664 122604 361720
rect 121453 361662 122604 361664
rect 121453 361659 121519 361662
rect 122598 361660 122604 361662
rect 122668 361722 122674 361724
rect 232497 361722 232563 361725
rect 122668 361720 232563 361722
rect 122668 361664 232502 361720
rect 232558 361664 232563 361720
rect 122668 361662 232563 361664
rect 122668 361660 122674 361662
rect 232497 361659 232563 361662
rect 96521 361042 96587 361045
rect 96521 361040 126898 361042
rect 96521 360984 96526 361040
rect 96582 360984 126898 361040
rect 96521 360982 126898 360984
rect 96521 360979 96587 360982
rect 70158 360844 70164 360908
rect 70228 360906 70234 360908
rect 123293 360906 123359 360909
rect 70228 360904 123359 360906
rect 70228 360848 123298 360904
rect 123354 360848 123359 360904
rect 70228 360846 123359 360848
rect 126838 360906 126898 360982
rect 126973 360906 127039 360909
rect 259453 360906 259519 360909
rect 126838 360904 259519 360906
rect 126838 360848 126978 360904
rect 127034 360848 259458 360904
rect 259514 360848 259519 360904
rect 126838 360846 259519 360848
rect 70228 360844 70234 360846
rect 123293 360843 123359 360846
rect 126973 360843 127039 360846
rect 259453 360843 259519 360846
rect 101489 360226 101555 360229
rect 101949 360226 102015 360229
rect 195329 360226 195395 360229
rect 101489 360224 195395 360226
rect 101489 360168 101494 360224
rect 101550 360168 101954 360224
rect 102010 360168 195334 360224
rect 195390 360168 195395 360224
rect 101489 360166 195395 360168
rect 101489 360163 101555 360166
rect 101949 360163 102015 360166
rect 195329 360163 195395 360166
rect 66110 359348 66116 359412
rect 66180 359410 66186 359412
rect 126973 359410 127039 359413
rect 66180 359408 127039 359410
rect 66180 359352 126978 359408
rect 127034 359352 127039 359408
rect 66180 359350 127039 359352
rect 66180 359348 66186 359350
rect 126973 359347 127039 359350
rect 91185 359276 91251 359277
rect 91134 359274 91140 359276
rect 91094 359214 91140 359274
rect 91204 359272 91251 359276
rect 91246 359216 91251 359272
rect 91134 359212 91140 359214
rect 91204 359212 91251 359216
rect 91185 359211 91251 359212
rect 109534 358940 109540 359004
rect 109604 359002 109610 359004
rect 109677 359002 109743 359005
rect 228357 359002 228423 359005
rect 109604 359000 228423 359002
rect 109604 358944 109682 359000
rect 109738 358944 228362 359000
rect 228418 358944 228423 359000
rect 109604 358942 228423 358944
rect 109604 358940 109610 358942
rect 109677 358939 109743 358942
rect 228357 358939 228423 358942
rect 125593 358866 125659 358869
rect 262213 358866 262279 358869
rect 125593 358864 262279 358866
rect 125593 358808 125598 358864
rect 125654 358808 262218 358864
rect 262274 358808 262279 358864
rect 125593 358806 262279 358808
rect 125593 358803 125659 358806
rect 262213 358803 262279 358806
rect -960 358458 480 358548
rect 3325 358458 3391 358461
rect -960 358456 3391 358458
rect -960 358400 3330 358456
rect 3386 358400 3391 358456
rect -960 358398 3391 358400
rect -960 358308 480 358398
rect 3325 358395 3391 358398
rect 77293 358050 77359 358053
rect 136030 358050 136036 358052
rect 77293 358048 136036 358050
rect 77293 357992 77298 358048
rect 77354 357992 136036 358048
rect 77293 357990 136036 357992
rect 77293 357987 77359 357990
rect 136030 357988 136036 357990
rect 136100 357988 136106 358052
rect 126973 357642 127039 357645
rect 188286 357642 188292 357644
rect 126973 357640 188292 357642
rect 126973 357584 126978 357640
rect 127034 357584 188292 357640
rect 126973 357582 188292 357584
rect 126973 357579 127039 357582
rect 188286 357580 188292 357582
rect 188356 357580 188362 357644
rect 80053 357506 80119 357509
rect 86953 357506 87019 357509
rect 249742 357506 249748 357508
rect 80053 357504 249748 357506
rect 80053 357448 80058 357504
rect 80114 357448 86958 357504
rect 87014 357448 249748 357504
rect 80053 357446 249748 357448
rect 80053 357443 80119 357446
rect 86953 357443 87019 357446
rect 249742 357444 249748 357446
rect 249812 357444 249818 357508
rect 125685 357370 125751 357373
rect 126237 357370 126303 357373
rect 125685 357368 126303 357370
rect 125685 357312 125690 357368
rect 125746 357312 126242 357368
rect 126298 357312 126303 357368
rect 125685 357310 126303 357312
rect 125685 357307 125751 357310
rect 126237 357307 126303 357310
rect 66161 356690 66227 356693
rect 111742 356690 111748 356692
rect 66161 356688 111748 356690
rect 66161 356632 66166 356688
rect 66222 356632 111748 356688
rect 66161 356630 111748 356632
rect 66161 356627 66227 356630
rect 111742 356628 111748 356630
rect 111812 356628 111818 356692
rect 95141 356282 95207 356285
rect 197854 356282 197860 356284
rect 95141 356280 197860 356282
rect 95141 356224 95146 356280
rect 95202 356224 197860 356280
rect 95141 356222 197860 356224
rect 95141 356219 95207 356222
rect 197854 356220 197860 356222
rect 197924 356220 197930 356284
rect 125685 356146 125751 356149
rect 233877 356146 233943 356149
rect 125685 356144 233943 356146
rect 125685 356088 125690 356144
rect 125746 356088 233882 356144
rect 233938 356088 233943 356144
rect 125685 356086 233943 356088
rect 125685 356083 125751 356086
rect 233877 356083 233943 356086
rect 129733 356010 129799 356013
rect 130469 356010 130535 356013
rect 129733 356008 130535 356010
rect 129733 355952 129738 356008
rect 129794 355952 130474 356008
rect 130530 355952 130535 356008
rect 129733 355950 130535 355952
rect 129733 355947 129799 355950
rect 130469 355947 130535 355950
rect 71037 355330 71103 355333
rect 122741 355330 122807 355333
rect 71037 355328 122807 355330
rect 71037 355272 71042 355328
rect 71098 355272 122746 355328
rect 122802 355272 122807 355328
rect 71037 355270 122807 355272
rect 71037 355267 71103 355270
rect 122741 355267 122807 355270
rect 111793 354922 111859 354925
rect 212574 354922 212580 354924
rect 111793 354920 212580 354922
rect 111793 354864 111798 354920
rect 111854 354864 212580 354920
rect 111793 354862 212580 354864
rect 111793 354859 111859 354862
rect 212574 354860 212580 354862
rect 212644 354860 212650 354924
rect 129733 354786 129799 354789
rect 232446 354786 232452 354788
rect 129733 354784 232452 354786
rect 129733 354728 129738 354784
rect 129794 354728 232452 354784
rect 129733 354726 232452 354728
rect 129733 354723 129799 354726
rect 232446 354724 232452 354726
rect 232516 354724 232522 354788
rect 60641 353970 60707 353973
rect 156689 353970 156755 353973
rect 60641 353968 156755 353970
rect 60641 353912 60646 353968
rect 60702 353912 156694 353968
rect 156750 353912 156755 353968
rect 60641 353910 156755 353912
rect 60641 353907 60707 353910
rect 156689 353907 156755 353910
rect 110413 353426 110479 353429
rect 111701 353426 111767 353429
rect 252553 353426 252619 353429
rect 110413 353424 252619 353426
rect 110413 353368 110418 353424
rect 110474 353368 111706 353424
rect 111762 353368 252558 353424
rect 252614 353368 252619 353424
rect 110413 353366 252619 353368
rect 110413 353363 110479 353366
rect 111701 353363 111767 353366
rect 252553 353363 252619 353366
rect 130377 352610 130443 352613
rect 139710 352610 139716 352612
rect 130377 352608 139716 352610
rect 130377 352552 130382 352608
rect 130438 352552 139716 352608
rect 130377 352550 139716 352552
rect 130377 352547 130443 352550
rect 139710 352548 139716 352550
rect 139780 352548 139786 352612
rect 144913 352202 144979 352205
rect 145557 352202 145623 352205
rect 206277 352202 206343 352205
rect 144913 352200 206343 352202
rect 144913 352144 144918 352200
rect 144974 352144 145562 352200
rect 145618 352144 206282 352200
rect 206338 352144 206343 352200
rect 144913 352142 206343 352144
rect 144913 352139 144979 352142
rect 145557 352139 145623 352142
rect 206277 352139 206343 352142
rect 59077 352066 59143 352069
rect 167637 352066 167703 352069
rect 59077 352064 167703 352066
rect 59077 352008 59082 352064
rect 59138 352008 167642 352064
rect 167698 352008 167703 352064
rect 59077 352006 167703 352008
rect 59077 352003 59143 352006
rect 167637 352003 167703 352006
rect 70393 351930 70459 351933
rect 71681 351930 71747 351933
rect 263593 351930 263659 351933
rect 70393 351928 263659 351930
rect 70393 351872 70398 351928
rect 70454 351872 71686 351928
rect 71742 351872 263598 351928
rect 263654 351872 263659 351928
rect 70393 351870 263659 351872
rect 70393 351867 70459 351870
rect 71681 351867 71747 351870
rect 263593 351867 263659 351870
rect 583017 351930 583083 351933
rect 583520 351930 584960 352020
rect 583017 351928 584960 351930
rect 583017 351872 583022 351928
rect 583078 351872 584960 351928
rect 583017 351870 584960 351872
rect 583017 351867 583083 351870
rect 583520 351780 584960 351870
rect 95141 351114 95207 351117
rect 124305 351114 124371 351117
rect 214649 351114 214715 351117
rect 95141 351112 214715 351114
rect 95141 351056 95146 351112
rect 95202 351056 124310 351112
rect 124366 351056 214654 351112
rect 214710 351056 214715 351112
rect 95141 351054 214715 351056
rect 95141 351051 95207 351054
rect 124305 351051 124371 351054
rect 214649 351051 214715 351054
rect 124857 350706 124923 350709
rect 186814 350706 186820 350708
rect 124857 350704 186820 350706
rect 124857 350648 124862 350704
rect 124918 350648 186820 350704
rect 124857 350646 186820 350648
rect 124857 350643 124923 350646
rect 186814 350644 186820 350646
rect 186884 350644 186890 350708
rect 118693 350570 118759 350573
rect 119337 350570 119403 350573
rect 248454 350570 248460 350572
rect 118693 350568 248460 350570
rect 118693 350512 118698 350568
rect 118754 350512 119342 350568
rect 119398 350512 248460 350568
rect 118693 350510 248460 350512
rect 118693 350507 118759 350510
rect 119337 350507 119403 350510
rect 248454 350508 248460 350510
rect 248524 350508 248530 350572
rect 582373 349754 582439 349757
rect 200070 349752 582439 349754
rect 200070 349696 582378 349752
rect 582434 349696 582439 349752
rect 200070 349694 582439 349696
rect 140865 349482 140931 349485
rect 197997 349482 198063 349485
rect 140865 349480 198063 349482
rect 140865 349424 140870 349480
rect 140926 349424 198002 349480
rect 198058 349424 198063 349480
rect 140865 349422 198063 349424
rect 140865 349419 140931 349422
rect 197997 349419 198063 349422
rect 85757 349346 85823 349349
rect 196934 349346 196940 349348
rect 85757 349344 196940 349346
rect 85757 349288 85762 349344
rect 85818 349288 196940 349344
rect 85757 349286 196940 349288
rect 85757 349283 85823 349286
rect 196934 349284 196940 349286
rect 197004 349346 197010 349348
rect 200070 349346 200130 349694
rect 582373 349691 582439 349694
rect 197004 349286 200130 349346
rect 197004 349284 197010 349286
rect 69606 349148 69612 349212
rect 69676 349210 69682 349212
rect 70158 349210 70164 349212
rect 69676 349150 70164 349210
rect 69676 349148 69682 349150
rect 70158 349148 70164 349150
rect 70228 349210 70234 349212
rect 223941 349210 224007 349213
rect 70228 349208 224007 349210
rect 70228 349152 223946 349208
rect 224002 349152 224007 349208
rect 70228 349150 224007 349152
rect 70228 349148 70234 349150
rect 223941 349147 224007 349150
rect 66662 349012 66668 349076
rect 66732 349074 66738 349076
rect 67357 349074 67423 349077
rect 66732 349072 67423 349074
rect 66732 349016 67362 349072
rect 67418 349016 67423 349072
rect 66732 349014 67423 349016
rect 66732 349012 66738 349014
rect 67357 349011 67423 349014
rect 115197 347986 115263 347989
rect 174629 347986 174695 347989
rect 115197 347984 174695 347986
rect 115197 347928 115202 347984
rect 115258 347928 174634 347984
rect 174690 347928 174695 347984
rect 115197 347926 174695 347928
rect 115197 347923 115263 347926
rect 174629 347923 174695 347926
rect 66662 347788 66668 347852
rect 66732 347850 66738 347852
rect 196709 347850 196775 347853
rect 66732 347848 196775 347850
rect 66732 347792 196714 347848
rect 196770 347792 196775 347848
rect 66732 347790 196775 347792
rect 66732 347788 66738 347790
rect 196709 347787 196775 347790
rect 117313 347714 117379 347717
rect 118550 347714 118556 347716
rect 117313 347712 118556 347714
rect 117313 347656 117318 347712
rect 117374 347656 118556 347712
rect 117313 347654 118556 347656
rect 117313 347651 117379 347654
rect 118550 347652 118556 347654
rect 118620 347652 118626 347716
rect 135161 347170 135227 347173
rect 156454 347170 156460 347172
rect 135161 347168 156460 347170
rect 135161 347112 135166 347168
rect 135222 347112 156460 347168
rect 135161 347110 156460 347112
rect 135161 347107 135227 347110
rect 156454 347108 156460 347110
rect 156524 347108 156530 347172
rect 67725 347034 67791 347037
rect 140865 347034 140931 347037
rect 67725 347032 140931 347034
rect 67725 346976 67730 347032
rect 67786 346976 140870 347032
rect 140926 346976 140931 347032
rect 67725 346974 140931 346976
rect 67725 346971 67791 346974
rect 140865 346971 140931 346974
rect 110321 346626 110387 346629
rect 124121 346626 124187 346629
rect 110321 346624 124187 346626
rect 110321 346568 110326 346624
rect 110382 346568 124126 346624
rect 124182 346568 124187 346624
rect 110321 346566 124187 346568
rect 110321 346563 110387 346566
rect 124121 346563 124187 346566
rect 140773 346626 140839 346629
rect 182817 346626 182883 346629
rect 140773 346624 182883 346626
rect 140773 346568 140778 346624
rect 140834 346568 182822 346624
rect 182878 346568 182883 346624
rect 140773 346566 182883 346568
rect 140773 346563 140839 346566
rect 182817 346563 182883 346566
rect 117313 346490 117379 346493
rect 267733 346490 267799 346493
rect 117313 346488 267799 346490
rect 117313 346432 117318 346488
rect 117374 346432 267738 346488
rect 267794 346432 267799 346488
rect 117313 346430 267799 346432
rect 117313 346427 117379 346430
rect 267733 346427 267799 346430
rect 67950 345748 67956 345812
rect 68020 345810 68026 345812
rect 115933 345810 115999 345813
rect 68020 345808 115999 345810
rect 68020 345752 115938 345808
rect 115994 345752 115999 345808
rect 68020 345750 115999 345752
rect 68020 345748 68026 345750
rect 115933 345747 115999 345750
rect 64137 345674 64203 345677
rect 67766 345674 67772 345676
rect 64137 345672 67772 345674
rect 64137 345616 64142 345672
rect 64198 345616 67772 345672
rect 64137 345614 67772 345616
rect 64137 345611 64203 345614
rect 67766 345612 67772 345614
rect 67836 345612 67842 345676
rect 105537 345674 105603 345677
rect 153837 345674 153903 345677
rect 105537 345672 153903 345674
rect 105537 345616 105542 345672
rect 105598 345616 153842 345672
rect 153898 345616 153903 345672
rect 105537 345614 153903 345616
rect 105537 345611 105603 345614
rect 153837 345611 153903 345614
rect -960 345402 480 345492
rect 3141 345402 3207 345405
rect -960 345400 3207 345402
rect -960 345344 3146 345400
rect 3202 345344 3207 345400
rect -960 345342 3207 345344
rect -960 345252 480 345342
rect 3141 345339 3207 345342
rect 122925 345266 122991 345269
rect 191097 345266 191163 345269
rect 122925 345264 191163 345266
rect 122925 345208 122930 345264
rect 122986 345208 191102 345264
rect 191158 345208 191163 345264
rect 122925 345206 191163 345208
rect 122925 345203 122991 345206
rect 191097 345203 191163 345206
rect 118601 345130 118667 345133
rect 357433 345130 357499 345133
rect 118601 345128 357499 345130
rect 118601 345072 118606 345128
rect 118662 345072 357438 345128
rect 357494 345072 357499 345128
rect 118601 345070 357499 345072
rect 118601 345067 118667 345070
rect 357433 345067 357499 345070
rect 121361 343906 121427 343909
rect 173157 343906 173223 343909
rect 121361 343904 173223 343906
rect 121361 343848 121366 343904
rect 121422 343848 173162 343904
rect 173218 343848 173223 343904
rect 121361 343846 173223 343848
rect 121361 343843 121427 343846
rect 173157 343843 173223 343846
rect 108941 343770 109007 343773
rect 582373 343770 582439 343773
rect 108941 343768 582439 343770
rect 108941 343712 108946 343768
rect 109002 343712 582378 343768
rect 582434 343712 582439 343768
rect 108941 343710 582439 343712
rect 108941 343707 109007 343710
rect 582373 343707 582439 343710
rect 139301 342546 139367 342549
rect 160185 342546 160251 342549
rect 139301 342544 160251 342546
rect 139301 342488 139306 342544
rect 139362 342488 160190 342544
rect 160246 342488 160251 342544
rect 139301 342486 160251 342488
rect 139301 342483 139367 342486
rect 160185 342483 160251 342486
rect 116577 342410 116643 342413
rect 176009 342410 176075 342413
rect 116577 342408 176075 342410
rect 116577 342352 116582 342408
rect 116638 342352 176014 342408
rect 176070 342352 176075 342408
rect 116577 342350 176075 342352
rect 116577 342347 116643 342350
rect 176009 342347 176075 342350
rect 70117 342274 70183 342277
rect 200757 342274 200823 342277
rect 70117 342272 200823 342274
rect 70117 342216 70122 342272
rect 70178 342216 200762 342272
rect 200818 342216 200823 342272
rect 70117 342214 200823 342216
rect 70117 342211 70183 342214
rect 200757 342211 200823 342214
rect 67265 341186 67331 341189
rect 178677 341186 178743 341189
rect 67265 341184 178743 341186
rect 67265 341128 67270 341184
rect 67326 341128 178682 341184
rect 178738 341128 178743 341184
rect 67265 341126 178743 341128
rect 67265 341123 67331 341126
rect 178677 341123 178743 341126
rect 80697 341050 80763 341053
rect 230422 341050 230428 341052
rect 80697 341048 230428 341050
rect 80697 340992 80702 341048
rect 80758 340992 230428 341048
rect 80697 340990 230428 340992
rect 80697 340987 80763 340990
rect 230422 340988 230428 340990
rect 230492 340988 230498 341052
rect 111701 340914 111767 340917
rect 335997 340914 336063 340917
rect 111701 340912 336063 340914
rect 111701 340856 111706 340912
rect 111762 340856 336002 340912
rect 336058 340856 336063 340912
rect 111701 340854 336063 340856
rect 111701 340851 111767 340854
rect 335997 340851 336063 340854
rect 142061 339826 142127 339829
rect 187049 339826 187115 339829
rect 142061 339824 187115 339826
rect 142061 339768 142066 339824
rect 142122 339768 187054 339824
rect 187110 339768 187115 339824
rect 142061 339766 187115 339768
rect 142061 339763 142127 339766
rect 187049 339763 187115 339766
rect 73061 339690 73127 339693
rect 209129 339690 209195 339693
rect 73061 339688 209195 339690
rect 73061 339632 73066 339688
rect 73122 339632 209134 339688
rect 209190 339632 209195 339688
rect 73061 339630 209195 339632
rect 73061 339627 73127 339630
rect 209129 339627 209195 339630
rect 98637 339554 98703 339557
rect 291142 339554 291148 339556
rect 98637 339552 291148 339554
rect 98637 339496 98642 339552
rect 98698 339496 291148 339552
rect 98637 339494 291148 339496
rect 98637 339491 98703 339494
rect 291142 339492 291148 339494
rect 291212 339492 291218 339556
rect 82721 338738 82787 338741
rect 109677 338738 109743 338741
rect 82721 338736 109743 338738
rect 82721 338680 82726 338736
rect 82782 338680 109682 338736
rect 109738 338680 109743 338736
rect 82721 338678 109743 338680
rect 82721 338675 82787 338678
rect 109677 338675 109743 338678
rect 120717 338466 120783 338469
rect 171869 338466 171935 338469
rect 120717 338464 171935 338466
rect 120717 338408 120722 338464
rect 120778 338408 171874 338464
rect 171930 338408 171935 338464
rect 583520 338452 584960 338692
rect 120717 338406 171935 338408
rect 120717 338403 120783 338406
rect 171869 338403 171935 338406
rect 64689 338330 64755 338333
rect 165061 338330 165127 338333
rect 64689 338328 165127 338330
rect 64689 338272 64694 338328
rect 64750 338272 165066 338328
rect 165122 338272 165127 338328
rect 64689 338270 165127 338272
rect 64689 338267 64755 338270
rect 165061 338267 165127 338270
rect 106181 338194 106247 338197
rect 222837 338194 222903 338197
rect 106181 338192 222903 338194
rect 106181 338136 106186 338192
rect 106242 338136 222842 338192
rect 222898 338136 222903 338192
rect 106181 338134 222903 338136
rect 106181 338131 106247 338134
rect 222837 338131 222903 338134
rect 87137 337106 87203 337109
rect 216029 337106 216095 337109
rect 87137 337104 216095 337106
rect 87137 337048 87142 337104
rect 87198 337048 216034 337104
rect 216090 337048 216095 337104
rect 87137 337046 216095 337048
rect 87137 337043 87203 337046
rect 216029 337043 216095 337046
rect 88609 336970 88675 336973
rect 220169 336970 220235 336973
rect 88609 336968 220235 336970
rect 88609 336912 88614 336968
rect 88670 336912 220174 336968
rect 220230 336912 220235 336968
rect 88609 336910 220235 336912
rect 88609 336907 88675 336910
rect 220169 336907 220235 336910
rect 74625 336834 74691 336837
rect 313917 336834 313983 336837
rect 74625 336832 313983 336834
rect 74625 336776 74630 336832
rect 74686 336776 313922 336832
rect 313978 336776 313983 336832
rect 74625 336774 313983 336776
rect 74625 336771 74691 336774
rect 313917 336771 313983 336774
rect 160185 336018 160251 336021
rect 239397 336018 239463 336021
rect 160185 336016 239463 336018
rect 160185 335960 160190 336016
rect 160246 335960 239402 336016
rect 239458 335960 239463 336016
rect 160185 335958 239463 335960
rect 160185 335955 160251 335958
rect 239397 335955 239463 335958
rect 135253 335746 135319 335749
rect 162301 335746 162367 335749
rect 135253 335744 162367 335746
rect 135253 335688 135258 335744
rect 135314 335688 162306 335744
rect 162362 335688 162367 335744
rect 135253 335686 162367 335688
rect 135253 335683 135319 335686
rect 162301 335683 162367 335686
rect 89805 335610 89871 335613
rect 166533 335610 166599 335613
rect 89805 335608 166599 335610
rect 89805 335552 89810 335608
rect 89866 335552 166538 335608
rect 166594 335552 166599 335608
rect 89805 335550 166599 335552
rect 89805 335547 89871 335550
rect 166533 335547 166599 335550
rect 60457 335474 60523 335477
rect 159541 335474 159607 335477
rect 60457 335472 159607 335474
rect 60457 335416 60462 335472
rect 60518 335416 159546 335472
rect 159602 335416 159607 335472
rect 60457 335414 159607 335416
rect 60457 335411 60523 335414
rect 159541 335411 159607 335414
rect 73705 334386 73771 334389
rect 189717 334386 189783 334389
rect 73705 334384 189783 334386
rect 73705 334328 73710 334384
rect 73766 334328 189722 334384
rect 189778 334328 189783 334384
rect 73705 334326 189783 334328
rect 73705 334323 73771 334326
rect 189717 334323 189783 334326
rect 71405 334250 71471 334253
rect 207657 334250 207723 334253
rect 71405 334248 207723 334250
rect 71405 334192 71410 334248
rect 71466 334192 207662 334248
rect 207718 334192 207723 334248
rect 71405 334190 207723 334192
rect 71405 334187 71471 334190
rect 207657 334187 207723 334190
rect 125317 334114 125383 334117
rect 339493 334114 339559 334117
rect 125317 334112 339559 334114
rect 125317 334056 125322 334112
rect 125378 334056 339498 334112
rect 339554 334056 339559 334112
rect 125317 334054 339559 334056
rect 125317 334051 125383 334054
rect 339493 334051 339559 334054
rect 97165 332890 97231 332893
rect 178953 332890 179019 332893
rect 97165 332888 179019 332890
rect 97165 332832 97170 332888
rect 97226 332832 178958 332888
rect 179014 332832 179019 332888
rect 97165 332830 179019 332832
rect 97165 332827 97231 332830
rect 178953 332827 179019 332830
rect 70669 332754 70735 332757
rect 208485 332754 208551 332757
rect 70669 332752 208551 332754
rect 70669 332696 70674 332752
rect 70730 332696 208490 332752
rect 208546 332696 208551 332752
rect 70669 332694 208551 332696
rect 70669 332691 70735 332694
rect 208485 332691 208551 332694
rect 77937 332618 78003 332621
rect 324313 332618 324379 332621
rect 77937 332616 324379 332618
rect 77937 332560 77942 332616
rect 77998 332560 324318 332616
rect 324374 332560 324379 332616
rect 77937 332558 324379 332560
rect 77937 332555 78003 332558
rect 324313 332555 324379 332558
rect 92381 332482 92447 332485
rect 93894 332482 93900 332484
rect 92381 332480 93900 332482
rect -960 332196 480 332436
rect 92381 332424 92386 332480
rect 92442 332424 93900 332480
rect 92381 332422 93900 332424
rect 92381 332419 92447 332422
rect 93894 332420 93900 332422
rect 93964 332420 93970 332484
rect 64781 331802 64847 331805
rect 135897 331802 135963 331805
rect 64781 331800 135963 331802
rect 64781 331744 64786 331800
rect 64842 331744 135902 331800
rect 135958 331744 135963 331800
rect 64781 331742 135963 331744
rect 64781 331739 64847 331742
rect 135897 331739 135963 331742
rect 136909 331530 136975 331533
rect 160686 331530 160692 331532
rect 136909 331528 160692 331530
rect 136909 331472 136914 331528
rect 136970 331472 160692 331528
rect 136909 331470 160692 331472
rect 136909 331467 136975 331470
rect 160686 331468 160692 331470
rect 160756 331468 160762 331532
rect 140865 331394 140931 331397
rect 226425 331394 226491 331397
rect 140865 331392 226491 331394
rect 140865 331336 140870 331392
rect 140926 331336 226430 331392
rect 226486 331336 226491 331392
rect 140865 331334 226491 331336
rect 140865 331331 140931 331334
rect 226425 331331 226491 331334
rect 92841 331258 92907 331261
rect 217317 331258 217383 331261
rect 92841 331256 217383 331258
rect 92841 331200 92846 331256
rect 92902 331200 217322 331256
rect 217378 331200 217383 331256
rect 92841 331198 217383 331200
rect 92841 331195 92907 331198
rect 217317 331195 217383 331198
rect 53833 331122 53899 331125
rect 54937 331122 55003 331125
rect 100109 331122 100175 331125
rect 53833 331120 100175 331122
rect 53833 331064 53838 331120
rect 53894 331064 54942 331120
rect 54998 331064 100114 331120
rect 100170 331064 100175 331120
rect 53833 331062 100175 331064
rect 53833 331059 53899 331062
rect 54937 331059 55003 331062
rect 100109 331059 100175 331062
rect 95049 330714 95115 330717
rect 108297 330714 108363 330717
rect 95049 330712 108363 330714
rect 95049 330656 95054 330712
rect 95110 330656 108302 330712
rect 108358 330656 108363 330712
rect 95049 330654 108363 330656
rect 95049 330651 95115 330654
rect 108297 330651 108363 330654
rect 99281 330578 99347 330581
rect 120717 330578 120783 330581
rect 99281 330576 120783 330578
rect 99281 330520 99286 330576
rect 99342 330520 120722 330576
rect 120778 330520 120783 330576
rect 99281 330518 120783 330520
rect 99281 330515 99347 330518
rect 120717 330515 120783 330518
rect 17217 330442 17283 330445
rect 53833 330442 53899 330445
rect 17217 330440 53899 330442
rect 17217 330384 17222 330440
rect 17278 330384 53838 330440
rect 53894 330384 53899 330440
rect 17217 330382 53899 330384
rect 17217 330379 17283 330382
rect 53833 330379 53899 330382
rect 97809 330442 97875 330445
rect 98637 330442 98703 330445
rect 140865 330442 140931 330445
rect 97809 330440 98703 330442
rect 97809 330384 97814 330440
rect 97870 330384 98642 330440
rect 98698 330384 98703 330440
rect 97809 330382 98703 330384
rect 97809 330379 97875 330382
rect 98637 330379 98703 330382
rect 103470 330440 140931 330442
rect 103470 330384 140870 330440
rect 140926 330384 140931 330440
rect 103470 330382 140931 330384
rect 98545 330306 98611 330309
rect 103470 330306 103530 330382
rect 140865 330379 140931 330382
rect 178677 330442 178743 330445
rect 230381 330442 230447 330445
rect 178677 330440 230447 330442
rect 178677 330384 178682 330440
rect 178738 330384 230386 330440
rect 230442 330384 230447 330440
rect 178677 330382 230447 330384
rect 178677 330379 178743 330382
rect 230381 330379 230447 330382
rect 98545 330304 103530 330306
rect 98545 330248 98550 330304
rect 98606 330248 103530 330304
rect 98545 330246 103530 330248
rect 98545 330243 98611 330246
rect 142889 330170 142955 330173
rect 174537 330170 174603 330173
rect 142889 330168 174603 330170
rect 142889 330112 142894 330168
rect 142950 330112 174542 330168
rect 174598 330112 174603 330168
rect 142889 330110 174603 330112
rect 142889 330107 142955 330110
rect 174537 330107 174603 330110
rect 61878 329972 61884 330036
rect 61948 330034 61954 330036
rect 88425 330034 88491 330037
rect 61948 330032 88491 330034
rect 61948 329976 88430 330032
rect 88486 329976 88491 330032
rect 61948 329974 88491 329976
rect 61948 329972 61954 329974
rect 88425 329971 88491 329974
rect 112805 330034 112871 330037
rect 154246 330034 154252 330036
rect 112805 330032 154252 330034
rect 112805 329976 112810 330032
rect 112866 329976 154252 330032
rect 112805 329974 154252 329976
rect 112805 329971 112871 329974
rect 154246 329972 154252 329974
rect 154316 329972 154322 330036
rect 131481 329898 131547 329901
rect 198089 329898 198155 329901
rect 131481 329896 198155 329898
rect 131481 329840 131486 329896
rect 131542 329840 198094 329896
rect 198150 329840 198155 329896
rect 131481 329838 198155 329840
rect 131481 329835 131547 329838
rect 198089 329835 198155 329838
rect 140773 329082 140839 329085
rect 202781 329082 202847 329085
rect 140773 329080 202847 329082
rect 140773 329024 140778 329080
rect 140834 329024 202786 329080
rect 202842 329024 202847 329080
rect 140773 329022 202847 329024
rect 140773 329019 140839 329022
rect 202781 329019 202847 329022
rect 135253 328946 135319 328949
rect 163681 328946 163747 328949
rect 135253 328944 163747 328946
rect 135253 328888 135258 328944
rect 135314 328888 163686 328944
rect 163742 328888 163747 328944
rect 135253 328886 163747 328888
rect 135253 328883 135319 328886
rect 163681 328883 163747 328886
rect 122097 328810 122163 328813
rect 140773 328810 140839 328813
rect 122097 328808 140839 328810
rect 122097 328752 122102 328808
rect 122158 328752 140778 328808
rect 140834 328752 140839 328808
rect 122097 328750 140839 328752
rect 122097 328747 122163 328750
rect 140773 328747 140839 328750
rect 68001 328674 68067 328677
rect 139761 328674 139827 328677
rect 68001 328672 139827 328674
rect 68001 328616 68006 328672
rect 68062 328616 139766 328672
rect 139822 328616 139827 328672
rect 68001 328614 139827 328616
rect 68001 328611 68067 328614
rect 139761 328611 139827 328614
rect 7557 328538 7623 328541
rect 123477 328538 123543 328541
rect 7557 328536 123543 328538
rect 7557 328480 7562 328536
rect 7618 328480 123482 328536
rect 123538 328480 123543 328536
rect 7557 328478 123543 328480
rect 7557 328475 7623 328478
rect 123477 328475 123543 328478
rect 148317 328538 148383 328541
rect 156229 328538 156295 328541
rect 148317 328536 156295 328538
rect 148317 328480 148322 328536
rect 148378 328480 156234 328536
rect 156290 328480 156295 328536
rect 148317 328478 156295 328480
rect 148317 328475 148383 328478
rect 156229 328475 156295 328478
rect 140773 327858 140839 327861
rect 159357 327858 159423 327861
rect 140773 327856 159423 327858
rect 140773 327800 140778 327856
rect 140834 327800 159362 327856
rect 159418 327800 159423 327856
rect 140773 327798 159423 327800
rect 140773 327795 140839 327798
rect 159357 327795 159423 327798
rect 111885 327722 111951 327725
rect 153694 327722 153700 327724
rect 111885 327720 153700 327722
rect 111885 327664 111890 327720
rect 111946 327664 153700 327720
rect 111885 327662 153700 327664
rect 111885 327659 111951 327662
rect 153694 327660 153700 327662
rect 153764 327660 153770 327724
rect 77293 327586 77359 327589
rect 78213 327586 78279 327589
rect 77293 327584 78279 327586
rect 77293 327528 77298 327584
rect 77354 327528 78218 327584
rect 78274 327528 78279 327584
rect 77293 327526 78279 327528
rect 77293 327523 77359 327526
rect 78213 327523 78279 327526
rect 82670 327524 82676 327588
rect 82740 327586 82746 327588
rect 82997 327586 83063 327589
rect 82740 327584 83063 327586
rect 82740 327528 83002 327584
rect 83058 327528 83063 327584
rect 82740 327526 83063 327528
rect 82740 327524 82746 327526
rect 82997 327523 83063 327526
rect 78581 327314 78647 327317
rect 212901 327314 212967 327317
rect 78581 327312 212967 327314
rect 78581 327256 78586 327312
rect 78642 327256 212906 327312
rect 212962 327256 212967 327312
rect 78581 327254 212967 327256
rect 78581 327251 78647 327254
rect 212901 327251 212967 327254
rect 145598 327116 145604 327180
rect 145668 327178 145674 327180
rect 147213 327178 147279 327181
rect 145668 327176 147279 327178
rect 145668 327120 147218 327176
rect 147274 327120 147279 327176
rect 145668 327118 147279 327120
rect 145668 327116 145674 327118
rect 147213 327115 147279 327118
rect 150382 327116 150388 327180
rect 150452 327178 150458 327180
rect 150709 327178 150775 327181
rect 150452 327176 150775 327178
rect 150452 327120 150714 327176
rect 150770 327120 150775 327176
rect 150452 327118 150775 327120
rect 150452 327116 150458 327118
rect 150709 327115 150775 327118
rect 153653 327178 153719 327181
rect 155350 327178 155356 327180
rect 153653 327176 155356 327178
rect 153653 327120 153658 327176
rect 153714 327120 155356 327176
rect 153653 327118 155356 327120
rect 153653 327115 153719 327118
rect 155350 327116 155356 327118
rect 155420 327116 155426 327180
rect 67265 327042 67331 327045
rect 67398 327042 67404 327044
rect 67265 327040 67404 327042
rect 67265 326984 67270 327040
rect 67326 326984 67404 327040
rect 67265 326982 67404 326984
rect 67265 326979 67331 326982
rect 67398 326980 67404 326982
rect 67468 326980 67474 327044
rect 70025 327042 70091 327045
rect 69430 327040 70091 327042
rect 69430 326984 70030 327040
rect 70086 326984 70091 327040
rect 69430 326982 70091 326984
rect 68093 326770 68159 326773
rect 69430 326770 69490 326982
rect 70025 326979 70091 326982
rect 154205 327042 154271 327045
rect 333973 327042 334039 327045
rect 154205 327040 334039 327042
rect 154205 326984 154210 327040
rect 154266 326984 333978 327040
rect 334034 326984 334039 327040
rect 154205 326982 334039 326984
rect 154205 326979 154271 326982
rect 333973 326979 334039 326982
rect 68093 326768 69490 326770
rect 68093 326712 68098 326768
rect 68154 326740 69490 326768
rect 68154 326712 69460 326740
rect 68093 326710 69460 326712
rect 68093 326707 68159 326710
rect 68645 326498 68711 326501
rect 160870 326498 160876 326500
rect 68645 326496 68938 326498
rect 68645 326440 68650 326496
rect 68706 326440 68938 326496
rect 68645 326438 68938 326440
rect 154652 326438 160876 326498
rect 68645 326435 68711 326438
rect 68878 325924 68938 326438
rect 160870 326436 160876 326438
rect 160940 326436 160946 326500
rect 156045 325410 156111 325413
rect 154652 325408 156111 325410
rect 154652 325352 156050 325408
rect 156106 325352 156111 325408
rect 154652 325350 156111 325352
rect 156045 325347 156111 325350
rect 582833 325274 582899 325277
rect 583520 325274 584960 325364
rect 582833 325272 584960 325274
rect 582833 325216 582838 325272
rect 582894 325216 584960 325272
rect 582833 325214 584960 325216
rect 582833 325211 582899 325214
rect 583520 325124 584960 325214
rect 154849 325002 154915 325005
rect 237414 325002 237420 325004
rect 154849 325000 237420 325002
rect 154849 324944 154854 325000
rect 154910 324944 237420 325000
rect 154849 324942 237420 324944
rect 154849 324939 154915 324942
rect 237414 324940 237420 324942
rect 237484 324940 237490 325004
rect 66897 324866 66963 324869
rect 66897 324864 68908 324866
rect 66897 324808 66902 324864
rect 66958 324808 68908 324864
rect 66897 324806 68908 324808
rect 66897 324803 66963 324806
rect 156045 324322 156111 324325
rect 154652 324320 156111 324322
rect 154652 324264 156050 324320
rect 156106 324264 156111 324320
rect 154652 324262 156111 324264
rect 156045 324259 156111 324262
rect 66713 323778 66779 323781
rect 66713 323776 68908 323778
rect 66713 323720 66718 323776
rect 66774 323720 68908 323776
rect 66713 323718 68908 323720
rect 66713 323715 66779 323718
rect 156137 323234 156203 323237
rect 154652 323232 156203 323234
rect 154652 323176 156142 323232
rect 156198 323176 156203 323232
rect 154652 323174 156203 323176
rect 156137 323171 156203 323174
rect 67173 322690 67239 322693
rect 67173 322688 68908 322690
rect 67173 322632 67178 322688
rect 67234 322632 68908 322688
rect 67173 322630 68908 322632
rect 67173 322627 67239 322630
rect 156045 322146 156111 322149
rect 154652 322144 156111 322146
rect 154652 322088 156050 322144
rect 156106 322088 156111 322144
rect 154652 322086 156111 322088
rect 156045 322083 156111 322086
rect 159541 322146 159607 322149
rect 199469 322146 199535 322149
rect 159541 322144 199535 322146
rect 159541 322088 159546 322144
rect 159602 322088 199474 322144
rect 199530 322088 199535 322144
rect 159541 322086 199535 322088
rect 159541 322083 159607 322086
rect 199469 322083 199535 322086
rect 67817 321602 67883 321605
rect 67817 321600 68908 321602
rect 67817 321544 67822 321600
rect 67878 321544 68908 321600
rect 67817 321542 68908 321544
rect 67817 321539 67883 321542
rect 156597 321058 156663 321061
rect 154652 321056 156663 321058
rect 154652 321000 156602 321056
rect 156658 321000 156663 321056
rect 154652 320998 156663 321000
rect 156597 320995 156663 320998
rect 154246 320724 154252 320788
rect 154316 320786 154322 320788
rect 178677 320786 178743 320789
rect 154316 320784 178743 320786
rect 154316 320728 178682 320784
rect 178738 320728 178743 320784
rect 154316 320726 178743 320728
rect 154316 320724 154322 320726
rect 178677 320723 178743 320726
rect 66621 320514 66687 320517
rect 66621 320512 68908 320514
rect 66621 320456 66626 320512
rect 66682 320456 68908 320512
rect 66621 320454 68908 320456
rect 66621 320451 66687 320454
rect 157241 319970 157307 319973
rect 154652 319968 157307 319970
rect 154652 319912 157246 319968
rect 157302 319912 157307 319968
rect 154652 319910 157307 319912
rect 157241 319907 157307 319910
rect 66897 319426 66963 319429
rect 195145 319426 195211 319429
rect 309133 319426 309199 319429
rect 66897 319424 68908 319426
rect -960 319290 480 319380
rect 66897 319368 66902 319424
rect 66958 319368 68908 319424
rect 66897 319366 68908 319368
rect 195145 319424 309199 319426
rect 195145 319368 195150 319424
rect 195206 319368 309138 319424
rect 309194 319368 309199 319424
rect 195145 319366 309199 319368
rect 66897 319363 66963 319366
rect 195145 319363 195211 319366
rect 309133 319363 309199 319366
rect 4061 319290 4127 319293
rect -960 319288 4127 319290
rect -960 319232 4066 319288
rect 4122 319232 4127 319288
rect -960 319230 4127 319232
rect -960 319140 480 319230
rect 4061 319227 4127 319230
rect 157241 318882 157307 318885
rect 154652 318880 157307 318882
rect 154652 318824 157246 318880
rect 157302 318824 157307 318880
rect 154652 318822 157307 318824
rect 157241 318819 157307 318822
rect 155166 318610 155172 318612
rect 154622 318550 155172 318610
rect 66713 318338 66779 318341
rect 66713 318336 68908 318338
rect 66713 318280 66718 318336
rect 66774 318280 68908 318336
rect 66713 318278 68908 318280
rect 66713 318275 66779 318278
rect 154622 318036 154682 318550
rect 155166 318548 155172 318550
rect 155236 318610 155242 318612
rect 156597 318610 156663 318613
rect 155236 318608 156663 318610
rect 155236 318552 156602 318608
rect 156658 318552 156663 318608
rect 155236 318550 156663 318552
rect 155236 318548 155242 318550
rect 156597 318547 156663 318550
rect 155350 318140 155356 318204
rect 155420 318202 155426 318204
rect 155420 318142 161490 318202
rect 155420 318140 155426 318142
rect 161430 318066 161490 318142
rect 332593 318066 332659 318069
rect 161430 318064 332659 318066
rect 161430 318008 332598 318064
rect 332654 318008 332659 318064
rect 161430 318006 332659 318008
rect 332593 318003 332659 318006
rect 66897 317522 66963 317525
rect 66897 317520 68908 317522
rect 66897 317464 66902 317520
rect 66958 317464 68908 317520
rect 66897 317462 68908 317464
rect 66897 317459 66963 317462
rect 191189 317386 191255 317389
rect 191598 317386 191604 317388
rect 191189 317384 191604 317386
rect 191189 317328 191194 317384
rect 191250 317328 191604 317384
rect 191189 317326 191604 317328
rect 191189 317323 191255 317326
rect 191598 317324 191604 317326
rect 191668 317324 191674 317388
rect 157241 316978 157307 316981
rect 154652 316976 157307 316978
rect 154652 316920 157246 316976
rect 157302 316920 157307 316976
rect 154652 316918 157307 316920
rect 157241 316915 157307 316918
rect 66662 316372 66668 316436
rect 66732 316434 66738 316436
rect 66732 316374 68908 316434
rect 66732 316372 66738 316374
rect 191598 316100 191604 316164
rect 191668 316162 191674 316164
rect 256693 316162 256759 316165
rect 191668 316160 256759 316162
rect 191668 316104 256698 316160
rect 256754 316104 256759 316160
rect 191668 316102 256759 316104
rect 191668 316100 191674 316102
rect 256693 316099 256759 316102
rect 157241 315890 157307 315893
rect 154652 315888 157307 315890
rect 154652 315832 157246 315888
rect 157302 315832 157307 315888
rect 154652 315830 157307 315832
rect 157241 315827 157307 315830
rect 69422 315556 69428 315620
rect 69492 315556 69498 315620
rect 67541 315346 67607 315349
rect 69430 315346 69490 315556
rect 67541 315344 69490 315346
rect 67541 315288 67546 315344
rect 67602 315316 69490 315344
rect 167637 315346 167703 315349
rect 211889 315346 211955 315349
rect 167637 315344 211955 315346
rect 67602 315288 69460 315316
rect 67541 315286 69460 315288
rect 167637 315288 167642 315344
rect 167698 315288 211894 315344
rect 211950 315288 211955 315344
rect 167637 315286 211955 315288
rect 67541 315283 67607 315286
rect 167637 315283 167703 315286
rect 211889 315283 211955 315286
rect 154246 315012 154252 315076
rect 154316 315074 154322 315076
rect 160921 315074 160987 315077
rect 154316 315072 160987 315074
rect 154316 315016 160926 315072
rect 160982 315016 160987 315072
rect 154316 315014 160987 315016
rect 154316 315012 154322 315014
rect 160921 315011 160987 315014
rect 155953 314802 156019 314805
rect 154652 314800 156019 314802
rect 154652 314744 155958 314800
rect 156014 314744 156019 314800
rect 154652 314742 156019 314744
rect 155953 314739 156019 314742
rect 65517 314258 65583 314261
rect 65517 314256 68908 314258
rect 65517 314200 65522 314256
rect 65578 314200 68908 314256
rect 65517 314198 68908 314200
rect 65517 314195 65583 314198
rect 160686 313924 160692 313988
rect 160756 313986 160762 313988
rect 327073 313986 327139 313989
rect 160756 313984 327139 313986
rect 160756 313928 327078 313984
rect 327134 313928 327139 313984
rect 160756 313926 327139 313928
rect 160756 313924 160762 313926
rect 327073 313923 327139 313926
rect 154622 313306 154682 313684
rect 195094 313306 195100 313308
rect 154622 313246 195100 313306
rect 195094 313244 195100 313246
rect 195164 313244 195170 313308
rect 66897 313170 66963 313173
rect 66897 313168 68908 313170
rect 66897 313112 66902 313168
rect 66958 313112 68908 313168
rect 66897 313110 68908 313112
rect 66897 313107 66963 313110
rect 157241 312626 157307 312629
rect 154652 312624 157307 312626
rect 154652 312568 157246 312624
rect 157302 312568 157307 312624
rect 154652 312566 157307 312568
rect 157241 312563 157307 312566
rect 67725 312082 67791 312085
rect 583385 312082 583451 312085
rect 583520 312082 584960 312172
rect 67725 312080 68908 312082
rect 67725 312024 67730 312080
rect 67786 312024 68908 312080
rect 67725 312022 68908 312024
rect 583385 312080 584960 312082
rect 583385 312024 583390 312080
rect 583446 312024 584960 312080
rect 583385 312022 584960 312024
rect 67725 312019 67791 312022
rect 583385 312019 583451 312022
rect 215845 311946 215911 311949
rect 216029 311946 216095 311949
rect 284334 311946 284340 311948
rect 215845 311944 284340 311946
rect 215845 311888 215850 311944
rect 215906 311888 216034 311944
rect 216090 311888 284340 311944
rect 215845 311886 284340 311888
rect 215845 311883 215911 311886
rect 216029 311883 216095 311886
rect 284334 311884 284340 311886
rect 284404 311884 284410 311948
rect 583520 311932 584960 312022
rect 157241 311538 157307 311541
rect 154652 311536 157307 311538
rect 154652 311480 157246 311536
rect 157302 311480 157307 311536
rect 154652 311478 157307 311480
rect 157241 311475 157307 311478
rect 160870 311068 160876 311132
rect 160940 311130 160946 311132
rect 338113 311130 338179 311133
rect 160940 311128 338179 311130
rect 160940 311072 338118 311128
rect 338174 311072 338179 311128
rect 160940 311070 338179 311072
rect 160940 311068 160946 311070
rect 338113 311067 338179 311070
rect 66897 310994 66963 310997
rect 66897 310992 68908 310994
rect 66897 310936 66902 310992
rect 66958 310936 68908 310992
rect 66897 310934 68908 310936
rect 66897 310931 66963 310934
rect 227621 310586 227687 310589
rect 266997 310586 267063 310589
rect 227621 310584 267063 310586
rect 227621 310528 227626 310584
rect 227682 310528 267002 310584
rect 267058 310528 267063 310584
rect 227621 310526 267063 310528
rect 227621 310523 227687 310526
rect 266997 310523 267063 310526
rect 157241 310450 157307 310453
rect 154652 310448 157307 310450
rect 154652 310392 157246 310448
rect 157302 310392 157307 310448
rect 154652 310390 157307 310392
rect 157241 310387 157307 310390
rect 66621 309906 66687 309909
rect 66621 309904 68908 309906
rect 66621 309848 66626 309904
rect 66682 309848 68908 309904
rect 66621 309846 68908 309848
rect 66621 309843 66687 309846
rect 157149 309634 157215 309637
rect 154652 309632 157215 309634
rect 154652 309576 157154 309632
rect 157210 309576 157215 309632
rect 154652 309574 157215 309576
rect 157149 309571 157215 309574
rect 157241 309226 157307 309229
rect 316033 309226 316099 309229
rect 157241 309224 316099 309226
rect 157241 309168 157246 309224
rect 157302 309168 316038 309224
rect 316094 309168 316099 309224
rect 157241 309166 316099 309168
rect 157241 309163 157307 309166
rect 316033 309163 316099 309166
rect 67081 309090 67147 309093
rect 67449 309090 67515 309093
rect 67081 309088 68908 309090
rect 67081 309032 67086 309088
rect 67142 309032 67454 309088
rect 67510 309032 68908 309088
rect 67081 309030 68908 309032
rect 67081 309027 67147 309030
rect 67449 309027 67515 309030
rect 156137 308546 156203 308549
rect 186998 308546 187004 308548
rect 154652 308544 187004 308546
rect 154652 308488 156142 308544
rect 156198 308488 187004 308544
rect 154652 308486 187004 308488
rect 156137 308483 156203 308486
rect 186998 308484 187004 308486
rect 187068 308484 187074 308548
rect 157149 308410 157215 308413
rect 214230 308410 214236 308412
rect 157149 308408 214236 308410
rect 157149 308352 157154 308408
rect 157210 308352 214236 308408
rect 157149 308350 214236 308352
rect 157149 308347 157215 308350
rect 214230 308348 214236 308350
rect 214300 308348 214306 308412
rect 67081 308002 67147 308005
rect 67398 308002 67404 308004
rect 67081 308000 67404 308002
rect 67081 307944 67086 308000
rect 67142 307944 67404 308000
rect 67081 307942 67404 307944
rect 67081 307939 67147 307942
rect 67398 307940 67404 307942
rect 67468 308002 67474 308004
rect 67468 307942 68908 308002
rect 67468 307940 67474 307942
rect 158069 307866 158135 307869
rect 249885 307866 249951 307869
rect 158069 307864 249951 307866
rect 158069 307808 158074 307864
rect 158130 307808 249890 307864
rect 249946 307808 249951 307864
rect 158069 307806 249951 307808
rect 158069 307803 158135 307806
rect 249885 307803 249951 307806
rect 156505 307458 156571 307461
rect 154652 307456 156571 307458
rect 154652 307400 156510 307456
rect 156566 307400 156571 307456
rect 154652 307398 156571 307400
rect 156505 307395 156571 307398
rect 66529 306914 66595 306917
rect 66529 306912 68908 306914
rect 66529 306856 66534 306912
rect 66590 306856 68908 306912
rect 66529 306854 68908 306856
rect 66529 306851 66595 306854
rect 170581 306506 170647 306509
rect 242934 306506 242940 306508
rect 170581 306504 242940 306506
rect 170581 306448 170586 306504
rect 170642 306448 242940 306504
rect 170581 306446 242940 306448
rect 170581 306443 170647 306446
rect 242934 306444 242940 306446
rect 243004 306444 243010 306508
rect 157241 306370 157307 306373
rect 154652 306368 157307 306370
rect -960 306234 480 306324
rect 154652 306312 157246 306368
rect 157302 306312 157307 306368
rect 154652 306310 157307 306312
rect 157241 306307 157307 306310
rect 3509 306234 3575 306237
rect -960 306232 3575 306234
rect -960 306176 3514 306232
rect 3570 306176 3575 306232
rect -960 306174 3575 306176
rect -960 306084 480 306174
rect 3509 306171 3575 306174
rect 66897 305826 66963 305829
rect 66897 305824 68908 305826
rect 66897 305768 66902 305824
rect 66958 305768 68908 305824
rect 66897 305766 68908 305768
rect 66897 305763 66963 305766
rect 157241 305282 157307 305285
rect 154652 305280 157307 305282
rect 154652 305224 157246 305280
rect 157302 305224 157307 305280
rect 154652 305222 157307 305224
rect 157241 305219 157307 305222
rect 220169 305010 220235 305013
rect 222101 305010 222167 305013
rect 298093 305010 298159 305013
rect 220169 305008 298159 305010
rect 220169 304952 220174 305008
rect 220230 304952 222106 305008
rect 222162 304952 298098 305008
rect 298154 304952 298159 305008
rect 220169 304950 298159 304952
rect 220169 304947 220235 304950
rect 222101 304947 222167 304950
rect 298093 304947 298159 304950
rect 67173 304738 67239 304741
rect 67173 304736 68908 304738
rect 67173 304680 67178 304736
rect 67234 304680 68908 304736
rect 67173 304678 68908 304680
rect 67173 304675 67239 304678
rect 156045 304194 156111 304197
rect 154652 304192 156111 304194
rect 154652 304136 156050 304192
rect 156106 304136 156111 304192
rect 154652 304134 156111 304136
rect 156045 304131 156111 304134
rect 66897 303650 66963 303653
rect 156689 303650 156755 303653
rect 253933 303650 253999 303653
rect 66897 303648 68908 303650
rect 66897 303592 66902 303648
rect 66958 303592 68908 303648
rect 66897 303590 68908 303592
rect 156689 303648 253999 303650
rect 156689 303592 156694 303648
rect 156750 303592 253938 303648
rect 253994 303592 253999 303648
rect 156689 303590 253999 303592
rect 66897 303587 66963 303590
rect 156689 303587 156755 303590
rect 253933 303587 253999 303590
rect 157241 303106 157307 303109
rect 154652 303104 157307 303106
rect 154652 303048 157246 303104
rect 157302 303048 157307 303104
rect 154652 303046 157307 303048
rect 157241 303043 157307 303046
rect 66989 302562 67055 302565
rect 66989 302560 68908 302562
rect 66989 302504 66994 302560
rect 67050 302504 68908 302560
rect 66989 302502 68908 302504
rect 66989 302499 67055 302502
rect 235165 302426 235231 302429
rect 299565 302426 299631 302429
rect 235165 302424 299631 302426
rect 235165 302368 235170 302424
rect 235226 302368 299570 302424
rect 299626 302368 299631 302424
rect 235165 302366 299631 302368
rect 235165 302363 235231 302366
rect 299565 302363 299631 302366
rect 192569 302290 192635 302293
rect 193121 302290 193187 302293
rect 262857 302290 262923 302293
rect 192569 302288 262923 302290
rect 192569 302232 192574 302288
rect 192630 302232 193126 302288
rect 193182 302232 262862 302288
rect 262918 302232 262923 302288
rect 192569 302230 262923 302232
rect 192569 302227 192635 302230
rect 193121 302227 193187 302230
rect 262857 302227 262923 302230
rect 156781 302018 156847 302021
rect 154652 302016 156847 302018
rect 154652 301960 156786 302016
rect 156842 301960 156847 302016
rect 154652 301958 156847 301960
rect 156781 301955 156847 301958
rect 65977 301474 66043 301477
rect 65977 301472 68908 301474
rect 65977 301416 65982 301472
rect 66038 301416 68908 301472
rect 65977 301414 68908 301416
rect 65977 301411 66043 301414
rect 200113 301338 200179 301341
rect 200757 301338 200823 301341
rect 200113 301336 209790 301338
rect 200113 301280 200118 301336
rect 200174 301280 200762 301336
rect 200818 301280 209790 301336
rect 200113 301278 209790 301280
rect 200113 301275 200179 301278
rect 200757 301275 200823 301278
rect 154622 300930 154682 301172
rect 209730 301066 209790 301278
rect 260097 301066 260163 301069
rect 209730 301064 260163 301066
rect 209730 301008 260102 301064
rect 260158 301008 260163 301064
rect 209730 301006 260163 301008
rect 260097 301003 260163 301006
rect 304257 300930 304323 300933
rect 154622 300928 304323 300930
rect 154622 300872 304262 300928
rect 304318 300872 304323 300928
rect 154622 300870 304323 300872
rect 304257 300867 304323 300870
rect 240869 300794 240935 300797
rect 241513 300794 241579 300797
rect 240869 300792 241579 300794
rect 240869 300736 240874 300792
rect 240930 300736 241518 300792
rect 241574 300736 241579 300792
rect 240869 300734 241579 300736
rect 240869 300731 240935 300734
rect 241513 300731 241579 300734
rect 66897 300658 66963 300661
rect 66897 300656 68908 300658
rect 66897 300600 66902 300656
rect 66958 300600 68908 300656
rect 66897 300598 68908 300600
rect 66897 300595 66963 300598
rect 163497 300250 163563 300253
rect 245837 300250 245903 300253
rect 163497 300248 245903 300250
rect 163497 300192 163502 300248
rect 163558 300192 245842 300248
rect 245898 300192 245903 300248
rect 163497 300190 245903 300192
rect 163497 300187 163563 300190
rect 245837 300187 245903 300190
rect 157149 300114 157215 300117
rect 154652 300112 157215 300114
rect 154652 300056 157154 300112
rect 157210 300056 157215 300112
rect 154652 300054 157215 300056
rect 157149 300051 157215 300054
rect 240869 300114 240935 300117
rect 583201 300114 583267 300117
rect 240869 300112 583267 300114
rect 240869 300056 240874 300112
rect 240930 300056 583206 300112
rect 583262 300056 583267 300112
rect 240869 300054 583267 300056
rect 240869 300051 240935 300054
rect 583201 300051 583267 300054
rect 67081 299570 67147 299573
rect 67081 299568 68908 299570
rect 67081 299512 67086 299568
rect 67142 299512 68908 299568
rect 67081 299510 68908 299512
rect 67081 299507 67147 299510
rect 157241 299026 157307 299029
rect 154652 299024 157307 299026
rect 154652 298968 157246 299024
rect 157302 298968 157307 299024
rect 154652 298966 157307 298968
rect 157241 298963 157307 298966
rect 580257 298754 580323 298757
rect 583520 298754 584960 298844
rect 580257 298752 584960 298754
rect 580257 298696 580262 298752
rect 580318 298696 584960 298752
rect 580257 298694 584960 298696
rect 580257 298691 580323 298694
rect 583520 298604 584960 298694
rect 67357 298482 67423 298485
rect 67357 298480 68908 298482
rect 67357 298424 67362 298480
rect 67418 298424 68908 298480
rect 67357 298422 68908 298424
rect 67357 298419 67423 298422
rect 209129 298346 209195 298349
rect 209405 298346 209471 298349
rect 269757 298346 269823 298349
rect 209129 298344 269823 298346
rect 209129 298288 209134 298344
rect 209190 298288 209410 298344
rect 209466 298288 269762 298344
rect 269818 298288 269823 298344
rect 209129 298286 269823 298288
rect 209129 298283 209195 298286
rect 209405 298283 209471 298286
rect 269757 298283 269823 298286
rect 173249 298210 173315 298213
rect 256877 298210 256943 298213
rect 173249 298208 256943 298210
rect 173249 298152 173254 298208
rect 173310 298152 256882 298208
rect 256938 298152 256943 298208
rect 173249 298150 256943 298152
rect 173249 298147 173315 298150
rect 256877 298147 256943 298150
rect 215293 298074 215359 298077
rect 215937 298074 216003 298077
rect 215293 298072 216003 298074
rect 215293 298016 215298 298072
rect 215354 298016 215942 298072
rect 215998 298016 216003 298072
rect 215293 298014 216003 298016
rect 215293 298011 215359 298014
rect 215937 298011 216003 298014
rect 156413 297938 156479 297941
rect 154652 297936 156479 297938
rect 154652 297880 156418 297936
rect 156474 297880 156479 297936
rect 154652 297878 156479 297880
rect 156413 297875 156479 297878
rect 67766 297332 67772 297396
rect 67836 297394 67842 297396
rect 185669 297394 185735 297397
rect 241646 297394 241652 297396
rect 67836 297334 68908 297394
rect 185669 297392 241652 297394
rect 185669 297336 185674 297392
rect 185730 297336 241652 297392
rect 185669 297334 241652 297336
rect 67836 297332 67842 297334
rect 185669 297331 185735 297334
rect 241646 297332 241652 297334
rect 241716 297332 241722 297396
rect 215293 296986 215359 296989
rect 251265 296986 251331 296989
rect 215293 296984 251331 296986
rect 215293 296928 215298 296984
rect 215354 296928 251270 296984
rect 251326 296928 251331 296984
rect 215293 296926 251331 296928
rect 215293 296923 215359 296926
rect 251265 296923 251331 296926
rect 156689 296850 156755 296853
rect 154652 296848 156755 296850
rect 154652 296792 156694 296848
rect 156750 296792 156755 296848
rect 154652 296790 156755 296792
rect 156689 296787 156755 296790
rect 218697 296850 218763 296853
rect 221038 296850 221044 296852
rect 218697 296848 221044 296850
rect 218697 296792 218702 296848
rect 218758 296792 221044 296848
rect 218697 296790 221044 296792
rect 218697 296787 218763 296790
rect 221038 296788 221044 296790
rect 221108 296788 221114 296852
rect 233693 296850 233759 296853
rect 583661 296850 583727 296853
rect 233693 296848 583727 296850
rect 233693 296792 233698 296848
rect 233754 296792 583666 296848
rect 583722 296792 583727 296848
rect 233693 296790 583727 296792
rect 233693 296787 233759 296790
rect 583661 296787 583727 296790
rect 66897 296306 66963 296309
rect 66897 296304 68908 296306
rect 66897 296248 66902 296304
rect 66958 296248 68908 296304
rect 66897 296246 68908 296248
rect 66897 296243 66963 296246
rect 180006 295972 180012 296036
rect 180076 296034 180082 296036
rect 201493 296034 201559 296037
rect 210417 296034 210483 296037
rect 180076 296032 210483 296034
rect 180076 295976 201498 296032
rect 201554 295976 210422 296032
rect 210478 295976 210483 296032
rect 180076 295974 210483 295976
rect 180076 295972 180082 295974
rect 201493 295971 201559 295974
rect 210417 295971 210483 295974
rect 154622 295354 154682 295732
rect 162117 295490 162183 295493
rect 225413 295490 225479 295493
rect 162117 295488 225479 295490
rect 162117 295432 162122 295488
rect 162178 295432 225418 295488
rect 225474 295432 225479 295488
rect 162117 295430 225479 295432
rect 162117 295427 162183 295430
rect 225413 295427 225479 295430
rect 225597 295490 225663 295493
rect 229737 295490 229803 295493
rect 225597 295488 229803 295490
rect 225597 295432 225602 295488
rect 225658 295432 229742 295488
rect 229798 295432 229803 295488
rect 225597 295430 229803 295432
rect 225597 295427 225663 295430
rect 229737 295427 229803 295430
rect 158621 295356 158687 295357
rect 158621 295354 158668 295356
rect 154622 295352 158668 295354
rect 158732 295354 158738 295356
rect 206277 295354 206343 295357
rect 206645 295354 206711 295357
rect 582925 295354 582991 295357
rect 154622 295296 158626 295352
rect 154622 295294 158668 295296
rect 158621 295292 158668 295294
rect 158732 295294 158778 295354
rect 206277 295352 582991 295354
rect 206277 295296 206282 295352
rect 206338 295296 206650 295352
rect 206706 295296 582930 295352
rect 582986 295296 582991 295352
rect 206277 295294 582991 295296
rect 158732 295292 158738 295294
rect 158621 295291 158687 295292
rect 206277 295291 206343 295294
rect 206645 295291 206711 295294
rect 582925 295291 582991 295294
rect 68878 295082 68938 295188
rect 69054 295082 69060 295084
rect 68878 295022 69060 295082
rect 68878 294538 68938 295022
rect 69054 295020 69060 295022
rect 69124 295020 69130 295084
rect 156321 294674 156387 294677
rect 154652 294672 156387 294674
rect 154652 294616 156326 294672
rect 156382 294616 156387 294672
rect 154652 294614 156387 294616
rect 156321 294611 156387 294614
rect 64830 294478 68938 294538
rect 199377 294538 199443 294541
rect 225965 294538 226031 294541
rect 199377 294536 226031 294538
rect 199377 294480 199382 294536
rect 199438 294480 225970 294536
rect 226026 294480 226031 294536
rect 199377 294478 226031 294480
rect 25497 293994 25563 293997
rect 64830 293994 64890 294478
rect 199377 294475 199443 294478
rect 225965 294475 226031 294478
rect 67081 294130 67147 294133
rect 185669 294130 185735 294133
rect 241421 294130 241487 294133
rect 67081 294128 68908 294130
rect 67081 294072 67086 294128
rect 67142 294072 68908 294128
rect 67081 294070 68908 294072
rect 185669 294128 241487 294130
rect 185669 294072 185674 294128
rect 185730 294072 241426 294128
rect 241482 294072 241487 294128
rect 185669 294070 241487 294072
rect 67081 294067 67147 294070
rect 185669 294067 185735 294070
rect 241421 294067 241487 294070
rect 25497 293992 64890 293994
rect 25497 293936 25502 293992
rect 25558 293936 64890 293992
rect 25497 293934 64890 293936
rect 238017 293994 238083 293997
rect 239029 293994 239095 293997
rect 583753 293994 583819 293997
rect 238017 293992 583819 293994
rect 238017 293936 238022 293992
rect 238078 293936 239034 293992
rect 239090 293936 583758 293992
rect 583814 293936 583819 293992
rect 238017 293934 583819 293936
rect 25497 293931 25563 293934
rect 238017 293931 238083 293934
rect 239029 293931 239095 293934
rect 583753 293931 583819 293934
rect -960 293178 480 293268
rect 2773 293178 2839 293181
rect -960 293176 2839 293178
rect -960 293120 2778 293176
rect 2834 293120 2839 293176
rect -960 293118 2839 293120
rect -960 293028 480 293118
rect 2773 293115 2839 293118
rect 66713 293042 66779 293045
rect 154622 293042 154682 293556
rect 66713 293040 68908 293042
rect 66713 292984 66718 293040
rect 66774 292984 68908 293040
rect 66713 292982 68908 292984
rect 154622 292982 157442 293042
rect 66713 292979 66779 292982
rect 157241 292770 157307 292773
rect 154652 292768 157307 292770
rect 154652 292712 157246 292768
rect 157302 292712 157307 292768
rect 154652 292710 157307 292712
rect 157241 292707 157307 292710
rect 157382 292634 157442 292982
rect 198089 292906 198155 292909
rect 254025 292906 254091 292909
rect 198089 292904 254091 292906
rect 198089 292848 198094 292904
rect 198150 292848 254030 292904
rect 254086 292848 254091 292904
rect 198089 292846 254091 292848
rect 198089 292843 198155 292846
rect 254025 292843 254091 292846
rect 157517 292770 157583 292773
rect 247217 292770 247283 292773
rect 157517 292768 247283 292770
rect 157517 292712 157522 292768
rect 157578 292712 247222 292768
rect 247278 292712 247283 292768
rect 157517 292710 247283 292712
rect 157517 292707 157583 292710
rect 247217 292707 247283 292710
rect 166206 292634 166212 292636
rect 157382 292574 166212 292634
rect 166206 292572 166212 292574
rect 166276 292572 166282 292636
rect 225321 292634 225387 292637
rect 228357 292634 228423 292637
rect 225321 292632 228423 292634
rect 225321 292576 225326 292632
rect 225382 292576 228362 292632
rect 228418 292576 228423 292632
rect 225321 292574 228423 292576
rect 225321 292571 225387 292574
rect 228357 292571 228423 292574
rect 233877 292634 233943 292637
rect 583109 292634 583175 292637
rect 233877 292632 583175 292634
rect 233877 292576 233882 292632
rect 233938 292576 583114 292632
rect 583170 292576 583175 292632
rect 233877 292574 583175 292576
rect 233877 292571 233943 292574
rect 583109 292571 583175 292574
rect 66897 292226 66963 292229
rect 66897 292224 68908 292226
rect 66897 292168 66902 292224
rect 66958 292168 68908 292224
rect 66897 292166 68908 292168
rect 66897 292163 66963 292166
rect 213177 291818 213243 291821
rect 582465 291818 582531 291821
rect 213177 291816 582531 291818
rect 213177 291760 213182 291816
rect 213238 291760 582470 291816
rect 582526 291760 582531 291816
rect 213177 291758 582531 291760
rect 213177 291755 213243 291758
rect 582465 291755 582531 291758
rect 156781 291682 156847 291685
rect 154652 291680 156847 291682
rect 154652 291624 156786 291680
rect 156842 291624 156847 291680
rect 154652 291622 156847 291624
rect 156781 291619 156847 291622
rect 195421 291546 195487 291549
rect 201401 291546 201467 291549
rect 195421 291544 201467 291546
rect 195421 291488 195426 291544
rect 195482 291488 201406 291544
rect 201462 291488 201467 291544
rect 195421 291486 201467 291488
rect 195421 291483 195487 291486
rect 201401 291483 201467 291486
rect 170397 291410 170463 291413
rect 197353 291410 197419 291413
rect 170397 291408 197419 291410
rect 170397 291352 170402 291408
rect 170458 291352 197358 291408
rect 197414 291352 197419 291408
rect 170397 291350 197419 291352
rect 170397 291347 170463 291350
rect 197353 291347 197419 291350
rect 199326 291348 199332 291412
rect 199396 291410 199402 291412
rect 232773 291410 232839 291413
rect 199396 291408 232839 291410
rect 199396 291352 232778 291408
rect 232834 291352 232839 291408
rect 199396 291350 232839 291352
rect 199396 291348 199402 291350
rect 232773 291347 232839 291350
rect 183001 291274 183067 291277
rect 217869 291274 217935 291277
rect 183001 291272 217935 291274
rect 183001 291216 183006 291272
rect 183062 291216 217874 291272
rect 217930 291216 217935 291272
rect 183001 291214 217935 291216
rect 183001 291211 183067 291214
rect 217869 291211 217935 291214
rect 218053 291274 218119 291277
rect 254117 291274 254183 291277
rect 218053 291272 254183 291274
rect 218053 291216 218058 291272
rect 218114 291216 254122 291272
rect 254178 291216 254183 291272
rect 218053 291214 254183 291216
rect 218053 291211 218119 291214
rect 254117 291211 254183 291214
rect 66989 291138 67055 291141
rect 66989 291136 68908 291138
rect 66989 291080 66994 291136
rect 67050 291080 68908 291136
rect 66989 291078 68908 291080
rect 66989 291075 67055 291078
rect 156454 291076 156460 291140
rect 156524 291138 156530 291140
rect 156689 291138 156755 291141
rect 156524 291136 156755 291138
rect 156524 291080 156694 291136
rect 156750 291080 156755 291136
rect 156524 291078 156755 291080
rect 156524 291076 156530 291078
rect 156689 291075 156755 291078
rect 159449 291138 159515 291141
rect 233693 291138 233759 291141
rect 159449 291136 233759 291138
rect 159449 291080 159454 291136
rect 159510 291080 233698 291136
rect 233754 291080 233759 291136
rect 159449 291078 233759 291080
rect 159449 291075 159515 291078
rect 233693 291075 233759 291078
rect 157241 290594 157307 290597
rect 154652 290592 157307 290594
rect 154652 290536 157246 290592
rect 157302 290536 157307 290592
rect 154652 290534 157307 290536
rect 157241 290531 157307 290534
rect 156689 290186 156755 290189
rect 247125 290186 247191 290189
rect 156689 290184 247191 290186
rect 156689 290128 156694 290184
rect 156750 290128 247130 290184
rect 247186 290128 247191 290184
rect 156689 290126 247191 290128
rect 156689 290123 156755 290126
rect 247125 290123 247191 290126
rect 66897 290050 66963 290053
rect 239489 290050 239555 290053
rect 280286 290050 280292 290052
rect 66897 290048 68908 290050
rect 66897 289992 66902 290048
rect 66958 289992 68908 290048
rect 66897 289990 68908 289992
rect 239489 290048 280292 290050
rect 239489 289992 239494 290048
rect 239550 289992 280292 290048
rect 239489 289990 280292 289992
rect 66897 289987 66963 289990
rect 239489 289987 239555 289990
rect 280286 289988 280292 289990
rect 280356 289988 280362 290052
rect 210417 289778 210483 289781
rect 583017 289778 583083 289781
rect 210417 289776 583083 289778
rect 210417 289720 210422 289776
rect 210478 289720 583022 289776
rect 583078 289720 583083 289776
rect 210417 289718 583083 289720
rect 210417 289715 210483 289718
rect 583017 289715 583083 289718
rect 222469 289642 222535 289645
rect 223021 289642 223087 289645
rect 222469 289640 223087 289642
rect 222469 289584 222474 289640
rect 222530 289584 223026 289640
rect 223082 289584 223087 289640
rect 222469 289582 223087 289584
rect 222469 289579 222535 289582
rect 223021 289579 223087 289582
rect 156781 289506 156847 289509
rect 154652 289504 156847 289506
rect 154652 289448 156786 289504
rect 156842 289448 156847 289504
rect 154652 289446 156847 289448
rect 156781 289443 156847 289446
rect 160921 289098 160987 289101
rect 160921 289096 180810 289098
rect 160921 289040 160926 289096
rect 160982 289040 180810 289096
rect 160921 289038 180810 289040
rect 160921 289035 160987 289038
rect 66897 288962 66963 288965
rect 66897 288960 68908 288962
rect 66897 288904 66902 288960
rect 66958 288904 68908 288960
rect 66897 288902 68908 288904
rect 66897 288899 66963 288902
rect 180750 288826 180810 289038
rect 191649 288826 191715 288829
rect 203149 288826 203215 288829
rect 180750 288824 203215 288826
rect 180750 288768 191654 288824
rect 191710 288768 203154 288824
rect 203210 288768 203215 288824
rect 180750 288766 203215 288768
rect 191649 288763 191715 288766
rect 203149 288763 203215 288766
rect 200614 288628 200620 288692
rect 200684 288690 200690 288692
rect 216765 288690 216831 288693
rect 200684 288688 216831 288690
rect 200684 288632 216770 288688
rect 216826 288632 216831 288688
rect 200684 288630 216831 288632
rect 200684 288628 200690 288630
rect 216765 288627 216831 288630
rect 222469 288690 222535 288693
rect 233182 288690 233188 288692
rect 222469 288688 233188 288690
rect 222469 288632 222474 288688
rect 222530 288632 233188 288688
rect 222469 288630 233188 288632
rect 222469 288627 222535 288630
rect 233182 288628 233188 288630
rect 233252 288628 233258 288692
rect 202229 288554 202295 288557
rect 288566 288554 288572 288556
rect 202229 288552 288572 288554
rect 202229 288496 202234 288552
rect 202290 288496 288572 288552
rect 202229 288494 288572 288496
rect 202229 288491 202295 288494
rect 288566 288492 288572 288494
rect 288636 288492 288642 288556
rect 156229 288418 156295 288421
rect 154652 288416 156295 288418
rect 154652 288360 156234 288416
rect 156290 288360 156295 288416
rect 154652 288358 156295 288360
rect 156229 288355 156295 288358
rect 66713 287874 66779 287877
rect 66713 287872 68908 287874
rect 66713 287816 66718 287872
rect 66774 287816 68908 287872
rect 66713 287814 68908 287816
rect 66713 287811 66779 287814
rect 197997 287466 198063 287469
rect 206093 287466 206159 287469
rect 197997 287464 206159 287466
rect 197997 287408 198002 287464
rect 198058 287408 206098 287464
rect 206154 287408 206159 287464
rect 197997 287406 206159 287408
rect 197997 287403 198063 287406
rect 206093 287403 206159 287406
rect 229737 287466 229803 287469
rect 249793 287466 249859 287469
rect 229737 287464 249859 287466
rect 229737 287408 229742 287464
rect 229798 287408 249798 287464
rect 249854 287408 249859 287464
rect 229737 287406 249859 287408
rect 229737 287403 229803 287406
rect 249793 287403 249859 287406
rect 156689 287330 156755 287333
rect 154652 287328 156755 287330
rect 154652 287272 156694 287328
rect 156750 287272 156755 287328
rect 154652 287270 156755 287272
rect 156689 287267 156755 287270
rect 198733 287330 198799 287333
rect 223021 287330 223087 287333
rect 198733 287328 223087 287330
rect 198733 287272 198738 287328
rect 198794 287272 223026 287328
rect 223082 287272 223087 287328
rect 198733 287270 223087 287272
rect 198733 287267 198799 287270
rect 223021 287267 223087 287270
rect 239949 287330 240015 287333
rect 287278 287330 287284 287332
rect 239949 287328 287284 287330
rect 239949 287272 239954 287328
rect 240010 287272 287284 287328
rect 239949 287270 287284 287272
rect 239949 287267 240015 287270
rect 287278 287268 287284 287270
rect 287348 287268 287354 287332
rect 199469 287194 199535 287197
rect 203701 287194 203767 287197
rect 199469 287192 203767 287194
rect 199469 287136 199474 287192
rect 199530 287136 203706 287192
rect 203762 287136 203767 287192
rect 199469 287134 203767 287136
rect 199469 287131 199535 287134
rect 203701 287131 203767 287134
rect 209037 287194 209103 287197
rect 211654 287194 211660 287196
rect 209037 287192 211660 287194
rect 209037 287136 209042 287192
rect 209098 287136 211660 287192
rect 209037 287134 211660 287136
rect 209037 287131 209103 287134
rect 211654 287132 211660 287134
rect 211724 287132 211730 287196
rect 211981 287194 212047 287197
rect 284293 287194 284359 287197
rect 211981 287192 284359 287194
rect 211981 287136 211986 287192
rect 212042 287136 284298 287192
rect 284354 287136 284359 287192
rect 211981 287134 284359 287136
rect 211981 287131 212047 287134
rect 284293 287131 284359 287134
rect 66897 286786 66963 286789
rect 66897 286784 68908 286786
rect 66897 286728 66902 286784
rect 66958 286728 68908 286784
rect 66897 286726 68908 286728
rect 66897 286723 66963 286726
rect 169017 286378 169083 286381
rect 213177 286378 213243 286381
rect 169017 286376 213243 286378
rect 169017 286320 169022 286376
rect 169078 286320 213182 286376
rect 213238 286320 213243 286376
rect 169017 286318 213243 286320
rect 169017 286315 169083 286318
rect 213177 286315 213243 286318
rect 157241 286242 157307 286245
rect 154652 286240 157307 286242
rect 154652 286184 157246 286240
rect 157302 286184 157307 286240
rect 154652 286182 157307 286184
rect 157241 286179 157307 286182
rect 226517 286106 226583 286109
rect 269849 286106 269915 286109
rect 226517 286104 269915 286106
rect 226517 286048 226522 286104
rect 226578 286048 269854 286104
rect 269910 286048 269915 286104
rect 226517 286046 269915 286048
rect 226517 286043 226583 286046
rect 269849 286043 269915 286046
rect 184473 285970 184539 285973
rect 210877 285970 210943 285973
rect 184473 285968 210943 285970
rect 184473 285912 184478 285968
rect 184534 285912 210882 285968
rect 210938 285912 210943 285968
rect 184473 285910 210943 285912
rect 184473 285907 184539 285910
rect 210877 285907 210943 285910
rect 219157 285970 219223 285973
rect 226926 285970 226932 285972
rect 219157 285968 226932 285970
rect 219157 285912 219162 285968
rect 219218 285912 226932 285968
rect 219157 285910 226932 285912
rect 219157 285907 219223 285910
rect 226926 285908 226932 285910
rect 226996 285908 227002 285972
rect 230565 285970 230631 285973
rect 240358 285970 240364 285972
rect 230565 285968 240364 285970
rect 230565 285912 230570 285968
rect 230626 285912 240364 285968
rect 230565 285910 240364 285912
rect 230565 285907 230631 285910
rect 240358 285908 240364 285910
rect 240428 285908 240434 285972
rect 225045 285834 225111 285837
rect 238518 285834 238524 285836
rect 225045 285832 238524 285834
rect 225045 285776 225050 285832
rect 225106 285776 238524 285832
rect 225045 285774 238524 285776
rect 225045 285771 225111 285774
rect 238518 285772 238524 285774
rect 238588 285772 238594 285836
rect 242249 285834 242315 285837
rect 243445 285834 243511 285837
rect 242249 285832 243511 285834
rect 242249 285776 242254 285832
rect 242310 285776 243450 285832
rect 243506 285776 243511 285832
rect 242249 285774 243511 285776
rect 242249 285771 242315 285774
rect 243445 285771 243511 285774
rect 66805 285698 66871 285701
rect 199561 285698 199627 285701
rect 202229 285698 202295 285701
rect 66805 285696 68908 285698
rect 66805 285640 66810 285696
rect 66866 285640 68908 285696
rect 66805 285638 68908 285640
rect 199561 285696 202295 285698
rect 199561 285640 199566 285696
rect 199622 285640 202234 285696
rect 202290 285640 202295 285696
rect 199561 285638 202295 285640
rect 66805 285635 66871 285638
rect 199561 285635 199627 285638
rect 202229 285635 202295 285638
rect 220077 285698 220143 285701
rect 224902 285698 224908 285700
rect 220077 285696 224908 285698
rect 220077 285640 220082 285696
rect 220138 285640 224908 285696
rect 220077 285638 224908 285640
rect 220077 285635 220143 285638
rect 224902 285636 224908 285638
rect 224972 285636 224978 285700
rect 235993 285698 236059 285701
rect 236494 285698 236500 285700
rect 235993 285696 236500 285698
rect 235993 285640 235998 285696
rect 236054 285640 236500 285696
rect 235993 285638 236500 285640
rect 235993 285635 236059 285638
rect 236494 285636 236500 285638
rect 236564 285636 236570 285700
rect 583520 285276 584960 285516
rect 156321 285154 156387 285157
rect 154652 285152 156387 285154
rect 154652 285096 156326 285152
rect 156382 285096 156387 285152
rect 154652 285094 156387 285096
rect 156321 285091 156387 285094
rect 66989 284610 67055 284613
rect 200021 284610 200087 284613
rect 211981 284610 212047 284613
rect 66989 284608 68908 284610
rect 66989 284552 66994 284608
rect 67050 284552 68908 284608
rect 66989 284550 68908 284552
rect 200021 284608 212047 284610
rect 200021 284552 200026 284608
rect 200082 284552 211986 284608
rect 212042 284552 212047 284608
rect 200021 284550 212047 284552
rect 66989 284547 67055 284550
rect 200021 284547 200087 284550
rect 211981 284547 212047 284550
rect 199653 284474 199719 284477
rect 217317 284474 217383 284477
rect 199653 284472 217383 284474
rect 199653 284416 199658 284472
rect 199714 284416 217322 284472
rect 217378 284416 217383 284472
rect 199653 284414 217383 284416
rect 199653 284411 199719 284414
rect 217317 284411 217383 284414
rect 230473 284474 230539 284477
rect 231669 284474 231735 284477
rect 281574 284474 281580 284476
rect 230473 284472 281580 284474
rect 230473 284416 230478 284472
rect 230534 284416 231674 284472
rect 231730 284416 281580 284472
rect 230473 284414 281580 284416
rect 230473 284411 230539 284414
rect 231669 284411 231735 284414
rect 281574 284412 281580 284414
rect 281644 284412 281650 284476
rect 157241 284338 157307 284341
rect 154652 284336 157307 284338
rect 154652 284280 157246 284336
rect 157302 284280 157307 284336
rect 154652 284278 157307 284280
rect 157241 284275 157307 284278
rect 167637 284338 167703 284341
rect 204253 284338 204319 284341
rect 167637 284336 204319 284338
rect 167637 284280 167642 284336
rect 167698 284280 204258 284336
rect 204314 284280 204319 284336
rect 167637 284278 204319 284280
rect 167637 284275 167703 284278
rect 204253 284275 204319 284278
rect 212349 284338 212415 284341
rect 582465 284338 582531 284341
rect 212349 284336 582531 284338
rect 212349 284280 212354 284336
rect 212410 284280 582470 284336
rect 582526 284280 582531 284336
rect 212349 284278 582531 284280
rect 212349 284275 212415 284278
rect 582465 284275 582531 284278
rect 243629 284066 243695 284069
rect 244089 284066 244155 284069
rect 243629 284064 244155 284066
rect 243629 284008 243634 284064
rect 243690 284008 244094 284064
rect 244150 284008 244155 284064
rect 243629 284006 244155 284008
rect 243629 284003 243695 284006
rect 244089 284003 244155 284006
rect 205357 283932 205423 283933
rect 205357 283930 205404 283932
rect 205312 283928 205404 283930
rect 205312 283872 205362 283928
rect 205312 283870 205404 283872
rect 205357 283868 205404 283870
rect 205468 283868 205474 283932
rect 206870 283868 206876 283932
rect 206940 283930 206946 283932
rect 207105 283930 207171 283933
rect 206940 283928 207171 283930
rect 206940 283872 207110 283928
rect 207166 283872 207171 283928
rect 206940 283870 207171 283872
rect 206940 283868 206946 283870
rect 205357 283867 205423 283868
rect 207105 283867 207171 283870
rect 208669 283930 208735 283933
rect 214097 283932 214163 283933
rect 209630 283930 209636 283932
rect 208669 283928 209636 283930
rect 208669 283872 208674 283928
rect 208730 283872 209636 283928
rect 208669 283870 209636 283872
rect 208669 283867 208735 283870
rect 209630 283868 209636 283870
rect 209700 283868 209706 283932
rect 214046 283930 214052 283932
rect 214006 283870 214052 283930
rect 214116 283928 214163 283932
rect 214158 283872 214163 283928
rect 214046 283868 214052 283870
rect 214116 283868 214163 283872
rect 215334 283868 215340 283932
rect 215404 283930 215410 283932
rect 215937 283930 216003 283933
rect 215404 283928 216003 283930
rect 215404 283872 215942 283928
rect 215998 283872 216003 283928
rect 215404 283870 216003 283872
rect 215404 283868 215410 283870
rect 214097 283867 214163 283868
rect 215937 283867 216003 283870
rect 217174 283868 217180 283932
rect 217244 283930 217250 283932
rect 217409 283930 217475 283933
rect 224677 283932 224743 283933
rect 224677 283930 224724 283932
rect 217244 283928 217475 283930
rect 217244 283872 217414 283928
rect 217470 283872 217475 283928
rect 217244 283870 217475 283872
rect 224632 283928 224724 283930
rect 224632 283872 224682 283928
rect 224632 283870 224724 283872
rect 217244 283868 217250 283870
rect 217409 283867 217475 283870
rect 224677 283868 224724 283870
rect 224788 283868 224794 283932
rect 226374 283868 226380 283932
rect 226444 283930 226450 283932
rect 226609 283930 226675 283933
rect 226444 283928 226675 283930
rect 226444 283872 226614 283928
rect 226670 283872 226675 283928
rect 226444 283870 226675 283872
rect 226444 283868 226450 283870
rect 224677 283867 224743 283868
rect 226609 283867 226675 283870
rect 227989 283930 228055 283933
rect 228766 283930 228772 283932
rect 227989 283928 228772 283930
rect 227989 283872 227994 283928
rect 228050 283872 228772 283928
rect 227989 283870 228772 283872
rect 227989 283867 228055 283870
rect 228766 283868 228772 283870
rect 228836 283868 228842 283932
rect 229461 283930 229527 283933
rect 229686 283930 229692 283932
rect 229461 283928 229692 283930
rect 229461 283872 229466 283928
rect 229522 283872 229692 283928
rect 229461 283870 229692 283872
rect 229461 283867 229527 283870
rect 229686 283868 229692 283870
rect 229756 283868 229762 283932
rect 231577 283930 231643 283933
rect 231710 283930 231716 283932
rect 231577 283928 231716 283930
rect 231577 283872 231582 283928
rect 231638 283872 231716 283928
rect 231577 283870 231716 283872
rect 231577 283867 231643 283870
rect 231710 283868 231716 283870
rect 231780 283868 231786 283932
rect 236494 283868 236500 283932
rect 236564 283930 236570 283932
rect 236729 283930 236795 283933
rect 236564 283928 236795 283930
rect 236564 283872 236734 283928
rect 236790 283872 236795 283928
rect 236564 283870 236795 283872
rect 236564 283868 236570 283870
rect 236729 283867 236795 283870
rect 66713 283794 66779 283797
rect 197353 283794 197419 283797
rect 248597 283794 248663 283797
rect 66713 283792 68908 283794
rect 66713 283736 66718 283792
rect 66774 283736 68908 283792
rect 66713 283734 68908 283736
rect 197353 283792 200284 283794
rect 197353 283736 197358 283792
rect 197414 283736 200284 283792
rect 197353 283734 200284 283736
rect 244076 283792 248663 283794
rect 244076 283736 248602 283792
rect 248658 283736 248663 283792
rect 244076 283734 248663 283736
rect 66713 283731 66779 283734
rect 197353 283731 197419 283734
rect 248597 283731 248663 283734
rect 189809 283522 189875 283525
rect 198733 283522 198799 283525
rect 189809 283520 198799 283522
rect 189809 283464 189814 283520
rect 189870 283464 198738 283520
rect 198794 283464 198799 283520
rect 189809 283462 198799 283464
rect 189809 283459 189875 283462
rect 198733 283459 198799 283462
rect 157241 283250 157307 283253
rect 246389 283250 246455 283253
rect 154652 283248 157307 283250
rect 154652 283192 157246 283248
rect 157302 283192 157307 283248
rect 154652 283190 157307 283192
rect 244076 283248 246455 283250
rect 244076 283192 246394 283248
rect 246450 283192 246455 283248
rect 244076 283190 246455 283192
rect 157241 283187 157307 283190
rect 246389 283187 246455 283190
rect 198549 282978 198615 282981
rect 244089 282978 244155 282981
rect 314653 282978 314719 282981
rect 198549 282976 200284 282978
rect 198549 282920 198554 282976
rect 198610 282920 200284 282976
rect 198549 282918 200284 282920
rect 244089 282976 314719 282978
rect 244089 282920 244094 282976
rect 244150 282920 314658 282976
rect 314714 282920 314719 282976
rect 244089 282918 314719 282920
rect 198549 282915 198615 282918
rect 244089 282915 244155 282918
rect 314653 282915 314719 282918
rect 66345 282706 66411 282709
rect 165153 282706 165219 282709
rect 200021 282706 200087 282709
rect 66345 282704 68908 282706
rect 66345 282648 66350 282704
rect 66406 282648 68908 282704
rect 66345 282646 68908 282648
rect 165153 282704 200087 282706
rect 165153 282648 165158 282704
rect 165214 282648 200026 282704
rect 200082 282648 200087 282704
rect 165153 282646 200087 282648
rect 66345 282643 66411 282646
rect 165153 282643 165219 282646
rect 200021 282643 200087 282646
rect 200062 282570 200068 282572
rect 180750 282510 200068 282570
rect 157149 282162 157215 282165
rect 154652 282160 157215 282162
rect 154652 282104 157154 282160
rect 157210 282104 157215 282160
rect 154652 282102 157215 282104
rect 157149 282099 157215 282102
rect 159541 282162 159607 282165
rect 180750 282162 180810 282510
rect 200062 282508 200068 282510
rect 200132 282508 200138 282572
rect 197353 282434 197419 282437
rect 245929 282434 245995 282437
rect 197353 282432 200284 282434
rect 197353 282376 197358 282432
rect 197414 282376 200284 282432
rect 197353 282374 200284 282376
rect 244076 282432 245995 282434
rect 244076 282376 245934 282432
rect 245990 282376 245995 282432
rect 244076 282374 245995 282376
rect 197353 282371 197419 282374
rect 245929 282371 245995 282374
rect 159541 282160 180810 282162
rect 159541 282104 159546 282160
rect 159602 282104 180810 282160
rect 159541 282102 180810 282104
rect 159541 282099 159607 282102
rect 67541 281618 67607 281621
rect 67541 281616 68908 281618
rect 67541 281560 67546 281616
rect 67602 281560 68908 281616
rect 67541 281558 68908 281560
rect 67541 281555 67607 281558
rect 197854 281556 197860 281620
rect 197924 281618 197930 281620
rect 246113 281618 246179 281621
rect 197924 281558 200284 281618
rect 244076 281616 246179 281618
rect 244076 281560 246118 281616
rect 246174 281560 246179 281616
rect 244076 281558 246179 281560
rect 197924 281556 197930 281558
rect 246113 281555 246179 281558
rect 157241 281074 157307 281077
rect 245929 281074 245995 281077
rect 154652 281072 157307 281074
rect 154652 281016 157246 281072
rect 157302 281016 157307 281072
rect 154652 281014 157307 281016
rect 244076 281072 245995 281074
rect 244076 281016 245934 281072
rect 245990 281016 245995 281072
rect 244076 281014 245995 281016
rect 157241 281011 157307 281014
rect 245929 281011 245995 281014
rect 197353 280802 197419 280805
rect 197353 280800 200284 280802
rect 197353 280744 197358 280800
rect 197414 280744 200284 280800
rect 197353 280742 200284 280744
rect 197353 280739 197419 280742
rect 66805 280530 66871 280533
rect 66805 280528 68908 280530
rect 66805 280472 66810 280528
rect 66866 280472 68908 280528
rect 66805 280470 68908 280472
rect 66805 280467 66871 280470
rect 197353 280258 197419 280261
rect 246113 280258 246179 280261
rect 197353 280256 200284 280258
rect -960 279972 480 280212
rect 197353 280200 197358 280256
rect 197414 280200 200284 280256
rect 197353 280198 200284 280200
rect 244076 280256 246179 280258
rect 244076 280200 246118 280256
rect 246174 280200 246179 280256
rect 244076 280198 246179 280200
rect 197353 280195 197419 280198
rect 246113 280195 246179 280198
rect 163446 280060 163452 280124
rect 163516 280122 163522 280124
rect 163589 280122 163655 280125
rect 195421 280122 195487 280125
rect 163516 280120 195487 280122
rect 163516 280064 163594 280120
rect 163650 280064 195426 280120
rect 195482 280064 195487 280120
rect 163516 280062 195487 280064
rect 163516 280060 163522 280062
rect 163589 280059 163655 280062
rect 195421 280059 195487 280062
rect 156965 279986 157031 279989
rect 154652 279984 157031 279986
rect 154652 279928 156970 279984
rect 157026 279928 157031 279984
rect 154652 279926 157031 279928
rect 156965 279923 157031 279926
rect 184565 279578 184631 279581
rect 199326 279578 199332 279580
rect 184565 279576 199332 279578
rect 184565 279520 184570 279576
rect 184626 279520 199332 279576
rect 184565 279518 199332 279520
rect 184565 279515 184631 279518
rect 199326 279516 199332 279518
rect 199396 279516 199402 279580
rect 67265 279442 67331 279445
rect 67950 279442 67956 279444
rect 67265 279440 67956 279442
rect 67265 279384 67270 279440
rect 67326 279384 67956 279440
rect 67265 279382 67956 279384
rect 67265 279379 67331 279382
rect 67950 279380 67956 279382
rect 68020 279442 68026 279444
rect 197445 279442 197511 279445
rect 245929 279442 245995 279445
rect 68020 279382 68908 279442
rect 197445 279440 200284 279442
rect 197445 279384 197450 279440
rect 197506 279384 200284 279440
rect 197445 279382 200284 279384
rect 244076 279440 245995 279442
rect 244076 279384 245934 279440
rect 245990 279384 245995 279440
rect 244076 279382 245995 279384
rect 68020 279380 68026 279382
rect 197445 279379 197511 279382
rect 245929 279379 245995 279382
rect 243486 279108 243492 279172
rect 243556 279108 243562 279172
rect 157241 278898 157307 278901
rect 154652 278896 157307 278898
rect 154652 278840 157246 278896
rect 157302 278840 157307 278896
rect 243494 278868 243554 279108
rect 154652 278838 157307 278840
rect 157241 278835 157307 278838
rect 197445 278626 197511 278629
rect 197445 278624 200284 278626
rect 197445 278568 197450 278624
rect 197506 278568 200284 278624
rect 197445 278566 200284 278568
rect 197445 278563 197511 278566
rect 66713 278354 66779 278357
rect 66713 278352 68908 278354
rect 66713 278296 66718 278352
rect 66774 278296 68908 278352
rect 66713 278294 68908 278296
rect 66713 278291 66779 278294
rect 198641 278082 198707 278085
rect 244273 278082 244339 278085
rect 198641 278080 200284 278082
rect 198641 278024 198646 278080
rect 198702 278024 200284 278080
rect 198641 278022 200284 278024
rect 244076 278080 244339 278082
rect 244076 278024 244278 278080
rect 244334 278024 244339 278080
rect 244076 278022 244339 278024
rect 198641 278019 198707 278022
rect 244273 278019 244339 278022
rect 193121 277946 193187 277949
rect 197353 277946 197419 277949
rect 193121 277944 197419 277946
rect 193121 277888 193126 277944
rect 193182 277888 197358 277944
rect 197414 277888 197419 277944
rect 193121 277886 197419 277888
rect 193121 277883 193187 277886
rect 197353 277883 197419 277886
rect 157241 277810 157307 277813
rect 154652 277808 157307 277810
rect 154652 277752 157246 277808
rect 157302 277752 157307 277808
rect 154652 277750 157307 277752
rect 157241 277747 157307 277750
rect 245929 277538 245995 277541
rect 244076 277536 245995 277538
rect 244076 277480 245934 277536
rect 245990 277480 245995 277536
rect 244076 277478 245995 277480
rect 245929 277475 245995 277478
rect 67081 277266 67147 277269
rect 197353 277266 197419 277269
rect 67081 277264 68908 277266
rect 67081 277208 67086 277264
rect 67142 277208 68908 277264
rect 67081 277206 68908 277208
rect 197353 277264 200284 277266
rect 197353 277208 197358 277264
rect 197414 277208 200284 277264
rect 197353 277206 200284 277208
rect 67081 277203 67147 277206
rect 197353 277203 197419 277206
rect 154665 276994 154731 276997
rect 154622 276992 154731 276994
rect 154622 276936 154670 276992
rect 154726 276936 154731 276992
rect 154622 276931 154731 276936
rect 154622 276722 154682 276931
rect 156873 276722 156939 276725
rect 154622 276720 156939 276722
rect 154622 276692 156878 276720
rect 154652 276664 156878 276692
rect 156934 276664 156939 276720
rect 154652 276662 156939 276664
rect 156873 276659 156939 276662
rect 197353 276722 197419 276725
rect 245745 276722 245811 276725
rect 197353 276720 200284 276722
rect 197353 276664 197358 276720
rect 197414 276664 200284 276720
rect 197353 276662 200284 276664
rect 244076 276720 245811 276722
rect 244076 276664 245750 276720
rect 245806 276664 245811 276720
rect 244076 276662 245811 276664
rect 197353 276659 197419 276662
rect 245745 276659 245811 276662
rect 65926 275980 65932 276044
rect 65996 276042 66002 276044
rect 66069 276042 66135 276045
rect 68878 276042 68938 276148
rect 65996 276040 68938 276042
rect 65996 275984 66074 276040
rect 66130 275984 68938 276040
rect 65996 275982 68938 275984
rect 65996 275980 66002 275982
rect 66069 275979 66135 275982
rect 157057 275906 157123 275909
rect 154652 275904 157123 275906
rect 154652 275848 157062 275904
rect 157118 275848 157123 275904
rect 154652 275846 157123 275848
rect 157057 275843 157123 275846
rect 197445 275906 197511 275909
rect 245929 275906 245995 275909
rect 197445 275904 200284 275906
rect 197445 275848 197450 275904
rect 197506 275848 200284 275904
rect 197445 275846 200284 275848
rect 244076 275904 245995 275906
rect 244076 275848 245934 275904
rect 245990 275848 245995 275904
rect 244076 275846 245995 275848
rect 197445 275843 197511 275846
rect 245929 275843 245995 275846
rect 244222 275634 244228 275636
rect 244046 275574 244228 275634
rect 66805 275362 66871 275365
rect 66805 275360 68908 275362
rect 66805 275304 66810 275360
rect 66866 275304 68908 275360
rect 66805 275302 68908 275304
rect 66805 275299 66871 275302
rect 155166 275300 155172 275364
rect 155236 275362 155242 275364
rect 169017 275362 169083 275365
rect 155236 275360 169083 275362
rect 155236 275304 169022 275360
rect 169078 275304 169083 275360
rect 244046 275332 244106 275574
rect 244222 275572 244228 275574
rect 244292 275572 244298 275636
rect 155236 275302 169083 275304
rect 155236 275300 155242 275302
rect 169017 275299 169083 275302
rect 156689 275226 156755 275229
rect 173014 275226 173020 275228
rect 156689 275224 173020 275226
rect 156689 275168 156694 275224
rect 156750 275168 173020 275224
rect 156689 275166 173020 275168
rect 156689 275163 156755 275166
rect 173014 275164 173020 275166
rect 173084 275164 173090 275228
rect 156873 274818 156939 274821
rect 154652 274816 156939 274818
rect 154652 274760 156878 274816
rect 156934 274760 156939 274816
rect 154652 274758 156939 274760
rect 156873 274755 156939 274758
rect 169201 274818 169267 274821
rect 200254 274818 200314 275060
rect 169201 274816 200314 274818
rect 169201 274760 169206 274816
rect 169262 274760 200314 274816
rect 169201 274758 200314 274760
rect 169201 274755 169267 274758
rect 197537 274546 197603 274549
rect 198641 274546 198707 274549
rect 245653 274546 245719 274549
rect 245837 274546 245903 274549
rect 197537 274544 200284 274546
rect 197537 274488 197542 274544
rect 197598 274488 198646 274544
rect 198702 274488 200284 274544
rect 197537 274486 200284 274488
rect 244076 274544 245903 274546
rect 244076 274488 245658 274544
rect 245714 274488 245842 274544
rect 245898 274488 245903 274544
rect 244076 274486 245903 274488
rect 197537 274483 197603 274486
rect 198641 274483 198707 274486
rect 245653 274483 245719 274486
rect 245837 274483 245903 274486
rect 66805 274274 66871 274277
rect 66805 274272 68908 274274
rect 66805 274216 66810 274272
rect 66866 274216 68908 274272
rect 66805 274214 68908 274216
rect 66805 274211 66871 274214
rect 162301 273866 162367 273869
rect 199561 273866 199627 273869
rect 162301 273864 199627 273866
rect 162301 273808 162306 273864
rect 162362 273808 199566 273864
rect 199622 273808 199627 273864
rect 162301 273806 199627 273808
rect 162301 273803 162367 273806
rect 199561 273803 199627 273806
rect 156505 273730 156571 273733
rect 154652 273728 156571 273730
rect 154652 273672 156510 273728
rect 156566 273672 156571 273728
rect 154652 273670 156571 273672
rect 156505 273667 156571 273670
rect 197353 273730 197419 273733
rect 245837 273730 245903 273733
rect 197353 273728 200284 273730
rect 197353 273672 197358 273728
rect 197414 273672 200284 273728
rect 197353 273670 200284 273672
rect 244076 273728 245903 273730
rect 244076 273672 245842 273728
rect 245898 273672 245903 273728
rect 244076 273670 245903 273672
rect 197353 273667 197419 273670
rect 245837 273667 245903 273670
rect 159357 273322 159423 273325
rect 160686 273322 160692 273324
rect 159357 273320 160692 273322
rect 159357 273264 159362 273320
rect 159418 273264 160692 273320
rect 159357 273262 160692 273264
rect 159357 273259 159423 273262
rect 160686 273260 160692 273262
rect 160756 273260 160762 273324
rect 66989 273186 67055 273189
rect 245745 273186 245811 273189
rect 66989 273184 68908 273186
rect 66989 273128 66994 273184
rect 67050 273128 68908 273184
rect 66989 273126 68908 273128
rect 244076 273184 245811 273186
rect 244076 273128 245750 273184
rect 245806 273128 245811 273184
rect 244076 273126 245811 273128
rect 66989 273123 67055 273126
rect 245745 273123 245811 273126
rect 197353 272914 197419 272917
rect 197353 272912 200284 272914
rect 197353 272856 197358 272912
rect 197414 272856 200284 272912
rect 197353 272854 200284 272856
rect 197353 272851 197419 272854
rect 157149 272642 157215 272645
rect 154652 272640 157215 272642
rect 154652 272584 157154 272640
rect 157210 272584 157215 272640
rect 154652 272582 157215 272584
rect 157149 272579 157215 272582
rect 193857 272370 193923 272373
rect 245929 272370 245995 272373
rect 246481 272370 246547 272373
rect 193857 272368 200284 272370
rect 193857 272312 193862 272368
rect 193918 272312 200284 272368
rect 193857 272310 200284 272312
rect 244076 272368 246547 272370
rect 244076 272312 245934 272368
rect 245990 272312 246486 272368
rect 246542 272312 246547 272368
rect 244076 272310 246547 272312
rect 193857 272307 193923 272310
rect 245929 272307 245995 272310
rect 246481 272307 246547 272310
rect 580349 272234 580415 272237
rect 583520 272234 584960 272324
rect 580349 272232 584960 272234
rect 580349 272176 580354 272232
rect 580410 272176 584960 272232
rect 580349 272174 584960 272176
rect 580349 272171 580415 272174
rect 66069 272098 66135 272101
rect 66069 272096 68908 272098
rect 66069 272040 66074 272096
rect 66130 272040 68908 272096
rect 583520 272084 584960 272174
rect 66069 272038 68908 272040
rect 66069 272035 66135 272038
rect 157241 271554 157307 271557
rect 154652 271552 157307 271554
rect 154652 271496 157246 271552
rect 157302 271496 157307 271552
rect 154652 271494 157307 271496
rect 157241 271491 157307 271494
rect 197813 271554 197879 271557
rect 245837 271554 245903 271557
rect 197813 271552 200284 271554
rect 197813 271496 197818 271552
rect 197874 271496 200284 271552
rect 197813 271494 200284 271496
rect 244076 271552 245903 271554
rect 244076 271496 245842 271552
rect 245898 271496 245903 271552
rect 244076 271494 245903 271496
rect 197813 271491 197879 271494
rect 245837 271491 245903 271494
rect 243997 271282 244063 271285
rect 243997 271280 244106 271282
rect 243997 271224 244002 271280
rect 244058 271224 244106 271280
rect 243997 271219 244106 271224
rect 66897 271010 66963 271013
rect 197353 271010 197419 271013
rect 66897 271008 68908 271010
rect 66897 270952 66902 271008
rect 66958 270952 68908 271008
rect 66897 270950 68908 270952
rect 197353 271008 200284 271010
rect 197353 270952 197358 271008
rect 197414 270952 200284 271008
rect 197353 270950 200284 270952
rect 66897 270947 66963 270950
rect 197353 270947 197419 270950
rect 244046 270602 244106 271219
rect 273294 270602 273300 270604
rect 244046 270542 273300 270602
rect 273294 270540 273300 270542
rect 273364 270540 273370 270604
rect 157241 270466 157307 270469
rect 154652 270464 157307 270466
rect 154652 270408 157246 270464
rect 157302 270408 157307 270464
rect 154652 270406 157307 270408
rect 157241 270403 157307 270406
rect 180793 270466 180859 270469
rect 181253 270466 181319 270469
rect 194869 270466 194935 270469
rect 180793 270464 194935 270466
rect 180793 270408 180798 270464
rect 180854 270408 181258 270464
rect 181314 270408 194874 270464
rect 194930 270408 194935 270464
rect 180793 270406 194935 270408
rect 180793 270403 180859 270406
rect 181253 270403 181319 270406
rect 194869 270403 194935 270406
rect 197353 270194 197419 270197
rect 245929 270194 245995 270197
rect 197353 270192 200284 270194
rect 197353 270136 197358 270192
rect 197414 270136 200284 270192
rect 197353 270134 200284 270136
rect 244076 270192 245995 270194
rect 244076 270136 245934 270192
rect 245990 270136 245995 270192
rect 244076 270134 245995 270136
rect 197353 270131 197419 270134
rect 245929 270131 245995 270134
rect 66713 269922 66779 269925
rect 66713 269920 68908 269922
rect 66713 269864 66718 269920
rect 66774 269864 68908 269920
rect 66713 269862 68908 269864
rect 66713 269859 66779 269862
rect 164969 269786 165035 269789
rect 181253 269786 181319 269789
rect 164969 269784 181319 269786
rect 164969 269728 164974 269784
rect 165030 269728 181258 269784
rect 181314 269728 181319 269784
rect 164969 269726 181319 269728
rect 164969 269723 165035 269726
rect 181253 269723 181319 269726
rect 246021 269650 246087 269653
rect 244076 269648 246087 269650
rect 244076 269592 246026 269648
rect 246082 269592 246087 269648
rect 244076 269590 246087 269592
rect 246021 269587 246087 269590
rect 161974 269378 161980 269380
rect 154652 269318 161980 269378
rect 161974 269316 161980 269318
rect 162044 269316 162050 269380
rect 197445 269378 197511 269381
rect 197445 269376 200284 269378
rect 197445 269320 197450 269376
rect 197506 269320 200284 269376
rect 197445 269318 200284 269320
rect 197445 269315 197511 269318
rect 244917 269106 244983 269109
rect 246665 269106 246731 269109
rect 244046 269104 246731 269106
rect 244046 269048 244922 269104
rect 244978 269048 246670 269104
rect 246726 269048 246731 269104
rect 244046 269046 246731 269048
rect 67633 268834 67699 268837
rect 197353 268834 197419 268837
rect 67633 268832 68908 268834
rect 67633 268776 67638 268832
rect 67694 268776 68908 268832
rect 67633 268774 68908 268776
rect 197353 268832 200284 268834
rect 197353 268776 197358 268832
rect 197414 268776 200284 268832
rect 244046 268804 244106 269046
rect 244917 269043 244983 269046
rect 246665 269043 246731 269046
rect 197353 268774 200284 268776
rect 67633 268771 67699 268774
rect 197353 268771 197419 268774
rect 157241 268290 157307 268293
rect 154652 268288 157307 268290
rect 154652 268232 157246 268288
rect 157302 268232 157307 268288
rect 154652 268230 157307 268232
rect 157241 268227 157307 268230
rect 245745 268018 245811 268021
rect 200070 267958 200284 268018
rect 244076 268016 245811 268018
rect 244076 267960 245750 268016
rect 245806 267960 245811 268016
rect 244076 267958 245811 267960
rect 177389 267882 177455 267885
rect 200070 267882 200130 267958
rect 245745 267955 245811 267958
rect 177389 267880 200130 267882
rect 177389 267824 177394 267880
rect 177450 267824 200130 267880
rect 177389 267822 200130 267824
rect 177389 267819 177455 267822
rect 66253 267746 66319 267749
rect 66253 267744 68908 267746
rect 66253 267688 66258 267744
rect 66314 267688 68908 267744
rect 66253 267686 68908 267688
rect 66253 267683 66319 267686
rect 157241 267474 157307 267477
rect 245837 267474 245903 267477
rect 154652 267472 157307 267474
rect 154652 267416 157246 267472
rect 157302 267416 157307 267472
rect 154652 267414 157307 267416
rect 244076 267472 245903 267474
rect 244076 267416 245842 267472
rect 245898 267416 245903 267472
rect 244076 267414 245903 267416
rect 157241 267411 157307 267414
rect 245837 267411 245903 267414
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 197997 267202 198063 267205
rect 197997 267200 200284 267202
rect 197997 267144 198002 267200
rect 198058 267144 200284 267200
rect 197997 267142 200284 267144
rect 197997 267139 198063 267142
rect 67398 266868 67404 266932
rect 67468 266930 67474 266932
rect 67468 266870 68908 266930
rect 67468 266868 67474 266870
rect 245929 266658 245995 266661
rect 200070 266598 200284 266658
rect 244076 266656 245995 266658
rect 244076 266600 245934 266656
rect 245990 266600 245995 266656
rect 244076 266598 245995 266600
rect 184381 266522 184447 266525
rect 200070 266522 200130 266598
rect 245929 266595 245995 266598
rect 184381 266520 200130 266522
rect 184381 266464 184386 266520
rect 184442 266464 200130 266520
rect 184381 266462 200130 266464
rect 184381 266459 184447 266462
rect 184197 266386 184263 266389
rect 154652 266384 184263 266386
rect 154652 266328 184202 266384
rect 184258 266328 184263 266384
rect 154652 266326 184263 266328
rect 184197 266323 184263 266326
rect 66805 265842 66871 265845
rect 197353 265842 197419 265845
rect 245929 265842 245995 265845
rect 66805 265840 68908 265842
rect 66805 265784 66810 265840
rect 66866 265784 68908 265840
rect 66805 265782 68908 265784
rect 197353 265840 200284 265842
rect 197353 265784 197358 265840
rect 197414 265784 200284 265840
rect 197353 265782 200284 265784
rect 244076 265840 245995 265842
rect 244076 265784 245934 265840
rect 245990 265784 245995 265840
rect 244076 265782 245995 265784
rect 66805 265779 66871 265782
rect 197353 265779 197419 265782
rect 245929 265779 245995 265782
rect 249977 265708 250043 265709
rect 249926 265644 249932 265708
rect 249996 265706 250043 265708
rect 249996 265704 250088 265706
rect 250038 265648 250088 265704
rect 249996 265646 250088 265648
rect 249996 265644 250043 265646
rect 249977 265643 250043 265644
rect 157241 265298 157307 265301
rect 246573 265298 246639 265301
rect 154652 265296 157307 265298
rect 154652 265240 157246 265296
rect 157302 265240 157307 265296
rect 154652 265238 157307 265240
rect 157241 265235 157307 265238
rect 200070 265238 200284 265298
rect 244076 265296 246639 265298
rect 244076 265240 246578 265296
rect 246634 265240 246639 265296
rect 244076 265238 246639 265240
rect 176101 265162 176167 265165
rect 200070 265162 200130 265238
rect 246573 265235 246639 265238
rect 176101 265160 200130 265162
rect 176101 265104 176106 265160
rect 176162 265104 200130 265160
rect 176101 265102 200130 265104
rect 176101 265099 176167 265102
rect 66805 264754 66871 264757
rect 154757 264754 154823 264757
rect 66805 264752 68908 264754
rect 66805 264696 66810 264752
rect 66866 264696 68908 264752
rect 66805 264694 68908 264696
rect 154622 264752 154823 264754
rect 154622 264696 154762 264752
rect 154818 264696 154823 264752
rect 154622 264694 154823 264696
rect 66805 264691 66871 264694
rect 154622 264180 154682 264694
rect 154757 264691 154823 264694
rect 196709 264482 196775 264485
rect 196709 264480 200284 264482
rect 196709 264424 196714 264480
rect 196770 264424 200284 264480
rect 196709 264422 200284 264424
rect 196709 264419 196775 264422
rect 155861 264210 155927 264213
rect 194041 264210 194107 264213
rect 155861 264208 194107 264210
rect 155861 264152 155866 264208
rect 155922 264152 194046 264208
rect 194102 264152 194107 264208
rect 155861 264150 194107 264152
rect 244046 264210 244106 264452
rect 244917 264210 244983 264213
rect 244046 264208 244983 264210
rect 244046 264152 244922 264208
rect 244978 264152 244983 264208
rect 244046 264150 244983 264152
rect 155861 264147 155927 264150
rect 194041 264147 194107 264150
rect 244917 264147 244983 264150
rect 249742 263938 249748 263940
rect 244076 263878 249748 263938
rect 249742 263876 249748 263878
rect 249812 263876 249818 263940
rect 66529 263666 66595 263669
rect 197353 263666 197419 263669
rect 66529 263664 68908 263666
rect 66529 263608 66534 263664
rect 66590 263608 68908 263664
rect 66529 263606 68908 263608
rect 197353 263664 200284 263666
rect 197353 263608 197358 263664
rect 197414 263608 200284 263664
rect 197353 263606 200284 263608
rect 66529 263603 66595 263606
rect 197353 263603 197419 263606
rect 157241 263122 157307 263125
rect 154652 263120 157307 263122
rect 154652 263064 157246 263120
rect 157302 263064 157307 263120
rect 154652 263062 157307 263064
rect 157241 263059 157307 263062
rect 197353 263122 197419 263125
rect 245837 263122 245903 263125
rect 197353 263120 200284 263122
rect 197353 263064 197358 263120
rect 197414 263064 200284 263120
rect 197353 263062 200284 263064
rect 244076 263120 245903 263122
rect 244076 263064 245842 263120
rect 245898 263064 245903 263120
rect 244076 263062 245903 263064
rect 197353 263059 197419 263062
rect 245837 263059 245903 263062
rect 66437 262578 66503 262581
rect 66437 262576 68908 262578
rect 66437 262520 66442 262576
rect 66498 262520 68908 262576
rect 66437 262518 68908 262520
rect 66437 262515 66503 262518
rect 198089 262306 198155 262309
rect 245929 262306 245995 262309
rect 198089 262304 200284 262306
rect 198089 262248 198094 262304
rect 198150 262248 200284 262304
rect 198089 262246 200284 262248
rect 244076 262304 245995 262306
rect 244076 262248 245934 262304
rect 245990 262248 245995 262304
rect 244076 262246 245995 262248
rect 198089 262243 198155 262246
rect 245929 262243 245995 262246
rect 154849 262034 154915 262037
rect 154652 262032 154915 262034
rect 154652 261976 154854 262032
rect 154910 261976 154915 262032
rect 154652 261974 154915 261976
rect 154849 261971 154915 261974
rect 248505 261762 248571 261765
rect 244076 261760 248571 261762
rect 244076 261704 248510 261760
rect 248566 261704 248571 261760
rect 244076 261702 248571 261704
rect 248505 261699 248571 261702
rect 66805 261490 66871 261493
rect 66805 261488 68908 261490
rect 66805 261432 66810 261488
rect 66866 261432 68908 261488
rect 66805 261430 68908 261432
rect 66805 261427 66871 261430
rect 169753 261218 169819 261221
rect 200254 261218 200314 261460
rect 169753 261216 200314 261218
rect 169753 261160 169758 261216
rect 169814 261160 200314 261216
rect 169753 261158 200314 261160
rect 169753 261155 169819 261158
rect 168373 260946 168439 260949
rect 154652 260944 168439 260946
rect 154652 260916 168378 260944
rect 154622 260888 168378 260916
rect 168434 260888 168439 260944
rect 154622 260886 168439 260888
rect 154622 260812 154682 260886
rect 168373 260883 168439 260886
rect 192753 260946 192819 260949
rect 246389 260946 246455 260949
rect 192753 260944 200284 260946
rect 192753 260888 192758 260944
rect 192814 260888 200284 260944
rect 192753 260886 200284 260888
rect 244076 260944 246455 260946
rect 244076 260888 246394 260944
rect 246450 260888 246455 260944
rect 244076 260886 246455 260888
rect 192753 260883 192819 260886
rect 246389 260883 246455 260886
rect 154614 260748 154620 260812
rect 154684 260748 154690 260812
rect 66805 260402 66871 260405
rect 66805 260400 68908 260402
rect 66805 260344 66810 260400
rect 66866 260344 68908 260400
rect 66805 260342 68908 260344
rect 66805 260339 66871 260342
rect 167821 260130 167887 260133
rect 191046 260130 191052 260132
rect 167821 260128 191052 260130
rect 167821 260072 167826 260128
rect 167882 260072 191052 260128
rect 167821 260070 191052 260072
rect 167821 260067 167887 260070
rect 191046 260068 191052 260070
rect 191116 260068 191122 260132
rect 197445 260130 197511 260133
rect 245929 260130 245995 260133
rect 197445 260128 200284 260130
rect 197445 260072 197450 260128
rect 197506 260072 200284 260128
rect 197445 260070 200284 260072
rect 244076 260128 245995 260130
rect 244076 260072 245934 260128
rect 245990 260072 245995 260128
rect 244076 260070 245995 260072
rect 197445 260067 197511 260070
rect 245929 260067 245995 260070
rect 156689 259858 156755 259861
rect 154652 259856 156755 259858
rect 154652 259800 156694 259856
rect 156750 259800 156755 259856
rect 154652 259798 156755 259800
rect 156689 259795 156755 259798
rect 244365 259586 244431 259589
rect 244076 259584 244431 259586
rect 244076 259528 244370 259584
rect 244426 259528 244431 259584
rect 244076 259526 244431 259528
rect 244365 259523 244431 259526
rect 68185 258770 68251 258773
rect 68878 258770 68938 259284
rect 156413 259042 156479 259045
rect 154652 259040 156479 259042
rect 154652 258984 156418 259040
rect 156474 258984 156479 259040
rect 154652 258982 156479 258984
rect 156413 258979 156479 258982
rect 191598 258980 191604 259044
rect 191668 259042 191674 259044
rect 200254 259042 200314 259284
rect 191668 258982 200314 259042
rect 191668 258980 191674 258982
rect 582465 258906 582531 258909
rect 583520 258906 584960 258996
rect 582465 258904 584960 258906
rect 582465 258848 582470 258904
rect 582526 258848 584960 258904
rect 582465 258846 584960 258848
rect 582465 258843 582531 258846
rect 68185 258768 68938 258770
rect 68185 258712 68190 258768
rect 68246 258712 68938 258768
rect 68185 258710 68938 258712
rect 197353 258770 197419 258773
rect 244457 258770 244523 258773
rect 245009 258770 245075 258773
rect 197353 258768 200284 258770
rect 197353 258712 197358 258768
rect 197414 258712 200284 258768
rect 197353 258710 200284 258712
rect 244076 258768 245075 258770
rect 244076 258712 244462 258768
rect 244518 258712 245014 258768
rect 245070 258712 245075 258768
rect 583520 258756 584960 258846
rect 244076 258710 245075 258712
rect 68185 258707 68251 258710
rect 197353 258707 197419 258710
rect 244457 258707 244523 258710
rect 245009 258707 245075 258710
rect 66713 258498 66779 258501
rect 66713 258496 68908 258498
rect 66713 258440 66718 258496
rect 66774 258440 68908 258496
rect 66713 258438 68908 258440
rect 66713 258435 66779 258438
rect 245929 258226 245995 258229
rect 244076 258224 245995 258226
rect 244076 258168 245934 258224
rect 245990 258168 245995 258224
rect 244076 258166 245995 258168
rect 245929 258163 245995 258166
rect 156873 257954 156939 257957
rect 154652 257952 156939 257954
rect 154652 257896 156878 257952
rect 156934 257896 156939 257952
rect 154652 257894 156939 257896
rect 156873 257891 156939 257894
rect 197353 257954 197419 257957
rect 197353 257952 200284 257954
rect 197353 257896 197358 257952
rect 197414 257896 200284 257952
rect 197353 257894 200284 257896
rect 197353 257891 197419 257894
rect 200021 257410 200087 257413
rect 247125 257410 247191 257413
rect 200021 257408 200284 257410
rect 69430 256868 69490 257380
rect 200021 257352 200026 257408
rect 200082 257352 200284 257408
rect 200021 257350 200284 257352
rect 244076 257408 247191 257410
rect 244076 257352 247130 257408
rect 247186 257352 247191 257408
rect 244076 257350 247191 257352
rect 200021 257347 200087 257350
rect 247125 257347 247191 257350
rect 69422 256804 69428 256868
rect 69492 256804 69498 256868
rect 157241 256866 157307 256869
rect 154652 256864 157307 256866
rect 154652 256808 157246 256864
rect 157302 256808 157307 256864
rect 154652 256806 157307 256808
rect 157241 256803 157307 256806
rect 198641 256594 198707 256597
rect 245653 256594 245719 256597
rect 198641 256592 200284 256594
rect 198641 256536 198646 256592
rect 198702 256536 200284 256592
rect 198641 256534 200284 256536
rect 244076 256592 245719 256594
rect 244076 256536 245658 256592
rect 245714 256536 245719 256592
rect 244076 256534 245719 256536
rect 198641 256531 198707 256534
rect 245653 256531 245719 256534
rect 67950 256260 67956 256324
rect 68020 256322 68026 256324
rect 68020 256262 68908 256322
rect 68020 256260 68026 256262
rect 246941 256050 247007 256053
rect 244076 256048 247007 256050
rect 244076 255992 246946 256048
rect 247002 255992 247007 256048
rect 244076 255990 247007 255992
rect 246941 255987 247007 255990
rect 157241 255778 157307 255781
rect 154652 255776 157307 255778
rect 154652 255720 157246 255776
rect 157302 255720 157307 255776
rect 154652 255718 157307 255720
rect 157241 255715 157307 255718
rect 197353 255778 197419 255781
rect 197353 255776 200284 255778
rect 197353 255720 197358 255776
rect 197414 255720 200284 255776
rect 197353 255718 200284 255720
rect 197353 255715 197419 255718
rect 67633 255234 67699 255237
rect 195973 255234 196039 255237
rect 197118 255234 197124 255236
rect 67633 255232 68908 255234
rect 67633 255176 67638 255232
rect 67694 255176 68908 255232
rect 67633 255174 68908 255176
rect 195973 255232 197124 255234
rect 195973 255176 195978 255232
rect 196034 255176 197124 255232
rect 195973 255174 197124 255176
rect 67633 255171 67699 255174
rect 195973 255171 196039 255174
rect 197118 255172 197124 255174
rect 197188 255234 197194 255236
rect 246941 255234 247007 255237
rect 197188 255174 200284 255234
rect 244076 255232 247007 255234
rect 244076 255176 246946 255232
rect 247002 255176 247007 255232
rect 244076 255174 247007 255176
rect 197188 255172 197194 255174
rect 246941 255171 247007 255174
rect 157241 254690 157307 254693
rect 154652 254688 157307 254690
rect 154652 254632 157246 254688
rect 157302 254632 157307 254688
rect 154652 254630 157307 254632
rect 157241 254627 157307 254630
rect 197353 254418 197419 254421
rect 197353 254416 200284 254418
rect 197353 254360 197358 254416
rect 197414 254360 200284 254416
rect 197353 254358 200284 254360
rect 197353 254355 197419 254358
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 66897 254146 66963 254149
rect 244046 254146 244106 254388
rect 255497 254146 255563 254149
rect 66897 254144 68908 254146
rect 66897 254088 66902 254144
rect 66958 254088 68908 254144
rect 66897 254086 68908 254088
rect 244046 254144 255563 254146
rect 244046 254088 255502 254144
rect 255558 254088 255563 254144
rect 244046 254086 255563 254088
rect 66897 254083 66963 254086
rect 255497 254083 255563 254086
rect 174629 253874 174695 253877
rect 181437 253874 181503 253877
rect 245929 253874 245995 253877
rect 174629 253872 181503 253874
rect 174629 253816 174634 253872
rect 174690 253816 181442 253872
rect 181498 253816 181503 253872
rect 174629 253814 181503 253816
rect 244076 253872 245995 253874
rect 244076 253816 245934 253872
rect 245990 253816 245995 253872
rect 244076 253814 245995 253816
rect 174629 253811 174695 253814
rect 181437 253811 181503 253814
rect 245929 253811 245995 253814
rect 156413 253602 156479 253605
rect 154652 253600 156479 253602
rect 154652 253544 156418 253600
rect 156474 253544 156479 253600
rect 154652 253542 156479 253544
rect 156413 253539 156479 253542
rect 197445 253602 197511 253605
rect 197445 253600 200284 253602
rect 197445 253544 197450 253600
rect 197506 253544 200284 253600
rect 197445 253542 200284 253544
rect 197445 253539 197511 253542
rect 66897 253058 66963 253061
rect 197353 253058 197419 253061
rect 245653 253058 245719 253061
rect 66897 253056 68908 253058
rect 66897 253000 66902 253056
rect 66958 253000 68908 253056
rect 66897 252998 68908 253000
rect 197353 253056 200284 253058
rect 197353 253000 197358 253056
rect 197414 253000 200284 253056
rect 197353 252998 200284 253000
rect 244076 253056 245719 253058
rect 244076 253000 245658 253056
rect 245714 253000 245719 253056
rect 244076 252998 245719 253000
rect 66897 252995 66963 252998
rect 197353 252995 197419 252998
rect 245653 252995 245719 252998
rect 66662 251908 66668 251972
rect 66732 251970 66738 251972
rect 154622 251970 154682 252484
rect 197353 252242 197419 252245
rect 245929 252242 245995 252245
rect 197353 252240 200284 252242
rect 197353 252184 197358 252240
rect 197414 252184 200284 252240
rect 197353 252182 200284 252184
rect 244076 252240 245995 252242
rect 244076 252184 245934 252240
rect 245990 252184 245995 252240
rect 244076 252182 245995 252184
rect 197353 252179 197419 252182
rect 245929 252179 245995 252182
rect 199878 251970 199884 251972
rect 66732 251910 68908 251970
rect 154622 251910 199884 251970
rect 66732 251908 66738 251910
rect 199878 251908 199884 251910
rect 199948 251908 199954 251972
rect 197445 251698 197511 251701
rect 246021 251698 246087 251701
rect 197445 251696 200284 251698
rect 197445 251640 197450 251696
rect 197506 251640 200284 251696
rect 197445 251638 200284 251640
rect 244076 251696 246087 251698
rect 244076 251640 246026 251696
rect 246082 251640 246087 251696
rect 244076 251638 246087 251640
rect 197445 251635 197511 251638
rect 246021 251635 246087 251638
rect 168414 251426 168420 251428
rect 154652 251366 168420 251426
rect 168414 251364 168420 251366
rect 168484 251364 168490 251428
rect 197353 250882 197419 250885
rect 244273 250882 244339 250885
rect 197353 250880 200284 250882
rect 67909 250338 67975 250341
rect 68878 250338 68938 250852
rect 197353 250824 197358 250880
rect 197414 250824 200284 250880
rect 197353 250822 200284 250824
rect 244076 250880 244339 250882
rect 244076 250824 244278 250880
rect 244334 250824 244339 250880
rect 244076 250822 244339 250824
rect 197353 250819 197419 250822
rect 244273 250819 244339 250822
rect 157241 250610 157307 250613
rect 154652 250608 157307 250610
rect 154652 250552 157246 250608
rect 157302 250552 157307 250608
rect 154652 250550 157307 250552
rect 157241 250547 157307 250550
rect 245653 250338 245719 250341
rect 67909 250336 68938 250338
rect 67909 250280 67914 250336
rect 67970 250280 68938 250336
rect 67909 250278 68938 250280
rect 244076 250336 245719 250338
rect 244076 250280 245658 250336
rect 245714 250280 245719 250336
rect 244076 250278 245719 250280
rect 67909 250275 67975 250278
rect 245653 250275 245719 250278
rect 65885 250066 65951 250069
rect 65885 250064 68908 250066
rect 65885 250008 65890 250064
rect 65946 250008 68908 250064
rect 65885 250006 68908 250008
rect 200070 250006 200284 250066
rect 65885 250003 65951 250006
rect 169109 249930 169175 249933
rect 200070 249930 200130 250006
rect 169109 249928 200130 249930
rect 169109 249872 169114 249928
rect 169170 249872 200130 249928
rect 169109 249870 200130 249872
rect 169109 249867 169175 249870
rect 199469 249796 199535 249797
rect 199469 249792 199516 249796
rect 199580 249794 199586 249796
rect 199469 249736 199474 249792
rect 199469 249732 199516 249736
rect 199580 249734 199626 249794
rect 199580 249732 199586 249734
rect 199469 249731 199535 249732
rect 156413 249522 156479 249525
rect 154652 249520 156479 249522
rect 154652 249464 156418 249520
rect 156474 249464 156479 249520
rect 154652 249462 156479 249464
rect 156413 249459 156479 249462
rect 197353 249522 197419 249525
rect 248454 249522 248460 249524
rect 197353 249520 200284 249522
rect 197353 249464 197358 249520
rect 197414 249464 200284 249520
rect 197353 249462 200284 249464
rect 244076 249462 248460 249522
rect 197353 249459 197419 249462
rect 248454 249460 248460 249462
rect 248524 249460 248530 249524
rect 178953 249114 179019 249117
rect 187509 249114 187575 249117
rect 178953 249112 187575 249114
rect 178953 249056 178958 249112
rect 179014 249056 187514 249112
rect 187570 249056 187575 249112
rect 178953 249054 187575 249056
rect 178953 249051 179019 249054
rect 187509 249051 187575 249054
rect 66805 248978 66871 248981
rect 66805 248976 68908 248978
rect 66805 248920 66810 248976
rect 66866 248920 68908 248976
rect 66805 248918 68908 248920
rect 66805 248915 66871 248918
rect 245745 248706 245811 248709
rect 200070 248646 200284 248706
rect 244076 248704 245811 248706
rect 244076 248648 245750 248704
rect 245806 248648 245811 248704
rect 244076 248646 245811 248648
rect 187509 248570 187575 248573
rect 200070 248570 200130 248646
rect 245745 248643 245811 248646
rect 187509 248568 200130 248570
rect 187509 248512 187514 248568
rect 187570 248512 200130 248568
rect 187509 248510 200130 248512
rect 187509 248507 187575 248510
rect 157149 248434 157215 248437
rect 154652 248432 157215 248434
rect 154652 248376 157154 248432
rect 157210 248376 157215 248432
rect 154652 248374 157215 248376
rect 157149 248371 157215 248374
rect 245929 248162 245995 248165
rect 244076 248160 245995 248162
rect 244076 248104 245934 248160
rect 245990 248104 245995 248160
rect 244076 248102 245995 248104
rect 245929 248099 245995 248102
rect 66621 247890 66687 247893
rect 197445 247890 197511 247893
rect 66621 247888 68908 247890
rect 66621 247832 66626 247888
rect 66682 247832 68908 247888
rect 66621 247830 68908 247832
rect 197445 247888 200284 247890
rect 197445 247832 197450 247888
rect 197506 247832 200284 247888
rect 197445 247830 200284 247832
rect 66621 247827 66687 247830
rect 197445 247827 197511 247830
rect 156781 247346 156847 247349
rect 244457 247346 244523 247349
rect 154652 247344 156847 247346
rect 154652 247288 156786 247344
rect 156842 247288 156847 247344
rect 154652 247286 156847 247288
rect 156781 247283 156847 247286
rect 200070 247286 200284 247346
rect 244076 247344 244523 247346
rect 244076 247288 244462 247344
rect 244518 247288 244523 247344
rect 244076 247286 244523 247288
rect 186998 247148 187004 247212
rect 187068 247210 187074 247212
rect 200070 247210 200130 247286
rect 244457 247283 244523 247286
rect 187068 247150 200130 247210
rect 187068 247148 187074 247150
rect 67265 246802 67331 246805
rect 67265 246800 68908 246802
rect 67265 246744 67270 246800
rect 67326 246744 68908 246800
rect 67265 246742 68908 246744
rect 67265 246739 67331 246742
rect 199878 246468 199884 246532
rect 199948 246530 199954 246532
rect 199948 246470 200284 246530
rect 199948 246468 199954 246470
rect 67725 245714 67791 245717
rect 154622 245714 154682 246228
rect 160686 246196 160692 246260
rect 160756 246258 160762 246260
rect 170397 246258 170463 246261
rect 243494 246260 243554 246500
rect 160756 246256 170463 246258
rect 160756 246200 170402 246256
rect 170458 246200 170463 246256
rect 160756 246198 170463 246200
rect 160756 246196 160762 246198
rect 170397 246195 170463 246198
rect 243486 246196 243492 246260
rect 243556 246196 243562 246260
rect 197353 245986 197419 245989
rect 245929 245986 245995 245989
rect 197353 245984 200284 245986
rect 197353 245928 197358 245984
rect 197414 245928 200284 245984
rect 197353 245926 200284 245928
rect 244076 245984 245995 245986
rect 244076 245928 245934 245984
rect 245990 245928 245995 245984
rect 244076 245926 245995 245928
rect 197353 245923 197419 245926
rect 245929 245923 245995 245926
rect 162209 245714 162275 245717
rect 67725 245712 68908 245714
rect 67725 245656 67730 245712
rect 67786 245656 68908 245712
rect 67725 245654 68908 245656
rect 154622 245712 162275 245714
rect 154622 245656 162214 245712
rect 162270 245656 162275 245712
rect 154622 245654 162275 245656
rect 67725 245651 67791 245654
rect 162209 245651 162275 245654
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 66621 245170 66687 245173
rect 69422 245170 69428 245172
rect 66621 245168 69428 245170
rect 66621 245112 66626 245168
rect 66682 245112 69428 245168
rect 66621 245110 69428 245112
rect 66621 245107 66687 245110
rect 69422 245108 69428 245110
rect 69492 245108 69498 245172
rect 156965 245170 157031 245173
rect 154652 245168 157031 245170
rect 154652 245112 156970 245168
rect 157026 245112 157031 245168
rect 154652 245110 157031 245112
rect 69430 244596 69490 245108
rect 156965 245107 157031 245110
rect 197353 245170 197419 245173
rect 245653 245170 245719 245173
rect 197353 245168 200284 245170
rect 197353 245112 197358 245168
rect 197414 245112 200284 245168
rect 197353 245110 200284 245112
rect 244076 245168 245719 245170
rect 244076 245112 245658 245168
rect 245714 245112 245719 245168
rect 244076 245110 245719 245112
rect 197353 245107 197419 245110
rect 245653 245107 245719 245110
rect 189717 244898 189783 244901
rect 194409 244898 194475 244901
rect 189717 244896 200314 244898
rect 189717 244840 189722 244896
rect 189778 244840 194414 244896
rect 194470 244840 200314 244896
rect 189717 244838 200314 244840
rect 189717 244835 189783 244838
rect 194409 244835 194475 244838
rect 154430 244428 154436 244492
rect 154500 244490 154506 244492
rect 191097 244490 191163 244493
rect 154500 244488 191163 244490
rect 154500 244432 191102 244488
rect 191158 244432 191163 244488
rect 154500 244430 191163 244432
rect 154500 244428 154506 244430
rect 191097 244427 191163 244430
rect 200254 244324 200314 244838
rect 247125 244626 247191 244629
rect 244076 244624 247191 244626
rect 244076 244568 247130 244624
rect 247186 244568 247191 244624
rect 244076 244566 247191 244568
rect 247125 244563 247191 244566
rect 156045 244082 156111 244085
rect 154652 244080 156111 244082
rect 154652 244024 156050 244080
rect 156106 244024 156111 244080
rect 154652 244022 156111 244024
rect 156045 244019 156111 244022
rect 196709 243810 196775 243813
rect 245929 243810 245995 243813
rect 196709 243808 200284 243810
rect 196709 243752 196714 243808
rect 196770 243752 200284 243808
rect 244076 243808 245995 243810
rect 244076 243780 245934 243808
rect 196709 243750 200284 243752
rect 244046 243752 245934 243780
rect 245990 243752 245995 243808
rect 244046 243750 245995 243752
rect 196709 243747 196775 243750
rect 66110 243476 66116 243540
rect 66180 243538 66186 243540
rect 162393 243538 162459 243541
rect 199878 243538 199884 243540
rect 66180 243478 68908 243538
rect 162393 243536 199884 243538
rect 162393 243480 162398 243536
rect 162454 243480 199884 243536
rect 162393 243478 199884 243480
rect 66180 243476 66186 243478
rect 162393 243475 162459 243478
rect 199878 243476 199884 243478
rect 199948 243476 199954 243540
rect 244046 243269 244106 243750
rect 245929 243747 245995 243750
rect 243997 243264 244106 243269
rect 243997 243208 244002 243264
rect 244058 243208 244106 243264
rect 243997 243206 244106 243208
rect 243997 243203 244063 243206
rect 155217 242994 155283 242997
rect 154652 242992 155283 242994
rect 154652 242936 155222 242992
rect 155278 242936 155283 242992
rect 154652 242934 155283 242936
rect 155217 242931 155283 242934
rect 195278 242932 195284 242996
rect 195348 242994 195354 242996
rect 245878 242994 245884 242996
rect 195348 242934 200284 242994
rect 244076 242934 245884 242994
rect 195348 242932 195354 242934
rect 245878 242932 245884 242934
rect 245948 242932 245954 242996
rect 67173 242858 67239 242861
rect 67398 242858 67404 242860
rect 67173 242856 67404 242858
rect 67173 242800 67178 242856
rect 67234 242800 67404 242856
rect 67173 242798 67404 242800
rect 67173 242795 67239 242798
rect 67398 242796 67404 242798
rect 67468 242796 67474 242860
rect 246389 242450 246455 242453
rect 244076 242448 246455 242450
rect 60457 242042 60523 242045
rect 69430 242042 69490 242420
rect 244076 242392 246394 242448
rect 246450 242392 246455 242448
rect 244076 242390 246455 242392
rect 246389 242387 246455 242390
rect 156873 242178 156939 242181
rect 154652 242176 156939 242178
rect 154652 242120 156878 242176
rect 156934 242120 156939 242176
rect 154652 242118 156939 242120
rect 156873 242115 156939 242118
rect 197261 242178 197327 242181
rect 197261 242176 200284 242178
rect 197261 242120 197266 242176
rect 197322 242120 200284 242176
rect 197261 242118 200284 242120
rect 197261 242115 197327 242118
rect 70301 242042 70367 242045
rect 135989 242044 136055 242045
rect 135989 242042 136036 242044
rect 60457 242040 64890 242042
rect 60457 241984 60462 242040
rect 60518 241984 64890 242040
rect 60457 241982 64890 241984
rect 69430 242040 70367 242042
rect 69430 241984 70306 242040
rect 70362 241984 70367 242040
rect 69430 241982 70367 241984
rect 135944 242040 136036 242042
rect 135944 241984 135994 242040
rect 135944 241982 136036 241984
rect 60457 241979 60523 241982
rect 64830 241906 64890 241982
rect 70301 241979 70367 241982
rect 135989 241980 136036 241982
rect 136100 241980 136106 242044
rect 136582 241980 136588 242044
rect 136652 242042 136658 242044
rect 136909 242042 136975 242045
rect 136652 242040 136975 242042
rect 136652 241984 136914 242040
rect 136970 241984 136975 242040
rect 136652 241982 136975 241984
rect 136652 241980 136658 241982
rect 135989 241979 136055 241980
rect 136909 241979 136975 241982
rect 138054 241980 138060 242044
rect 138124 242042 138130 242044
rect 138197 242042 138263 242045
rect 138124 242040 138263 242042
rect 138124 241984 138202 242040
rect 138258 241984 138263 242040
rect 138124 241982 138263 241984
rect 138124 241980 138130 241982
rect 138197 241979 138263 241982
rect 146753 242042 146819 242045
rect 147438 242042 147444 242044
rect 146753 242040 147444 242042
rect 146753 241984 146758 242040
rect 146814 241984 147444 242040
rect 146753 241982 147444 241984
rect 146753 241979 146819 241982
rect 147438 241980 147444 241982
rect 147508 241980 147514 242044
rect 69657 241906 69723 241909
rect 64830 241904 69723 241906
rect 64830 241848 69662 241904
rect 69718 241848 69723 241904
rect 64830 241846 69723 241848
rect 69657 241843 69723 241846
rect 154021 241770 154087 241773
rect 198089 241770 198155 241773
rect 154021 241768 198155 241770
rect 154021 241712 154026 241768
rect 154082 241712 198094 241768
rect 198150 241712 198155 241768
rect 154021 241710 198155 241712
rect 154021 241707 154087 241710
rect 198089 241707 198155 241710
rect 197353 241634 197419 241637
rect 197353 241632 200284 241634
rect 197353 241576 197358 241632
rect 197414 241576 200284 241632
rect 197353 241574 200284 241576
rect 197353 241571 197419 241574
rect 64505 241498 64571 241501
rect 154849 241498 154915 241501
rect 64505 241496 154915 241498
rect 64505 241440 64510 241496
rect 64566 241440 154854 241496
rect 154910 241440 154915 241496
rect 64505 241438 154915 241440
rect 64505 241435 64571 241438
rect 154849 241435 154915 241438
rect 244046 241365 244106 241604
rect 57789 241362 57855 241365
rect 82951 241362 83017 241365
rect 57789 241360 83290 241362
rect 57789 241304 57794 241360
rect 57850 241304 82956 241360
rect 83012 241304 83290 241360
rect 57789 241302 83290 241304
rect 57789 241299 57855 241302
rect 82951 241299 83017 241302
rect 83230 241226 83290 241302
rect 83406 241300 83412 241364
rect 83476 241362 83482 241364
rect 93853 241362 93919 241365
rect 94359 241362 94425 241365
rect 83476 241360 94425 241362
rect 83476 241304 93858 241360
rect 93914 241304 94364 241360
rect 94420 241304 94425 241360
rect 83476 241302 94425 241304
rect 83476 241300 83482 241302
rect 93853 241299 93919 241302
rect 94359 241299 94425 241302
rect 118647 241362 118713 241365
rect 198641 241362 198707 241365
rect 118647 241360 198707 241362
rect 118647 241304 118652 241360
rect 118708 241304 198646 241360
rect 198702 241304 198707 241360
rect 118647 241302 198707 241304
rect 118647 241299 118713 241302
rect 198641 241299 198707 241302
rect 243997 241360 244106 241365
rect 243997 241304 244002 241360
rect 244058 241304 244106 241360
rect 243997 241302 244106 241304
rect 243997 241299 244063 241302
rect 84101 241226 84167 241229
rect 83230 241224 84167 241226
rect -960 241090 480 241180
rect 83230 241168 84106 241224
rect 84162 241168 84167 241224
rect 83230 241166 84167 241168
rect 84101 241163 84167 241166
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 156873 240818 156939 240821
rect 169293 240818 169359 240821
rect 156873 240816 169359 240818
rect 156873 240760 156878 240816
rect 156934 240760 169298 240816
rect 169354 240760 169359 240816
rect 156873 240758 169359 240760
rect 156873 240755 156939 240758
rect 169293 240755 169359 240758
rect 193949 240818 194015 240821
rect 199929 240818 199995 240821
rect 244365 240818 244431 240821
rect 193949 240816 200284 240818
rect 193949 240760 193954 240816
rect 194010 240760 199934 240816
rect 199990 240760 200284 240816
rect 193949 240758 200284 240760
rect 244076 240816 244431 240818
rect 244076 240760 244370 240816
rect 244426 240760 244431 240816
rect 244076 240758 244431 240760
rect 193949 240755 194015 240758
rect 199929 240755 199995 240758
rect 244365 240755 244431 240758
rect 199561 240274 199627 240277
rect 245694 240274 245700 240276
rect 199561 240272 200866 240274
rect 199561 240216 199566 240272
rect 199622 240216 200866 240272
rect 199561 240214 200866 240216
rect 244076 240214 245700 240274
rect 199561 240211 199627 240214
rect 50889 240138 50955 240141
rect 75177 240138 75243 240141
rect 75453 240138 75519 240141
rect 50889 240136 75519 240138
rect 50889 240080 50894 240136
rect 50950 240080 75182 240136
rect 75238 240080 75458 240136
rect 75514 240080 75519 240136
rect 50889 240078 75519 240080
rect 200806 240138 200866 240214
rect 245694 240212 245700 240214
rect 245764 240212 245770 240276
rect 201125 240138 201191 240141
rect 200806 240136 201191 240138
rect 200806 240080 201130 240136
rect 201186 240080 201191 240136
rect 200806 240078 201191 240080
rect 50889 240075 50955 240078
rect 75177 240075 75243 240078
rect 75453 240075 75519 240078
rect 201125 240075 201191 240078
rect 214230 240076 214236 240140
rect 214300 240138 214306 240140
rect 215109 240138 215175 240141
rect 221089 240140 221155 240141
rect 224953 240140 225019 240141
rect 229737 240140 229803 240141
rect 221038 240138 221044 240140
rect 214300 240136 215175 240138
rect 214300 240080 215114 240136
rect 215170 240080 215175 240136
rect 214300 240078 215175 240080
rect 220998 240078 221044 240138
rect 221108 240136 221155 240140
rect 224902 240138 224908 240140
rect 221150 240080 221155 240136
rect 214300 240076 214306 240078
rect 215109 240075 215175 240078
rect 221038 240076 221044 240078
rect 221108 240076 221155 240080
rect 224862 240078 224908 240138
rect 224972 240136 225019 240140
rect 229686 240138 229692 240140
rect 225014 240080 225019 240136
rect 224902 240076 224908 240078
rect 224972 240076 225019 240080
rect 229646 240078 229692 240138
rect 229756 240136 229803 240140
rect 229798 240080 229803 240136
rect 229686 240076 229692 240078
rect 229756 240076 229803 240080
rect 230422 240076 230428 240140
rect 230492 240138 230498 240140
rect 230565 240138 230631 240141
rect 230492 240136 230631 240138
rect 230492 240080 230570 240136
rect 230626 240080 230631 240136
rect 230492 240078 230631 240080
rect 230492 240076 230498 240078
rect 221089 240075 221155 240076
rect 224953 240075 225019 240076
rect 229737 240075 229803 240076
rect 230565 240075 230631 240078
rect 237414 240076 237420 240140
rect 237484 240138 237490 240140
rect 237925 240138 237991 240141
rect 262213 240138 262279 240141
rect 580165 240138 580231 240141
rect 237484 240136 237991 240138
rect 237484 240080 237930 240136
rect 237986 240080 237991 240136
rect 237484 240078 237991 240080
rect 237484 240076 237490 240078
rect 237925 240075 237991 240078
rect 258030 240136 580231 240138
rect 258030 240080 262218 240136
rect 262274 240080 580170 240136
rect 580226 240080 580231 240136
rect 258030 240078 580231 240080
rect 56317 240002 56383 240005
rect 154430 240002 154436 240004
rect 56317 240000 154436 240002
rect 56317 239944 56322 240000
rect 56378 239944 154436 240000
rect 56317 239942 154436 239944
rect 56317 239939 56383 239942
rect 154430 239940 154436 239942
rect 154500 239940 154506 240004
rect 182725 240002 182791 240005
rect 204437 240002 204503 240005
rect 182725 240000 204503 240002
rect 182725 239944 182730 240000
rect 182786 239944 204442 240000
rect 204498 239944 204503 240000
rect 182725 239942 204503 239944
rect 182725 239939 182791 239942
rect 204437 239939 204503 239942
rect 239213 240002 239279 240005
rect 258030 240002 258090 240078
rect 262213 240075 262279 240078
rect 580165 240075 580231 240078
rect 239213 240000 258090 240002
rect 239213 239944 239218 240000
rect 239274 239944 258090 240000
rect 239213 239942 258090 239944
rect 239213 239939 239279 239942
rect 67357 239866 67423 239869
rect 72417 239866 72483 239869
rect 67357 239864 72483 239866
rect 67357 239808 67362 239864
rect 67418 239808 72422 239864
rect 72478 239808 72483 239864
rect 67357 239806 72483 239808
rect 67357 239803 67423 239806
rect 72417 239803 72483 239806
rect 141785 239866 141851 239869
rect 173801 239866 173867 239869
rect 141785 239864 173867 239866
rect 141785 239808 141790 239864
rect 141846 239808 173806 239864
rect 173862 239808 173867 239864
rect 141785 239806 173867 239808
rect 141785 239803 141851 239806
rect 173801 239803 173867 239806
rect 240869 239866 240935 239869
rect 243997 239866 244063 239869
rect 240869 239864 244063 239866
rect 240869 239808 240874 239864
rect 240930 239808 244002 239864
rect 244058 239808 244063 239864
rect 240869 239806 244063 239808
rect 240869 239803 240935 239806
rect 243997 239803 244063 239806
rect 126145 239730 126211 239733
rect 228725 239730 228791 239733
rect 229001 239730 229067 239733
rect 126145 239728 229067 239730
rect 126145 239672 126150 239728
rect 126206 239672 228730 239728
rect 228786 239672 229006 239728
rect 229062 239672 229067 239728
rect 126145 239670 229067 239672
rect 126145 239667 126211 239670
rect 228725 239667 228791 239670
rect 229001 239667 229067 239670
rect 72601 239458 72667 239461
rect 84837 239458 84903 239461
rect 72601 239456 84903 239458
rect 72601 239400 72606 239456
rect 72662 239400 84842 239456
rect 84898 239400 84903 239456
rect 72601 239398 84903 239400
rect 72601 239395 72667 239398
rect 84837 239395 84903 239398
rect 199878 239396 199884 239460
rect 199948 239458 199954 239460
rect 204161 239458 204227 239461
rect 199948 239456 204227 239458
rect 199948 239400 204166 239456
rect 204222 239400 204227 239456
rect 199948 239398 204227 239400
rect 199948 239396 199954 239398
rect 204161 239395 204227 239398
rect 208301 239458 208367 239461
rect 238017 239458 238083 239461
rect 208301 239456 238083 239458
rect 208301 239400 208306 239456
rect 208362 239400 238022 239456
rect 238078 239400 238083 239456
rect 208301 239398 238083 239400
rect 208301 239395 208367 239398
rect 238017 239395 238083 239398
rect 200205 238778 200271 238781
rect 199886 238776 200271 238778
rect 199886 238720 200210 238776
rect 200266 238720 200271 238776
rect 199886 238718 200271 238720
rect 71405 238642 71471 238645
rect 199886 238642 199946 238718
rect 200205 238715 200271 238718
rect 71405 238640 199946 238642
rect 71405 238584 71410 238640
rect 71466 238584 199946 238640
rect 71405 238582 199946 238584
rect 200113 238642 200179 238645
rect 208301 238642 208367 238645
rect 200113 238640 208367 238642
rect 200113 238584 200118 238640
rect 200174 238584 208306 238640
rect 208362 238584 208367 238640
rect 200113 238582 208367 238584
rect 71405 238579 71471 238582
rect 200113 238579 200179 238582
rect 208301 238579 208367 238582
rect 212574 238580 212580 238644
rect 212644 238642 212650 238644
rect 213637 238642 213703 238645
rect 212644 238640 213703 238642
rect 212644 238584 213642 238640
rect 213698 238584 213703 238640
rect 212644 238582 213703 238584
rect 212644 238580 212650 238582
rect 213637 238579 213703 238582
rect 219525 238642 219591 238645
rect 222326 238642 222332 238644
rect 219525 238640 222332 238642
rect 219525 238584 219530 238640
rect 219586 238584 222332 238640
rect 219525 238582 222332 238584
rect 219525 238579 219591 238582
rect 222326 238580 222332 238582
rect 222396 238580 222402 238644
rect 232446 238580 232452 238644
rect 232516 238642 232522 238644
rect 235901 238642 235967 238645
rect 232516 238640 235967 238642
rect 232516 238584 235906 238640
rect 235962 238584 235967 238640
rect 232516 238582 235967 238584
rect 232516 238580 232522 238582
rect 235901 238579 235967 238582
rect 241646 238580 241652 238644
rect 241716 238642 241722 238644
rect 242157 238642 242223 238645
rect 241716 238640 242223 238642
rect 241716 238584 242162 238640
rect 242218 238584 242223 238640
rect 241716 238582 242223 238584
rect 241716 238580 241722 238582
rect 242157 238579 242223 238582
rect 53649 238506 53715 238509
rect 76557 238506 76623 238509
rect 53649 238504 76623 238506
rect 53649 238448 53654 238504
rect 53710 238448 76562 238504
rect 76618 238448 76623 238504
rect 53649 238446 76623 238448
rect 53649 238443 53715 238446
rect 76557 238443 76623 238446
rect 122925 238506 122991 238509
rect 226701 238506 226767 238509
rect 242801 238506 242867 238509
rect 122925 238504 242867 238506
rect 122925 238448 122930 238504
rect 122986 238448 226706 238504
rect 226762 238448 242806 238504
rect 242862 238448 242867 238504
rect 122925 238446 242867 238448
rect 122925 238443 122991 238446
rect 226701 238443 226767 238446
rect 242801 238443 242867 238446
rect 211654 238308 211660 238372
rect 211724 238370 211730 238372
rect 214557 238370 214623 238373
rect 211724 238368 214623 238370
rect 211724 238312 214562 238368
rect 214618 238312 214623 238368
rect 211724 238310 214623 238312
rect 211724 238308 211730 238310
rect 214557 238307 214623 238310
rect 235349 238370 235415 238373
rect 255405 238370 255471 238373
rect 235349 238368 255471 238370
rect 235349 238312 235354 238368
rect 235410 238312 255410 238368
rect 255466 238312 255471 238368
rect 235349 238310 255471 238312
rect 235349 238307 235415 238310
rect 255405 238307 255471 238310
rect 200614 237900 200620 237964
rect 200684 237962 200690 237964
rect 231761 237962 231827 237965
rect 200684 237960 231827 237962
rect 200684 237904 231766 237960
rect 231822 237904 231827 237960
rect 200684 237902 231827 237904
rect 200684 237900 200690 237902
rect 231761 237899 231827 237902
rect 255405 237962 255471 237965
rect 582833 237962 582899 237965
rect 255405 237960 582899 237962
rect 255405 237904 255410 237960
rect 255466 237904 582838 237960
rect 582894 237904 582899 237960
rect 255405 237902 582899 237904
rect 255405 237899 255471 237902
rect 582833 237899 582899 237902
rect 200205 237418 200271 237421
rect 200757 237418 200823 237421
rect 213085 237420 213151 237421
rect 213085 237418 213132 237420
rect 200205 237416 200823 237418
rect 200205 237360 200210 237416
rect 200266 237360 200762 237416
rect 200818 237360 200823 237416
rect 200205 237358 200823 237360
rect 213040 237416 213132 237418
rect 213040 237360 213090 237416
rect 213040 237358 213132 237360
rect 200205 237355 200271 237358
rect 200757 237355 200823 237358
rect 213085 237356 213132 237358
rect 213196 237356 213202 237420
rect 230565 237418 230631 237421
rect 231669 237418 231735 237421
rect 230565 237416 231735 237418
rect 230565 237360 230570 237416
rect 230626 237360 231674 237416
rect 231730 237360 231735 237416
rect 230565 237358 231735 237360
rect 213085 237355 213151 237356
rect 230565 237355 230631 237358
rect 231669 237355 231735 237358
rect 241605 237418 241671 237421
rect 242157 237418 242223 237421
rect 241605 237416 242223 237418
rect 241605 237360 241610 237416
rect 241666 237360 242162 237416
rect 242218 237360 242223 237416
rect 241605 237358 242223 237360
rect 241605 237355 241671 237358
rect 242157 237355 242223 237358
rect 4797 237282 4863 237285
rect 136725 237282 136791 237285
rect 4797 237280 136791 237282
rect 4797 237224 4802 237280
rect 4858 237224 136730 237280
rect 136786 237224 136791 237280
rect 4797 237222 136791 237224
rect 4797 237219 4863 237222
rect 136725 237219 136791 237222
rect 149053 237282 149119 237285
rect 155166 237282 155172 237284
rect 149053 237280 155172 237282
rect 149053 237224 149058 237280
rect 149114 237224 155172 237280
rect 149053 237222 155172 237224
rect 149053 237219 149119 237222
rect 155166 237220 155172 237222
rect 155236 237220 155242 237284
rect 196934 237220 196940 237284
rect 197004 237282 197010 237284
rect 202045 237282 202111 237285
rect 197004 237280 202111 237282
rect 197004 237224 202050 237280
rect 202106 237224 202111 237280
rect 197004 237222 202111 237224
rect 197004 237220 197010 237222
rect 202045 237219 202111 237222
rect 216029 237282 216095 237285
rect 260189 237282 260255 237285
rect 216029 237280 260255 237282
rect 216029 237224 216034 237280
rect 216090 237224 260194 237280
rect 260250 237224 260255 237280
rect 216029 237222 260255 237224
rect 216029 237219 216095 237222
rect 260189 237219 260255 237222
rect 67817 237146 67883 237149
rect 162117 237146 162183 237149
rect 67817 237144 162183 237146
rect 67817 237088 67822 237144
rect 67878 237088 162122 237144
rect 162178 237088 162183 237144
rect 67817 237086 162183 237088
rect 67817 237083 67883 237086
rect 162117 237083 162183 237086
rect 186814 237084 186820 237148
rect 186884 237146 186890 237148
rect 225229 237146 225295 237149
rect 186884 237144 225295 237146
rect 186884 237088 225234 237144
rect 225290 237088 225295 237144
rect 186884 237086 225295 237088
rect 186884 237084 186890 237086
rect 225229 237083 225295 237086
rect 166257 236738 166323 236741
rect 169753 236738 169819 236741
rect 166257 236736 169819 236738
rect 166257 236680 166262 236736
rect 166318 236680 169758 236736
rect 169814 236680 169819 236736
rect 166257 236678 169819 236680
rect 166257 236675 166323 236678
rect 169753 236675 169819 236678
rect 202781 236738 202847 236741
rect 205081 236738 205147 236741
rect 202781 236736 205147 236738
rect 202781 236680 202786 236736
rect 202842 236680 205086 236736
rect 205142 236680 205147 236736
rect 202781 236678 205147 236680
rect 202781 236675 202847 236678
rect 205081 236675 205147 236678
rect 74717 236602 74783 236605
rect 238937 236602 239003 236605
rect 248597 236602 248663 236605
rect 74717 236600 248663 236602
rect 74717 236544 74722 236600
rect 74778 236544 238942 236600
rect 238998 236544 248602 236600
rect 248658 236544 248663 236600
rect 74717 236542 248663 236544
rect 74717 236539 74783 236542
rect 238937 236539 239003 236542
rect 248597 236539 248663 236542
rect 136725 236058 136791 236061
rect 137277 236058 137343 236061
rect 136725 236056 137343 236058
rect 136725 236000 136730 236056
rect 136786 236000 137282 236056
rect 137338 236000 137343 236056
rect 136725 235998 137343 236000
rect 136725 235995 136791 235998
rect 137277 235995 137343 235998
rect 176009 236058 176075 236061
rect 180149 236058 180215 236061
rect 176009 236056 180215 236058
rect 176009 236000 176014 236056
rect 176070 236000 180154 236056
rect 180210 236000 180215 236056
rect 176009 235998 180215 236000
rect 176009 235995 176075 235998
rect 180149 235995 180215 235998
rect 56409 235922 56475 235925
rect 176101 235922 176167 235925
rect 56409 235920 176167 235922
rect 56409 235864 56414 235920
rect 56470 235864 176106 235920
rect 176162 235864 176167 235920
rect 56409 235862 176167 235864
rect 56409 235859 56475 235862
rect 176101 235859 176167 235862
rect 179321 235922 179387 235925
rect 242709 235922 242775 235925
rect 179321 235920 242775 235922
rect 179321 235864 179326 235920
rect 179382 235864 242714 235920
rect 242770 235864 242775 235920
rect 179321 235862 242775 235864
rect 179321 235859 179387 235862
rect 242709 235859 242775 235862
rect 150525 235786 150591 235789
rect 180006 235786 180012 235788
rect 150525 235784 180012 235786
rect 150525 235728 150530 235784
rect 150586 235728 180012 235784
rect 150525 235726 180012 235728
rect 150525 235723 150591 235726
rect 180006 235724 180012 235726
rect 180076 235724 180082 235788
rect 188286 235724 188292 235788
rect 188356 235786 188362 235788
rect 236453 235786 236519 235789
rect 188356 235784 236519 235786
rect 188356 235728 236458 235784
rect 236514 235728 236519 235784
rect 188356 235726 236519 235728
rect 188356 235724 188362 235726
rect 236453 235723 236519 235726
rect 116025 235650 116091 235653
rect 155677 235650 155743 235653
rect 116025 235648 155743 235650
rect 116025 235592 116030 235648
rect 116086 235592 155682 235648
rect 155738 235592 155743 235648
rect 116025 235590 155743 235592
rect 116025 235587 116091 235590
rect 155677 235587 155743 235590
rect 196617 235650 196683 235653
rect 210325 235650 210391 235653
rect 196617 235648 210391 235650
rect 196617 235592 196622 235648
rect 196678 235592 210330 235648
rect 210386 235592 210391 235648
rect 196617 235590 210391 235592
rect 196617 235587 196683 235590
rect 210325 235587 210391 235590
rect 157977 235242 158043 235245
rect 158713 235242 158779 235245
rect 195278 235242 195284 235244
rect 157977 235240 195284 235242
rect 157977 235184 157982 235240
rect 158038 235184 158718 235240
rect 158774 235184 195284 235240
rect 157977 235182 195284 235184
rect 157977 235179 158043 235182
rect 158713 235179 158779 235182
rect 195278 235180 195284 235182
rect 195348 235180 195354 235244
rect 213729 234698 213795 234701
rect 214046 234698 214052 234700
rect 213729 234696 214052 234698
rect 213729 234640 213734 234696
rect 213790 234640 214052 234696
rect 213729 234638 214052 234640
rect 213729 234635 213795 234638
rect 214046 234636 214052 234638
rect 214116 234636 214122 234700
rect 59169 234562 59235 234565
rect 245878 234562 245884 234564
rect 59169 234560 245884 234562
rect 59169 234504 59174 234560
rect 59230 234504 245884 234560
rect 59169 234502 245884 234504
rect 59169 234499 59235 234502
rect 245878 234500 245884 234502
rect 245948 234500 245954 234564
rect 252502 234562 252508 234564
rect 248370 234502 252508 234562
rect 142337 234426 142403 234429
rect 163589 234426 163655 234429
rect 142337 234424 163655 234426
rect 142337 234368 142342 234424
rect 142398 234368 163594 234424
rect 163650 234368 163655 234424
rect 142337 234366 163655 234368
rect 142337 234363 142403 234366
rect 163589 234363 163655 234366
rect 191046 234364 191052 234428
rect 191116 234426 191122 234428
rect 208853 234426 208919 234429
rect 191116 234424 208919 234426
rect 191116 234368 208858 234424
rect 208914 234368 208919 234424
rect 191116 234366 208919 234368
rect 191116 234364 191122 234366
rect 208853 234363 208919 234366
rect 216581 234426 216647 234429
rect 248370 234426 248430 234502
rect 252502 234500 252508 234502
rect 252572 234562 252578 234564
rect 580257 234562 580323 234565
rect 252572 234560 580323 234562
rect 252572 234504 580262 234560
rect 580318 234504 580323 234560
rect 252572 234502 580323 234504
rect 252572 234500 252578 234502
rect 580257 234499 580323 234502
rect 216581 234424 248430 234426
rect 216581 234368 216586 234424
rect 216642 234368 248430 234424
rect 216581 234366 248430 234368
rect 216581 234363 216647 234366
rect 65926 233820 65932 233884
rect 65996 233882 66002 233884
rect 122097 233882 122163 233885
rect 65996 233880 122163 233882
rect 65996 233824 122102 233880
rect 122158 233824 122163 233880
rect 65996 233822 122163 233824
rect 65996 233820 66002 233822
rect 122097 233819 122163 233822
rect 151169 233882 151235 233885
rect 233509 233882 233575 233885
rect 151169 233880 233575 233882
rect 151169 233824 151174 233880
rect 151230 233824 233514 233880
rect 233570 233824 233575 233880
rect 151169 233822 233575 233824
rect 151169 233819 151235 233822
rect 233509 233819 233575 233822
rect 125317 233338 125383 233341
rect 140773 233338 140839 233341
rect 125317 233336 140839 233338
rect 125317 233280 125322 233336
rect 125378 233280 140778 233336
rect 140834 233280 140839 233336
rect 125317 233278 140839 233280
rect 125317 233275 125383 233278
rect 140773 233275 140839 233278
rect 103513 233202 103579 233205
rect 169109 233202 169175 233205
rect 103513 233200 169175 233202
rect 103513 233144 103518 233200
rect 103574 233144 169114 233200
rect 169170 233144 169175 233200
rect 103513 233142 169175 233144
rect 103513 233139 103579 233142
rect 169109 233139 169175 233142
rect 192477 233202 192543 233205
rect 228173 233202 228239 233205
rect 192477 233200 228239 233202
rect 192477 233144 192482 233200
rect 192538 233144 228178 233200
rect 228234 233144 228239 233200
rect 192477 233142 228239 233144
rect 192477 233139 192543 233142
rect 228173 233139 228239 233142
rect 231710 233140 231716 233204
rect 231780 233202 231786 233204
rect 233366 233202 233372 233204
rect 231780 233142 233372 233202
rect 231780 233140 231786 233142
rect 233366 233140 233372 233142
rect 233436 233140 233442 233204
rect 138657 233066 138723 233069
rect 139710 233066 139716 233068
rect 138657 233064 139716 233066
rect 138657 233008 138662 233064
rect 138718 233008 139716 233064
rect 138657 233006 139716 233008
rect 138657 233003 138723 233006
rect 139710 233004 139716 233006
rect 139780 233004 139786 233068
rect 144913 233066 144979 233069
rect 177389 233066 177455 233069
rect 144913 233064 177455 233066
rect 144913 233008 144918 233064
rect 144974 233008 177394 233064
rect 177450 233008 177455 233064
rect 144913 233006 177455 233008
rect 144913 233003 144979 233006
rect 177389 233003 177455 233006
rect 173249 232794 173315 232797
rect 221917 232794 221983 232797
rect 173249 232792 221983 232794
rect 173249 232736 173254 232792
rect 173310 232736 221922 232792
rect 221978 232736 221983 232792
rect 173249 232734 221983 232736
rect 173249 232731 173315 232734
rect 221917 232731 221983 232734
rect 64597 232658 64663 232661
rect 115197 232658 115263 232661
rect 64597 232656 115263 232658
rect 64597 232600 64602 232656
rect 64658 232600 115202 232656
rect 115258 232600 115263 232656
rect 64597 232598 115263 232600
rect 64597 232595 64663 232598
rect 115197 232595 115263 232598
rect 200849 232658 200915 232661
rect 221365 232658 221431 232661
rect 200849 232656 221431 232658
rect 200849 232600 200854 232656
rect 200910 232600 221370 232656
rect 221426 232600 221431 232656
rect 200849 232598 221431 232600
rect 200849 232595 200915 232598
rect 221365 232595 221431 232598
rect 69606 232460 69612 232524
rect 69676 232522 69682 232524
rect 151077 232522 151143 232525
rect 69676 232520 151143 232522
rect 69676 232464 151082 232520
rect 151138 232464 151143 232520
rect 69676 232462 151143 232464
rect 69676 232460 69682 232462
rect 151077 232459 151143 232462
rect 221549 232522 221615 232525
rect 242934 232522 242940 232524
rect 221549 232520 242940 232522
rect 221549 232464 221554 232520
rect 221610 232464 242940 232520
rect 221549 232462 242940 232464
rect 221549 232459 221615 232462
rect 242934 232460 242940 232462
rect 243004 232460 243010 232524
rect 582649 232386 582715 232389
rect 583520 232386 584960 232476
rect 582649 232384 584960 232386
rect 582649 232328 582654 232384
rect 582710 232328 584960 232384
rect 582649 232326 584960 232328
rect 582649 232323 582715 232326
rect 583520 232236 584960 232326
rect 198733 231978 198799 231981
rect 155910 231976 198799 231978
rect 155910 231920 198738 231976
rect 198794 231920 198799 231976
rect 155910 231918 198799 231920
rect 58985 231842 59051 231845
rect 155910 231842 155970 231918
rect 198733 231915 198799 231918
rect 58985 231840 155970 231842
rect 58985 231784 58990 231840
rect 59046 231784 155970 231840
rect 58985 231782 155970 231784
rect 58985 231779 59051 231782
rect 217174 231780 217180 231844
rect 217244 231842 217250 231844
rect 217317 231842 217383 231845
rect 217244 231840 217383 231842
rect 217244 231784 217322 231840
rect 217378 231784 217383 231840
rect 217244 231782 217383 231784
rect 217244 231780 217250 231782
rect 217317 231779 217383 231782
rect 76414 231644 76420 231708
rect 76484 231706 76490 231708
rect 102133 231706 102199 231709
rect 76484 231704 102199 231706
rect 76484 231648 102138 231704
rect 102194 231648 102199 231704
rect 76484 231646 102199 231648
rect 76484 231644 76490 231646
rect 102133 231643 102199 231646
rect 106733 231706 106799 231709
rect 133597 231706 133663 231709
rect 106733 231704 133663 231706
rect 106733 231648 106738 231704
rect 106794 231648 133602 231704
rect 133658 231648 133663 231704
rect 106733 231646 133663 231648
rect 106733 231643 106799 231646
rect 133597 231643 133663 231646
rect 140773 231570 140839 231573
rect 185945 231570 186011 231573
rect 186221 231570 186287 231573
rect 140773 231568 186287 231570
rect 140773 231512 140778 231568
rect 140834 231512 185950 231568
rect 186006 231512 186226 231568
rect 186282 231512 186287 231568
rect 140773 231510 186287 231512
rect 140773 231507 140839 231510
rect 185945 231507 186011 231510
rect 186221 231507 186287 231510
rect 133086 231372 133092 231436
rect 133156 231434 133162 231436
rect 133505 231434 133571 231437
rect 209221 231434 209287 231437
rect 133156 231432 209287 231434
rect 133156 231376 133510 231432
rect 133566 231376 209226 231432
rect 209282 231376 209287 231432
rect 133156 231374 209287 231376
rect 133156 231372 133162 231374
rect 133505 231371 133571 231374
rect 209221 231371 209287 231374
rect 180241 231298 180307 231301
rect 231485 231298 231551 231301
rect 180241 231296 231551 231298
rect 180241 231240 180246 231296
rect 180302 231240 231490 231296
rect 231546 231240 231551 231296
rect 180241 231238 231551 231240
rect 180241 231235 180307 231238
rect 231485 231235 231551 231238
rect 185945 231162 186011 231165
rect 201585 231162 201651 231165
rect 185945 231160 201651 231162
rect 185945 231104 185950 231160
rect 186006 231104 201590 231160
rect 201646 231104 201651 231160
rect 185945 231102 201651 231104
rect 185945 231099 186011 231102
rect 201585 231099 201651 231102
rect 222101 231162 222167 231165
rect 307753 231162 307819 231165
rect 222101 231160 307819 231162
rect 222101 231104 222106 231160
rect 222162 231104 307758 231160
rect 307814 231104 307819 231160
rect 222101 231102 307819 231104
rect 222101 231099 222167 231102
rect 307753 231099 307819 231102
rect 69790 230420 69796 230484
rect 69860 230482 69866 230484
rect 183001 230482 183067 230485
rect 69860 230480 183067 230482
rect 69860 230424 183006 230480
rect 183062 230424 183067 230480
rect 69860 230422 183067 230424
rect 69860 230420 69866 230422
rect 183001 230419 183067 230422
rect 129549 230346 129615 230349
rect 160001 230346 160067 230349
rect 244457 230346 244523 230349
rect 129549 230344 244523 230346
rect 129549 230288 129554 230344
rect 129610 230288 160006 230344
rect 160062 230288 244462 230344
rect 244518 230288 244523 230344
rect 129549 230286 244523 230288
rect 129549 230283 129615 230286
rect 160001 230283 160067 230286
rect 244457 230283 244523 230286
rect 67950 229740 67956 229804
rect 68020 229802 68026 229804
rect 140037 229802 140103 229805
rect 68020 229800 140103 229802
rect 68020 229744 140042 229800
rect 140098 229744 140103 229800
rect 68020 229742 140103 229744
rect 68020 229740 68026 229742
rect 140037 229739 140103 229742
rect 195881 229122 195947 229125
rect 289813 229122 289879 229125
rect 195838 229120 289879 229122
rect 195838 229064 195886 229120
rect 195942 229064 289818 229120
rect 289874 229064 289879 229120
rect 195838 229062 289879 229064
rect 195838 229059 195947 229062
rect 289813 229059 289879 229062
rect 75821 228986 75887 228989
rect 195838 228986 195898 229059
rect 75821 228984 195898 228986
rect 75821 228928 75826 228984
rect 75882 228928 195898 228984
rect 75821 228926 195898 228928
rect 75821 228923 75887 228926
rect 122097 228850 122163 228853
rect 151169 228850 151235 228853
rect 122097 228848 151235 228850
rect 122097 228792 122102 228848
rect 122158 228792 151174 228848
rect 151230 228792 151235 228848
rect 122097 228790 151235 228792
rect 122097 228787 122163 228790
rect 151169 228787 151235 228790
rect 192753 228850 192819 228853
rect 237373 228850 237439 228853
rect 192753 228848 237439 228850
rect 192753 228792 192758 228848
rect 192814 228792 237378 228848
rect 237434 228792 237439 228848
rect 192753 228790 237439 228792
rect 192753 228787 192819 228790
rect 237373 228787 237439 228790
rect 61878 228380 61884 228444
rect 61948 228442 61954 228444
rect 70485 228442 70551 228445
rect 61948 228440 70551 228442
rect 61948 228384 70490 228440
rect 70546 228384 70551 228440
rect 61948 228382 70551 228384
rect 61948 228380 61954 228382
rect 70485 228379 70551 228382
rect 191649 228442 191715 228445
rect 205081 228442 205147 228445
rect 191649 228440 205147 228442
rect 191649 228384 191654 228440
rect 191710 228384 205086 228440
rect 205142 228384 205147 228440
rect 191649 228382 205147 228384
rect 191649 228379 191715 228382
rect 205081 228379 205147 228382
rect 66161 228306 66227 228309
rect 187693 228306 187759 228309
rect 66161 228304 187759 228306
rect 66161 228248 66166 228304
rect 66222 228248 187698 228304
rect 187754 228248 187759 228304
rect 66161 228246 187759 228248
rect 66161 228243 66227 228246
rect 187693 228243 187759 228246
rect 203609 228306 203675 228309
rect 243721 228306 243787 228309
rect 203609 228304 243787 228306
rect 203609 228248 203614 228304
rect 203670 228248 243726 228304
rect 243782 228248 243787 228304
rect 203609 228246 243787 228248
rect 203609 228243 203675 228246
rect 243721 228243 243787 228246
rect -960 227884 480 228124
rect 237373 227762 237439 227765
rect 238109 227762 238175 227765
rect 237373 227760 238175 227762
rect 237373 227704 237378 227760
rect 237434 227704 238114 227760
rect 238170 227704 238175 227760
rect 237373 227702 238175 227704
rect 237373 227699 237439 227702
rect 238109 227699 238175 227702
rect 82670 227564 82676 227628
rect 82740 227626 82746 227628
rect 245694 227626 245700 227628
rect 82740 227566 245700 227626
rect 82740 227564 82746 227566
rect 245694 227564 245700 227566
rect 245764 227564 245770 227628
rect 156597 227490 156663 227493
rect 225689 227490 225755 227493
rect 156597 227488 225755 227490
rect 156597 227432 156602 227488
rect 156658 227432 225694 227488
rect 225750 227432 225755 227488
rect 156597 227430 225755 227432
rect 156597 227427 156663 227430
rect 225689 227427 225755 227430
rect 135161 227354 135227 227357
rect 166257 227354 166323 227357
rect 135161 227352 166323 227354
rect 135161 227296 135166 227352
rect 135222 227296 166262 227352
rect 166318 227296 166323 227352
rect 135161 227294 166323 227296
rect 135161 227291 135227 227294
rect 166257 227291 166323 227294
rect 108941 227218 109007 227221
rect 158161 227218 158227 227221
rect 108941 227216 158227 227218
rect 108941 227160 108946 227216
rect 109002 227160 158166 227216
rect 158222 227160 158227 227216
rect 108941 227158 158227 227160
rect 108941 227155 109007 227158
rect 158161 227155 158227 227158
rect 61837 226266 61903 226269
rect 234981 226266 235047 226269
rect 61837 226264 235047 226266
rect 61837 226208 61842 226264
rect 61898 226208 234986 226264
rect 235042 226208 235047 226264
rect 61837 226206 235047 226208
rect 61837 226203 61903 226206
rect 234981 226203 235047 226206
rect 190821 226130 190887 226133
rect 225597 226130 225663 226133
rect 190821 226128 225663 226130
rect 190821 226072 190826 226128
rect 190882 226072 225602 226128
rect 225658 226072 225663 226128
rect 190821 226070 225663 226072
rect 190821 226067 190887 226070
rect 225597 226067 225663 226070
rect 84837 225994 84903 225997
rect 152457 225994 152523 225997
rect 84837 225992 152523 225994
rect 84837 225936 84842 225992
rect 84898 225936 152462 225992
rect 152518 225936 152523 225992
rect 84837 225934 152523 225936
rect 84837 225931 84903 225934
rect 152457 225931 152523 225934
rect 69657 225858 69723 225861
rect 192661 225858 192727 225861
rect 69657 225856 192727 225858
rect 69657 225800 69662 225856
rect 69718 225800 192666 225856
rect 192722 225800 192727 225856
rect 69657 225798 192727 225800
rect 69657 225795 69723 225798
rect 192661 225795 192727 225798
rect 212165 225042 212231 225045
rect 582649 225042 582715 225045
rect 212165 225040 582715 225042
rect 212165 224984 212170 225040
rect 212226 224984 582654 225040
rect 582710 224984 582715 225040
rect 212165 224982 582715 224984
rect 212165 224979 212231 224982
rect 582649 224979 582715 224982
rect 84101 224906 84167 224909
rect 239765 224906 239831 224909
rect 84101 224904 239831 224906
rect 84101 224848 84106 224904
rect 84162 224848 239770 224904
rect 239826 224848 239831 224904
rect 84101 224846 239831 224848
rect 84101 224843 84167 224846
rect 239765 224843 239831 224846
rect 161381 224770 161447 224773
rect 232589 224770 232655 224773
rect 161381 224768 232655 224770
rect 161381 224712 161386 224768
rect 161442 224712 232594 224768
rect 232650 224712 232655 224768
rect 161381 224710 232655 224712
rect 161381 224707 161447 224710
rect 232589 224707 232655 224710
rect 137277 224634 137343 224637
rect 196709 224634 196775 224637
rect 137277 224632 196775 224634
rect 137277 224576 137282 224632
rect 137338 224576 196714 224632
rect 196770 224576 196775 224632
rect 137277 224574 196775 224576
rect 137277 224571 137343 224574
rect 196709 224571 196775 224574
rect 51717 224226 51783 224229
rect 150382 224226 150388 224228
rect 51717 224224 150388 224226
rect 51717 224168 51722 224224
rect 51778 224168 150388 224224
rect 51717 224166 150388 224168
rect 51717 224163 51783 224166
rect 150382 224164 150388 224166
rect 150452 224164 150458 224228
rect 209037 224226 209103 224229
rect 210693 224226 210759 224229
rect 285806 224226 285812 224228
rect 209037 224224 285812 224226
rect 209037 224168 209042 224224
rect 209098 224168 210698 224224
rect 210754 224168 285812 224224
rect 209037 224166 285812 224168
rect 209037 224163 209103 224166
rect 210693 224163 210759 224166
rect 285806 224164 285812 224166
rect 285876 224164 285882 224228
rect 77201 223546 77267 223549
rect 203517 223546 203583 223549
rect 77201 223544 203583 223546
rect 77201 223488 77206 223544
rect 77262 223488 203522 223544
rect 203578 223488 203583 223544
rect 77201 223486 203583 223488
rect 77201 223483 77267 223486
rect 203517 223483 203583 223486
rect 119337 223410 119403 223413
rect 189809 223410 189875 223413
rect 119337 223408 189875 223410
rect 119337 223352 119342 223408
rect 119398 223352 189814 223408
rect 189870 223352 189875 223408
rect 119337 223350 189875 223352
rect 119337 223347 119403 223350
rect 189809 223347 189875 223350
rect 191046 222940 191052 223004
rect 191116 223002 191122 223004
rect 245837 223002 245903 223005
rect 191116 223000 245903 223002
rect 191116 222944 245842 223000
rect 245898 222944 245903 223000
rect 191116 222942 245903 222944
rect 191116 222940 191122 222942
rect 245837 222939 245903 222942
rect 67265 222866 67331 222869
rect 356053 222866 356119 222869
rect 67265 222864 356119 222866
rect 67265 222808 67270 222864
rect 67326 222808 356058 222864
rect 356114 222808 356119 222864
rect 67265 222806 356119 222808
rect 67265 222803 67331 222806
rect 356053 222803 356119 222806
rect 115197 222186 115263 222189
rect 212165 222186 212231 222189
rect 115197 222184 212231 222186
rect 115197 222128 115202 222184
rect 115258 222128 212170 222184
rect 212226 222128 212231 222184
rect 115197 222126 212231 222128
rect 115197 222123 115263 222126
rect 212165 222123 212231 222126
rect 204897 222050 204963 222053
rect 205357 222050 205423 222053
rect 204897 222048 205423 222050
rect 204897 221992 204902 222048
rect 204958 221992 205362 222048
rect 205418 221992 205423 222048
rect 204897 221990 205423 221992
rect 204897 221987 204963 221990
rect 205357 221987 205423 221990
rect 101949 221506 102015 221509
rect 196617 221506 196683 221509
rect 101949 221504 196683 221506
rect 101949 221448 101954 221504
rect 102010 221448 196622 221504
rect 196678 221448 196683 221504
rect 101949 221446 196683 221448
rect 101949 221443 102015 221446
rect 196617 221443 196683 221446
rect 191925 220962 191991 220965
rect 204897 220962 204963 220965
rect 191925 220960 204963 220962
rect 191925 220904 191930 220960
rect 191986 220904 204902 220960
rect 204958 220904 204963 220960
rect 191925 220902 204963 220904
rect 191925 220899 191991 220902
rect 204897 220899 204963 220902
rect 209773 220962 209839 220965
rect 583753 220962 583819 220965
rect 209773 220960 583819 220962
rect 209773 220904 209778 220960
rect 209834 220904 583758 220960
rect 583814 220904 583819 220960
rect 209773 220902 583819 220904
rect 209773 220899 209839 220902
rect 583753 220899 583819 220902
rect 57605 220826 57671 220829
rect 184565 220826 184631 220829
rect 57605 220824 184631 220826
rect 57605 220768 57610 220824
rect 57666 220768 184570 220824
rect 184626 220768 184631 220824
rect 57605 220766 184631 220768
rect 57605 220763 57671 220766
rect 184565 220763 184631 220766
rect 187693 220826 187759 220829
rect 248689 220826 248755 220829
rect 187693 220824 248755 220826
rect 187693 220768 187698 220824
rect 187754 220768 248694 220824
rect 248750 220768 248755 220824
rect 187693 220766 248755 220768
rect 187693 220763 187759 220766
rect 248689 220763 248755 220766
rect 136541 220690 136607 220693
rect 167821 220690 167887 220693
rect 136541 220688 167887 220690
rect 136541 220632 136546 220688
rect 136602 220632 167826 220688
rect 167882 220632 167887 220688
rect 136541 220630 167887 220632
rect 136541 220627 136607 220630
rect 167821 220627 167887 220630
rect 90909 220146 90975 220149
rect 299473 220146 299539 220149
rect 90909 220144 299539 220146
rect 90909 220088 90914 220144
rect 90970 220088 299478 220144
rect 299534 220088 299539 220144
rect 90909 220086 299539 220088
rect 90909 220083 90975 220086
rect 299473 220083 299539 220086
rect 114461 219330 114527 219333
rect 209129 219330 209195 219333
rect 114461 219328 209195 219330
rect 114461 219272 114466 219328
rect 114522 219272 209134 219328
rect 209190 219272 209195 219328
rect 114461 219270 209195 219272
rect 114461 219267 114527 219270
rect 209129 219267 209195 219270
rect 155166 219132 155172 219196
rect 155236 219194 155242 219196
rect 230197 219194 230263 219197
rect 155236 219192 230263 219194
rect 155236 219136 230202 219192
rect 230258 219136 230263 219192
rect 155236 219134 230263 219136
rect 155236 219132 155242 219134
rect 230197 219131 230263 219134
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 93669 218650 93735 218653
rect 298686 218650 298692 218652
rect 93669 218648 298692 218650
rect 93669 218592 93674 218648
rect 93730 218592 298692 218648
rect 93669 218590 298692 218592
rect 93669 218587 93735 218590
rect 298686 218588 298692 218590
rect 298756 218588 298762 218652
rect 110321 217970 110387 217973
rect 219525 217970 219591 217973
rect 110321 217968 219591 217970
rect 110321 217912 110326 217968
rect 110382 217912 219530 217968
rect 219586 217912 219591 217968
rect 110321 217910 219591 217912
rect 110321 217907 110387 217910
rect 219525 217907 219591 217910
rect 86953 217834 87019 217837
rect 184289 217834 184355 217837
rect 86953 217832 184355 217834
rect 86953 217776 86958 217832
rect 87014 217776 184294 217832
rect 184350 217776 184355 217832
rect 86953 217774 184355 217776
rect 86953 217771 87019 217774
rect 184289 217771 184355 217774
rect 67173 217290 67239 217293
rect 583385 217290 583451 217293
rect 67173 217288 583451 217290
rect 67173 217232 67178 217288
rect 67234 217232 583390 217288
rect 583446 217232 583451 217288
rect 67173 217230 583451 217232
rect 67173 217227 67239 217230
rect 583385 217227 583451 217230
rect 60549 216610 60615 216613
rect 218789 216610 218855 216613
rect 60549 216608 218855 216610
rect 60549 216552 60554 216608
rect 60610 216552 218794 216608
rect 218850 216552 218855 216608
rect 60549 216550 218855 216552
rect 60549 216547 60615 216550
rect 218789 216547 218855 216550
rect 189717 216066 189783 216069
rect 206277 216066 206343 216069
rect 189717 216064 206343 216066
rect 189717 216008 189722 216064
rect 189778 216008 206282 216064
rect 206338 216008 206343 216064
rect 189717 216006 206343 216008
rect 189717 216003 189783 216006
rect 206277 216003 206343 216006
rect 92289 215930 92355 215933
rect 193949 215930 194015 215933
rect 92289 215928 194015 215930
rect 92289 215872 92294 215928
rect 92350 215872 193954 215928
rect 194010 215872 194015 215928
rect 92289 215870 194015 215872
rect 92289 215867 92355 215870
rect 193949 215867 194015 215870
rect 209630 215868 209636 215932
rect 209700 215930 209706 215932
rect 283097 215930 283163 215933
rect 209700 215928 283163 215930
rect 209700 215872 283102 215928
rect 283158 215872 283163 215928
rect 209700 215870 283163 215872
rect 209700 215868 209706 215870
rect 283097 215867 283163 215870
rect 122649 215250 122715 215253
rect 224953 215250 225019 215253
rect 122649 215248 225019 215250
rect 122649 215192 122654 215248
rect 122710 215192 224958 215248
rect 225014 215192 225019 215248
rect 122649 215190 225019 215192
rect 122649 215187 122715 215190
rect 224953 215187 225019 215190
rect -960 214978 480 215068
rect 3417 214978 3483 214981
rect -960 214976 3483 214978
rect -960 214920 3422 214976
rect 3478 214920 3483 214976
rect -960 214918 3483 214920
rect -960 214828 480 214918
rect 3417 214915 3483 214918
rect 224953 214842 225019 214845
rect 225689 214842 225755 214845
rect 224953 214840 225755 214842
rect 224953 214784 224958 214840
rect 225014 214784 225694 214840
rect 225750 214784 225755 214840
rect 224953 214782 225755 214784
rect 224953 214779 225019 214782
rect 225689 214779 225755 214782
rect 132309 214570 132375 214573
rect 186814 214570 186820 214572
rect 132309 214568 186820 214570
rect 132309 214512 132314 214568
rect 132370 214512 186820 214568
rect 132309 214510 186820 214512
rect 132309 214507 132375 214510
rect 186814 214508 186820 214510
rect 186884 214508 186890 214572
rect 194409 214570 194475 214573
rect 291377 214570 291443 214573
rect 194409 214568 291443 214570
rect 194409 214512 194414 214568
rect 194470 214512 291382 214568
rect 291438 214512 291443 214568
rect 194409 214510 291443 214512
rect 194409 214507 194475 214510
rect 291377 214507 291443 214510
rect 147673 214026 147739 214029
rect 197353 214026 197419 214029
rect 147673 214024 197419 214026
rect 147673 213968 147678 214024
rect 147734 213968 197358 214024
rect 197414 213968 197419 214024
rect 147673 213966 197419 213968
rect 147673 213963 147739 213966
rect 197353 213963 197419 213966
rect 54937 213890 55003 213893
rect 209773 213890 209839 213893
rect 54937 213888 209839 213890
rect 54937 213832 54942 213888
rect 54998 213832 209778 213888
rect 209834 213832 209839 213888
rect 54937 213830 209839 213832
rect 54937 213827 55003 213830
rect 209773 213827 209839 213830
rect 214833 213890 214899 213893
rect 215334 213890 215340 213892
rect 214833 213888 215340 213890
rect 214833 213832 214838 213888
rect 214894 213832 215340 213888
rect 214833 213830 215340 213832
rect 214833 213827 214899 213830
rect 215334 213828 215340 213830
rect 215404 213828 215410 213892
rect 126881 213754 126947 213757
rect 220261 213754 220327 213757
rect 126881 213752 220327 213754
rect 126881 213696 126886 213752
rect 126942 213696 220266 213752
rect 220322 213696 220327 213752
rect 126881 213694 220327 213696
rect 126881 213691 126947 213694
rect 220261 213691 220327 213694
rect 224718 213284 224724 213348
rect 224788 213346 224794 213348
rect 240133 213346 240199 213349
rect 224788 213344 240199 213346
rect 224788 213288 240138 213344
rect 240194 213288 240199 213344
rect 224788 213286 240199 213288
rect 224788 213284 224794 213286
rect 240133 213283 240199 213286
rect 210417 213210 210483 213213
rect 213126 213210 213132 213212
rect 210417 213208 213132 213210
rect 210417 213152 210422 213208
rect 210478 213152 213132 213208
rect 210417 213150 213132 213152
rect 210417 213147 210483 213150
rect 213126 213148 213132 213150
rect 213196 213210 213202 213212
rect 289997 213210 290063 213213
rect 213196 213208 290063 213210
rect 213196 213152 290002 213208
rect 290058 213152 290063 213208
rect 213196 213150 290063 213152
rect 213196 213148 213202 213150
rect 289997 213147 290063 213150
rect 59077 212530 59143 212533
rect 196249 212530 196315 212533
rect 59077 212528 196315 212530
rect 59077 212472 59082 212528
rect 59138 212472 196254 212528
rect 196310 212472 196315 212528
rect 59077 212470 196315 212472
rect 59077 212467 59143 212470
rect 196249 212467 196315 212470
rect 102041 212394 102107 212397
rect 172421 212394 172487 212397
rect 102041 212392 172487 212394
rect 102041 212336 102046 212392
rect 102102 212336 172426 212392
rect 172482 212336 172487 212392
rect 102041 212334 172487 212336
rect 102041 212331 102107 212334
rect 172421 212331 172487 212334
rect 172789 212394 172855 212397
rect 217041 212394 217107 212397
rect 217501 212394 217567 212397
rect 172789 212392 217567 212394
rect 172789 212336 172794 212392
rect 172850 212336 217046 212392
rect 217102 212336 217506 212392
rect 217562 212336 217567 212392
rect 172789 212334 217567 212336
rect 172789 212331 172855 212334
rect 217041 212331 217107 212334
rect 217501 212331 217567 212334
rect 206461 211986 206527 211989
rect 231894 211986 231900 211988
rect 206461 211984 231900 211986
rect 206461 211928 206466 211984
rect 206522 211928 231900 211984
rect 206461 211926 231900 211928
rect 206461 211923 206527 211926
rect 231894 211924 231900 211926
rect 231964 211924 231970 211988
rect 162209 211850 162275 211853
rect 180057 211850 180123 211853
rect 162209 211848 180123 211850
rect 162209 211792 162214 211848
rect 162270 211792 180062 211848
rect 180118 211792 180123 211848
rect 162209 211790 180123 211792
rect 162209 211787 162275 211790
rect 180057 211787 180123 211790
rect 196249 211850 196315 211853
rect 197261 211850 197327 211853
rect 209129 211850 209195 211853
rect 196249 211848 209195 211850
rect 196249 211792 196254 211848
rect 196310 211792 197266 211848
rect 197322 211792 209134 211848
rect 209190 211792 209195 211848
rect 196249 211790 209195 211792
rect 196249 211787 196315 211790
rect 197261 211787 197327 211790
rect 209129 211787 209195 211790
rect 226977 211850 227043 211853
rect 276657 211850 276723 211853
rect 226977 211848 276723 211850
rect 226977 211792 226982 211848
rect 227038 211792 276662 211848
rect 276718 211792 276723 211848
rect 226977 211790 276723 211792
rect 226977 211787 227043 211790
rect 276657 211787 276723 211790
rect 217041 211170 217107 211173
rect 220261 211170 220327 211173
rect 217041 211168 220327 211170
rect 217041 211112 217046 211168
rect 217102 211112 220266 211168
rect 220322 211112 220327 211168
rect 217041 211110 220327 211112
rect 217041 211107 217107 211110
rect 220261 211107 220327 211110
rect 128353 211034 128419 211037
rect 206369 211034 206435 211037
rect 128353 211032 206435 211034
rect 128353 210976 128358 211032
rect 128414 210976 206374 211032
rect 206430 210976 206435 211032
rect 128353 210974 206435 210976
rect 128353 210971 128419 210974
rect 206369 210971 206435 210974
rect 153101 210898 153167 210901
rect 162853 210898 162919 210901
rect 237373 210898 237439 210901
rect 153101 210896 237439 210898
rect 153101 210840 153106 210896
rect 153162 210840 162858 210896
rect 162914 210840 237378 210896
rect 237434 210840 237439 210896
rect 153101 210838 237439 210840
rect 153101 210835 153167 210838
rect 162853 210835 162919 210838
rect 237373 210835 237439 210838
rect 3417 210354 3483 210357
rect 155166 210354 155172 210356
rect 3417 210352 155172 210354
rect 3417 210296 3422 210352
rect 3478 210296 155172 210352
rect 3417 210294 155172 210296
rect 3417 210291 3483 210294
rect 155166 210292 155172 210294
rect 155236 210292 155242 210356
rect 166206 210292 166212 210356
rect 166276 210354 166282 210356
rect 345013 210354 345079 210357
rect 166276 210352 345079 210354
rect 166276 210296 345018 210352
rect 345074 210296 345079 210352
rect 166276 210294 345079 210296
rect 166276 210292 166282 210294
rect 345013 210291 345079 210294
rect 92381 209674 92447 209677
rect 211245 209674 211311 209677
rect 92381 209672 211311 209674
rect 92381 209616 92386 209672
rect 92442 209616 211250 209672
rect 211306 209616 211311 209672
rect 92381 209614 211311 209616
rect 92381 209611 92447 209614
rect 211245 209611 211311 209614
rect 85481 209130 85547 209133
rect 257337 209130 257403 209133
rect 85481 209128 257403 209130
rect 85481 209072 85486 209128
rect 85542 209072 257342 209128
rect 257398 209072 257403 209128
rect 85481 209070 257403 209072
rect 85481 209067 85547 209070
rect 257337 209067 257403 209070
rect 140681 208994 140747 208997
rect 332685 208994 332751 208997
rect 140681 208992 332751 208994
rect 140681 208936 140686 208992
rect 140742 208936 332690 208992
rect 332746 208936 332751 208992
rect 140681 208934 332751 208936
rect 140681 208931 140747 208934
rect 332685 208931 332751 208934
rect 211245 208450 211311 208453
rect 211889 208450 211955 208453
rect 211245 208448 211955 208450
rect 211245 208392 211250 208448
rect 211306 208392 211894 208448
rect 211950 208392 211955 208448
rect 211245 208390 211955 208392
rect 211245 208387 211311 208390
rect 211889 208387 211955 208390
rect 52177 208314 52243 208317
rect 218053 208314 218119 208317
rect 52177 208312 218119 208314
rect 52177 208256 52182 208312
rect 52238 208256 218058 208312
rect 218114 208256 218119 208312
rect 52177 208254 218119 208256
rect 52177 208251 52243 208254
rect 218053 208251 218119 208254
rect 133689 207770 133755 207773
rect 314009 207770 314075 207773
rect 133689 207768 314075 207770
rect 133689 207712 133694 207768
rect 133750 207712 314014 207768
rect 314070 207712 314075 207768
rect 133689 207710 314075 207712
rect 133689 207707 133755 207710
rect 314009 207707 314075 207710
rect 100661 207634 100727 207637
rect 300853 207634 300919 207637
rect 100661 207632 300919 207634
rect 100661 207576 100666 207632
rect 100722 207576 300858 207632
rect 300914 207576 300919 207632
rect 100661 207574 300919 207576
rect 100661 207571 100727 207574
rect 300853 207571 300919 207574
rect 218053 207090 218119 207093
rect 218697 207090 218763 207093
rect 218053 207088 218763 207090
rect 218053 207032 218058 207088
rect 218114 207032 218702 207088
rect 218758 207032 218763 207088
rect 218053 207030 218763 207032
rect 218053 207027 218119 207030
rect 218697 207027 218763 207030
rect 124121 206954 124187 206957
rect 240869 206954 240935 206957
rect 124121 206952 240935 206954
rect 124121 206896 124126 206952
rect 124182 206896 240874 206952
rect 240930 206896 240935 206952
rect 124121 206894 240935 206896
rect 124121 206891 124187 206894
rect 240869 206891 240935 206894
rect 66662 206212 66668 206276
rect 66732 206274 66738 206276
rect 583569 206274 583635 206277
rect 66732 206272 583635 206274
rect 66732 206216 583574 206272
rect 583630 206216 583635 206272
rect 66732 206214 583635 206216
rect 66732 206212 66738 206214
rect 583569 206211 583635 206214
rect 583109 205730 583175 205733
rect 583520 205730 584960 205820
rect 583109 205728 584960 205730
rect 583109 205672 583114 205728
rect 583170 205672 584960 205728
rect 583109 205670 584960 205672
rect 583109 205667 583175 205670
rect 67633 205594 67699 205597
rect 207381 205594 207447 205597
rect 67633 205592 209790 205594
rect 67633 205536 67638 205592
rect 67694 205536 207386 205592
rect 207442 205536 209790 205592
rect 583520 205580 584960 205670
rect 67633 205534 209790 205536
rect 67633 205531 67699 205534
rect 207381 205531 207447 205534
rect 154389 205050 154455 205053
rect 195237 205050 195303 205053
rect 154389 205048 195303 205050
rect 154389 204992 154394 205048
rect 154450 204992 195242 205048
rect 195298 204992 195303 205048
rect 154389 204990 195303 204992
rect 209730 205050 209790 205534
rect 244273 205188 244339 205189
rect 244222 205124 244228 205188
rect 244292 205186 244339 205188
rect 244292 205184 244384 205186
rect 244334 205128 244384 205184
rect 244292 205126 244384 205128
rect 244292 205124 244339 205126
rect 244273 205123 244339 205124
rect 225873 205050 225939 205053
rect 209730 205048 225939 205050
rect 209730 204992 225878 205048
rect 225934 204992 225939 205048
rect 209730 204990 225939 204992
rect 154389 204987 154455 204990
rect 195237 204987 195303 204990
rect 225873 204987 225939 204990
rect 122741 204914 122807 204917
rect 188429 204914 188495 204917
rect 122741 204912 188495 204914
rect 122741 204856 122746 204912
rect 122802 204856 188434 204912
rect 188490 204856 188495 204912
rect 122741 204854 188495 204856
rect 122741 204851 122807 204854
rect 188429 204851 188495 204854
rect 193949 204914 194015 204917
rect 340873 204914 340939 204917
rect 193949 204912 340939 204914
rect 193949 204856 193954 204912
rect 194010 204856 340878 204912
rect 340934 204856 340939 204912
rect 193949 204854 340939 204856
rect 193949 204851 194015 204854
rect 340873 204851 340939 204854
rect 73797 204234 73863 204237
rect 201493 204234 201559 204237
rect 202229 204234 202295 204237
rect 240225 204234 240291 204237
rect 240961 204234 241027 204237
rect 73797 204232 202295 204234
rect 73797 204176 73802 204232
rect 73858 204176 201498 204232
rect 201554 204176 202234 204232
rect 202290 204176 202295 204232
rect 73797 204174 202295 204176
rect 73797 204171 73863 204174
rect 201493 204171 201559 204174
rect 202229 204171 202295 204174
rect 219390 204232 241027 204234
rect 219390 204176 240230 204232
rect 240286 204176 240966 204232
rect 241022 204176 241027 204232
rect 219390 204174 241027 204176
rect 186957 204098 187023 204101
rect 219390 204098 219450 204174
rect 240225 204171 240291 204174
rect 240961 204171 241027 204174
rect 186957 204096 219450 204098
rect 186957 204040 186962 204096
rect 187018 204040 219450 204096
rect 186957 204038 219450 204040
rect 186957 204035 187023 204038
rect 36537 203690 36603 203693
rect 164969 203690 165035 203693
rect 36537 203688 165035 203690
rect 36537 203632 36542 203688
rect 36598 203632 164974 203688
rect 165030 203632 165035 203688
rect 36537 203630 165035 203632
rect 36537 203627 36603 203630
rect 164969 203627 165035 203630
rect 111609 203554 111675 203557
rect 306465 203554 306531 203557
rect 111609 203552 306531 203554
rect 111609 203496 111614 203552
rect 111670 203496 306470 203552
rect 306526 203496 306531 203552
rect 111609 203494 306531 203496
rect 111609 203491 111675 203494
rect 306465 203491 306531 203494
rect 121361 202874 121427 202877
rect 160921 202874 160987 202877
rect 121361 202872 160987 202874
rect 121361 202816 121366 202872
rect 121422 202816 160926 202872
rect 160982 202816 160987 202872
rect 121361 202814 160987 202816
rect 121361 202811 121427 202814
rect 160921 202811 160987 202814
rect 115749 202738 115815 202741
rect 138657 202738 138723 202741
rect 115749 202736 138723 202738
rect 115749 202680 115754 202736
rect 115810 202680 138662 202736
rect 138718 202680 138723 202736
rect 115749 202678 138723 202680
rect 115749 202675 115815 202678
rect 138657 202675 138723 202678
rect 198733 202466 198799 202469
rect 212717 202466 212783 202469
rect 198733 202464 212783 202466
rect 198733 202408 198738 202464
rect 198794 202408 212722 202464
rect 212778 202408 212783 202464
rect 198733 202406 212783 202408
rect 198733 202403 198799 202406
rect 212717 202403 212783 202406
rect 154481 202330 154547 202333
rect 169109 202330 169175 202333
rect 154481 202328 169175 202330
rect 154481 202272 154486 202328
rect 154542 202272 169114 202328
rect 169170 202272 169175 202328
rect 154481 202270 169175 202272
rect 154481 202267 154547 202270
rect 169109 202267 169175 202270
rect 185761 202330 185827 202333
rect 225597 202330 225663 202333
rect 185761 202328 225663 202330
rect 185761 202272 185766 202328
rect 185822 202272 225602 202328
rect 225658 202272 225663 202328
rect 185761 202270 225663 202272
rect 185761 202267 185827 202270
rect 225597 202267 225663 202270
rect 129641 202194 129707 202197
rect 288382 202194 288388 202196
rect 129641 202192 288388 202194
rect 129641 202136 129646 202192
rect 129702 202136 288388 202192
rect 129641 202134 288388 202136
rect 129641 202131 129707 202134
rect 288382 202132 288388 202134
rect 288452 202132 288458 202196
rect -960 201922 480 202012
rect 3049 201922 3115 201925
rect -960 201920 3115 201922
rect -960 201864 3054 201920
rect 3110 201864 3115 201920
rect -960 201862 3115 201864
rect -960 201772 480 201862
rect 3049 201859 3115 201862
rect 140037 201378 140103 201381
rect 276013 201378 276079 201381
rect 276749 201378 276815 201381
rect 140037 201376 276815 201378
rect 140037 201320 140042 201376
rect 140098 201320 276018 201376
rect 276074 201320 276754 201376
rect 276810 201320 276815 201376
rect 140037 201318 276815 201320
rect 140037 201315 140103 201318
rect 276013 201315 276079 201318
rect 276749 201315 276815 201318
rect 111701 200698 111767 200701
rect 253054 200698 253060 200700
rect 111701 200696 253060 200698
rect 111701 200640 111706 200696
rect 111762 200640 253060 200696
rect 111701 200638 253060 200640
rect 111701 200635 111767 200638
rect 253054 200636 253060 200638
rect 253124 200636 253130 200700
rect 75177 200018 75243 200021
rect 224401 200018 224467 200021
rect 75177 200016 224467 200018
rect 75177 199960 75182 200016
rect 75238 199960 224406 200016
rect 224462 199960 224467 200016
rect 75177 199958 224467 199960
rect 75177 199955 75243 199958
rect 224401 199955 224467 199958
rect 156689 199338 156755 199341
rect 353293 199338 353359 199341
rect 156689 199336 353359 199338
rect 156689 199280 156694 199336
rect 156750 199280 353298 199336
rect 353354 199280 353359 199336
rect 156689 199278 353359 199280
rect 156689 199275 156755 199278
rect 353293 199275 353359 199278
rect 202597 198794 202663 198797
rect 236729 198794 236795 198797
rect 202597 198792 236795 198794
rect 202597 198736 202602 198792
rect 202658 198736 236734 198792
rect 236790 198736 236795 198792
rect 202597 198734 236795 198736
rect 202597 198731 202663 198734
rect 236729 198731 236795 198734
rect 176009 198250 176075 198253
rect 196709 198250 196775 198253
rect 176009 198248 196775 198250
rect 176009 198192 176014 198248
rect 176070 198192 196714 198248
rect 196770 198192 196775 198248
rect 176009 198190 196775 198192
rect 176009 198187 176075 198190
rect 196709 198187 196775 198190
rect 133781 198114 133847 198117
rect 166257 198114 166323 198117
rect 133781 198112 166323 198114
rect 133781 198056 133786 198112
rect 133842 198056 166262 198112
rect 166318 198056 166323 198112
rect 133781 198054 166323 198056
rect 133781 198051 133847 198054
rect 166257 198051 166323 198054
rect 187601 198114 187667 198117
rect 278129 198114 278195 198117
rect 187601 198112 278195 198114
rect 187601 198056 187606 198112
rect 187662 198056 278134 198112
rect 278190 198056 278195 198112
rect 187601 198054 278195 198056
rect 187601 198051 187667 198054
rect 278129 198051 278195 198054
rect 73061 197978 73127 197981
rect 358813 197978 358879 197981
rect 73061 197976 358879 197978
rect 73061 197920 73066 197976
rect 73122 197920 358818 197976
rect 358874 197920 358879 197976
rect 73061 197918 358879 197920
rect 73061 197915 73127 197918
rect 358813 197915 358879 197918
rect 138657 197298 138723 197301
rect 221549 197298 221615 197301
rect 138657 197296 221615 197298
rect 138657 197240 138662 197296
rect 138718 197240 221554 197296
rect 221610 197240 221615 197296
rect 138657 197238 221615 197240
rect 138657 197235 138723 197238
rect 221549 197235 221615 197238
rect 182909 196754 182975 196757
rect 284385 196754 284451 196757
rect 182909 196752 284451 196754
rect 182909 196696 182914 196752
rect 182970 196696 284390 196752
rect 284446 196696 284451 196752
rect 182909 196694 284451 196696
rect 182909 196691 182975 196694
rect 284385 196691 284451 196694
rect 88241 196618 88307 196621
rect 315297 196618 315363 196621
rect 88241 196616 315363 196618
rect 88241 196560 88246 196616
rect 88302 196560 315302 196616
rect 315358 196560 315363 196616
rect 88241 196558 315363 196560
rect 88241 196555 88307 196558
rect 315297 196555 315363 196558
rect 226333 196074 226399 196077
rect 226926 196074 226932 196076
rect 226333 196072 226932 196074
rect 226333 196016 226338 196072
rect 226394 196016 226932 196072
rect 226333 196014 226932 196016
rect 226333 196011 226399 196014
rect 226926 196012 226932 196014
rect 226996 196074 227002 196076
rect 228449 196074 228515 196077
rect 226996 196072 228515 196074
rect 226996 196016 228454 196072
rect 228510 196016 228515 196072
rect 226996 196014 228515 196016
rect 226996 196012 227002 196014
rect 228449 196011 228515 196014
rect 231761 196074 231827 196077
rect 234654 196074 234660 196076
rect 231761 196072 234660 196074
rect 231761 196016 231766 196072
rect 231822 196016 234660 196072
rect 231761 196014 234660 196016
rect 231761 196011 231827 196014
rect 234654 196012 234660 196014
rect 234724 196012 234730 196076
rect 128261 195938 128327 195941
rect 160737 195938 160803 195941
rect 128261 195936 160803 195938
rect 128261 195880 128266 195936
rect 128322 195880 160742 195936
rect 160798 195880 160803 195936
rect 128261 195878 160803 195880
rect 128261 195875 128327 195878
rect 160737 195875 160803 195878
rect 202229 195394 202295 195397
rect 280286 195394 280292 195396
rect 202229 195392 280292 195394
rect 202229 195336 202234 195392
rect 202290 195336 280292 195392
rect 202229 195334 280292 195336
rect 202229 195331 202295 195334
rect 280286 195332 280292 195334
rect 280356 195332 280362 195396
rect 151721 195258 151787 195261
rect 316125 195258 316191 195261
rect 151721 195256 316191 195258
rect 151721 195200 151726 195256
rect 151782 195200 316130 195256
rect 316186 195200 316191 195256
rect 151721 195198 316191 195200
rect 151721 195195 151787 195198
rect 316125 195195 316191 195198
rect 187049 194034 187115 194037
rect 225689 194034 225755 194037
rect 187049 194032 225755 194034
rect 187049 193976 187054 194032
rect 187110 193976 225694 194032
rect 225750 193976 225755 194032
rect 187049 193974 225755 193976
rect 187049 193971 187115 193974
rect 225689 193971 225755 193974
rect 225873 194034 225939 194037
rect 296897 194034 296963 194037
rect 225873 194032 296963 194034
rect 225873 193976 225878 194032
rect 225934 193976 296902 194032
rect 296958 193976 296963 194032
rect 225873 193974 296963 193976
rect 225873 193971 225939 193974
rect 296897 193971 296963 193974
rect 107561 193898 107627 193901
rect 287094 193898 287100 193900
rect 107561 193896 287100 193898
rect 107561 193840 107566 193896
rect 107622 193840 287100 193896
rect 107561 193838 287100 193840
rect 107561 193835 107627 193838
rect 287094 193836 287100 193838
rect 287164 193836 287170 193900
rect 104157 193218 104223 193221
rect 232957 193218 233023 193221
rect 104157 193216 233023 193218
rect 104157 193160 104162 193216
rect 104218 193160 232962 193216
rect 233018 193160 233023 193216
rect 104157 193158 233023 193160
rect 104157 193155 104223 193158
rect 232957 193155 233023 193158
rect 583477 193082 583543 193085
rect 583477 193080 583586 193082
rect 583477 193024 583482 193080
rect 583538 193024 583586 193080
rect 583477 193019 583586 193024
rect 583526 192674 583586 193019
rect 583342 192628 583586 192674
rect 583342 192614 584960 192628
rect 79961 192538 80027 192541
rect 299657 192538 299723 192541
rect 79961 192536 299723 192538
rect 79961 192480 79966 192536
rect 80022 192480 299662 192536
rect 299718 192480 299723 192536
rect 79961 192478 299723 192480
rect 583342 192538 583402 192614
rect 583520 192538 584960 192614
rect 583342 192478 584960 192538
rect 79961 192475 80027 192478
rect 299657 192475 299723 192478
rect 583520 192388 584960 192478
rect 93761 191722 93827 191725
rect 171869 191722 171935 191725
rect 93761 191720 171935 191722
rect 93761 191664 93766 191720
rect 93822 191664 171874 191720
rect 171930 191664 171935 191720
rect 93761 191662 171935 191664
rect 93761 191659 93827 191662
rect 171869 191659 171935 191662
rect 181621 191178 181687 191181
rect 229686 191178 229692 191180
rect 181621 191176 229692 191178
rect 181621 191120 181626 191176
rect 181682 191120 229692 191176
rect 181621 191118 229692 191120
rect 181621 191115 181687 191118
rect 229686 191116 229692 191118
rect 229756 191116 229762 191180
rect 103421 191042 103487 191045
rect 318793 191042 318859 191045
rect 103421 191040 318859 191042
rect 103421 190984 103426 191040
rect 103482 190984 318798 191040
rect 318854 190984 318859 191040
rect 103421 190982 318859 190984
rect 103421 190979 103487 190982
rect 318793 190979 318859 190982
rect 217225 189954 217291 189957
rect 226374 189954 226380 189956
rect 217225 189952 226380 189954
rect 217225 189896 217230 189952
rect 217286 189896 226380 189952
rect 217225 189894 226380 189896
rect 217225 189891 217291 189894
rect 226374 189892 226380 189894
rect 226444 189892 226450 189956
rect 161974 189756 161980 189820
rect 162044 189818 162050 189820
rect 169753 189818 169819 189821
rect 162044 189816 169819 189818
rect 162044 189760 169758 189816
rect 169814 189760 169819 189816
rect 162044 189758 169819 189760
rect 162044 189756 162050 189758
rect 169753 189755 169819 189758
rect 190361 189818 190427 189821
rect 228214 189818 228220 189820
rect 190361 189816 228220 189818
rect 190361 189760 190366 189816
rect 190422 189760 228220 189816
rect 190361 189758 228220 189760
rect 190361 189755 190427 189758
rect 228214 189756 228220 189758
rect 228284 189756 228290 189820
rect 228357 189818 228423 189821
rect 240542 189818 240548 189820
rect 228357 189816 240548 189818
rect 228357 189760 228362 189816
rect 228418 189760 240548 189816
rect 228357 189758 240548 189760
rect 228357 189755 228423 189758
rect 240542 189756 240548 189758
rect 240612 189756 240618 189820
rect 95141 189682 95207 189685
rect 186957 189682 187023 189685
rect 95141 189680 187023 189682
rect 95141 189624 95146 189680
rect 95202 189624 186962 189680
rect 187018 189624 187023 189680
rect 95141 189622 187023 189624
rect 95141 189619 95207 189622
rect 186957 189619 187023 189622
rect 196709 189682 196775 189685
rect 284518 189682 284524 189684
rect 196709 189680 284524 189682
rect 196709 189624 196714 189680
rect 196770 189624 284524 189680
rect 196709 189622 284524 189624
rect 196709 189619 196775 189622
rect 284518 189620 284524 189622
rect 284588 189620 284594 189684
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 215937 188594 216003 188597
rect 241462 188594 241468 188596
rect 215937 188592 241468 188594
rect 215937 188536 215942 188592
rect 215998 188536 241468 188592
rect 215937 188534 241468 188536
rect 215937 188531 216003 188534
rect 241462 188532 241468 188534
rect 241532 188532 241538 188596
rect 206277 188458 206343 188461
rect 232078 188458 232084 188460
rect 206277 188456 232084 188458
rect 206277 188400 206282 188456
rect 206338 188400 232084 188456
rect 206277 188398 232084 188400
rect 206277 188395 206343 188398
rect 232078 188396 232084 188398
rect 232148 188396 232154 188460
rect 99281 188322 99347 188325
rect 303613 188322 303679 188325
rect 99281 188320 303679 188322
rect 99281 188264 99286 188320
rect 99342 188264 303618 188320
rect 303674 188264 303679 188320
rect 99281 188262 303679 188264
rect 99281 188259 99347 188262
rect 303613 188259 303679 188262
rect 241421 187778 241487 187781
rect 242433 187778 242499 187781
rect 241421 187776 242499 187778
rect 241421 187720 241426 187776
rect 241482 187720 242438 187776
rect 242494 187720 242499 187776
rect 241421 187718 242499 187720
rect 241421 187715 241487 187718
rect 242433 187715 242499 187718
rect 115841 187642 115907 187645
rect 222101 187642 222167 187645
rect 115841 187640 222167 187642
rect 115841 187584 115846 187640
rect 115902 187584 222106 187640
rect 222162 187584 222167 187640
rect 115841 187582 222167 187584
rect 115841 187579 115907 187582
rect 222101 187579 222167 187582
rect 238109 187234 238175 187237
rect 251214 187234 251220 187236
rect 238109 187232 251220 187234
rect 238109 187176 238114 187232
rect 238170 187176 251220 187232
rect 238109 187174 251220 187176
rect 238109 187171 238175 187174
rect 251214 187172 251220 187174
rect 251284 187172 251290 187236
rect 220721 187098 220787 187101
rect 244406 187098 244412 187100
rect 220721 187096 244412 187098
rect 220721 187040 220726 187096
rect 220782 187040 244412 187096
rect 220721 187038 244412 187040
rect 220721 187035 220787 187038
rect 244406 187036 244412 187038
rect 244476 187036 244482 187100
rect 203517 186962 203583 186965
rect 280245 186962 280311 186965
rect 203517 186960 280311 186962
rect 203517 186904 203522 186960
rect 203578 186904 280250 186960
rect 280306 186904 280311 186960
rect 203517 186902 280311 186904
rect 203517 186899 203583 186902
rect 280245 186899 280311 186902
rect 286317 186962 286383 186965
rect 295374 186962 295380 186964
rect 286317 186960 295380 186962
rect 286317 186904 286322 186960
rect 286378 186904 295380 186960
rect 286317 186902 295380 186904
rect 286317 186899 286383 186902
rect 295374 186900 295380 186902
rect 295444 186900 295450 186964
rect 145598 185676 145604 185740
rect 145668 185738 145674 185740
rect 177246 185738 177252 185740
rect 145668 185678 177252 185738
rect 145668 185676 145674 185678
rect 177246 185676 177252 185678
rect 177316 185676 177322 185740
rect 206870 185676 206876 185740
rect 206940 185738 206946 185740
rect 227662 185738 227668 185740
rect 206940 185678 227668 185738
rect 206940 185676 206946 185678
rect 227662 185676 227668 185678
rect 227732 185676 227738 185740
rect 228766 185676 228772 185740
rect 228836 185738 228842 185740
rect 279325 185738 279391 185741
rect 228836 185736 279391 185738
rect 228836 185680 279330 185736
rect 279386 185680 279391 185736
rect 228836 185678 279391 185680
rect 228836 185676 228842 185678
rect 279325 185675 279391 185678
rect 91001 185602 91067 185605
rect 246246 185602 246252 185604
rect 91001 185600 246252 185602
rect 91001 185544 91006 185600
rect 91062 185544 246252 185600
rect 91001 185542 246252 185544
rect 91001 185539 91067 185542
rect 246246 185540 246252 185542
rect 246316 185540 246322 185604
rect 269757 185602 269823 185605
rect 290590 185602 290596 185604
rect 269757 185600 290596 185602
rect 269757 185544 269762 185600
rect 269818 185544 290596 185600
rect 269757 185542 290596 185544
rect 269757 185539 269823 185542
rect 290590 185540 290596 185542
rect 290660 185540 290666 185604
rect 225597 184378 225663 184381
rect 285949 184378 286015 184381
rect 225597 184376 286015 184378
rect 225597 184320 225602 184376
rect 225658 184320 285954 184376
rect 286010 184320 286015 184376
rect 225597 184318 286015 184320
rect 225597 184315 225663 184318
rect 285949 184315 286015 184318
rect 67766 184180 67772 184244
rect 67836 184242 67842 184244
rect 342253 184242 342319 184245
rect 67836 184240 342319 184242
rect 67836 184184 342258 184240
rect 342314 184184 342319 184240
rect 67836 184182 342319 184184
rect 67836 184180 67842 184182
rect 342253 184179 342319 184182
rect 97901 183018 97967 183021
rect 249006 183018 249012 183020
rect 97901 183016 249012 183018
rect 97901 182960 97906 183016
rect 97962 182960 249012 183016
rect 97901 182958 249012 182960
rect 97901 182955 97967 182958
rect 249006 182956 249012 182958
rect 249076 182956 249082 183020
rect 170489 182882 170555 182885
rect 329833 182882 329899 182885
rect 170489 182880 329899 182882
rect 170489 182824 170494 182880
rect 170550 182824 329838 182880
rect 329894 182824 329899 182880
rect 170489 182822 329899 182824
rect 170489 182819 170555 182822
rect 329833 182819 329899 182822
rect 98913 182202 98979 182205
rect 178953 182202 179019 182205
rect 98913 182200 179019 182202
rect 98913 182144 98918 182200
rect 98974 182144 178958 182200
rect 179014 182144 179019 182200
rect 98913 182142 179019 182144
rect 98913 182139 98979 182142
rect 178953 182139 179019 182142
rect 218697 181658 218763 181661
rect 230422 181658 230428 181660
rect 218697 181656 230428 181658
rect 218697 181600 218702 181656
rect 218758 181600 230428 181656
rect 218697 181598 230428 181600
rect 218697 181595 218763 181598
rect 230422 181596 230428 181598
rect 230492 181596 230498 181660
rect 197997 181522 198063 181525
rect 237598 181522 237604 181524
rect 197997 181520 237604 181522
rect 197997 181464 198002 181520
rect 198058 181464 237604 181520
rect 197997 181462 237604 181464
rect 197997 181459 198063 181462
rect 237598 181460 237604 181462
rect 237668 181460 237674 181524
rect 262857 181522 262923 181525
rect 291326 181522 291332 181524
rect 262857 181520 291332 181522
rect 262857 181464 262862 181520
rect 262918 181464 291332 181520
rect 262857 181462 291332 181464
rect 262857 181459 262923 181462
rect 291326 181460 291332 181462
rect 291396 181460 291402 181524
rect 160829 181386 160895 181389
rect 285622 181386 285628 181388
rect 160829 181384 285628 181386
rect 160829 181328 160834 181384
rect 160890 181328 285628 181384
rect 160829 181326 285628 181328
rect 160829 181323 160895 181326
rect 285622 181324 285628 181326
rect 285692 181324 285698 181388
rect 124949 180978 125015 180981
rect 167821 180978 167887 180981
rect 124949 180976 167887 180978
rect 124949 180920 124954 180976
rect 125010 180920 167826 180976
rect 167882 180920 167887 180976
rect 124949 180918 167887 180920
rect 124949 180915 125015 180918
rect 167821 180915 167887 180918
rect 118509 180842 118575 180845
rect 170489 180842 170555 180845
rect 118509 180840 170555 180842
rect 118509 180784 118514 180840
rect 118570 180784 170494 180840
rect 170550 180784 170555 180840
rect 118509 180782 170555 180784
rect 118509 180779 118575 180782
rect 170489 180779 170555 180782
rect 225689 180162 225755 180165
rect 233417 180162 233483 180165
rect 225689 180160 233483 180162
rect 225689 180104 225694 180160
rect 225750 180104 233422 180160
rect 233478 180104 233483 180160
rect 225689 180102 233483 180104
rect 225689 180099 225755 180102
rect 233417 180099 233483 180102
rect 177941 180026 178007 180029
rect 280337 180026 280403 180029
rect 177941 180024 280403 180026
rect 177941 179968 177946 180024
rect 178002 179968 280342 180024
rect 280398 179968 280403 180024
rect 177941 179966 280403 179968
rect 177941 179963 178007 179966
rect 280337 179963 280403 179966
rect 282177 180026 282243 180029
rect 290089 180026 290155 180029
rect 282177 180024 290155 180026
rect 282177 179968 282182 180024
rect 282238 179968 290094 180024
rect 290150 179968 290155 180024
rect 282177 179966 290155 179968
rect 282177 179963 282243 179966
rect 290089 179963 290155 179966
rect 113357 179618 113423 179621
rect 169201 179618 169267 179621
rect 113357 179616 169267 179618
rect 113357 179560 113362 179616
rect 113418 179560 169206 179616
rect 169262 179560 169267 179616
rect 113357 179558 169267 179560
rect 113357 179555 113423 179558
rect 169201 179555 169267 179558
rect 100753 179482 100819 179485
rect 166349 179482 166415 179485
rect 100753 179480 166415 179482
rect 100753 179424 100758 179480
rect 100814 179424 166354 179480
rect 166410 179424 166415 179480
rect 100753 179422 166415 179424
rect 100753 179419 100819 179422
rect 166349 179419 166415 179422
rect 220261 179482 220327 179485
rect 245837 179482 245903 179485
rect 220261 179480 245903 179482
rect 220261 179424 220266 179480
rect 220322 179424 245842 179480
rect 245898 179424 245903 179480
rect 220261 179422 245903 179424
rect 220261 179419 220327 179422
rect 245837 179419 245903 179422
rect 266353 179482 266419 179485
rect 267089 179482 267155 179485
rect 281625 179482 281691 179485
rect 266353 179480 281691 179482
rect 266353 179424 266358 179480
rect 266414 179424 267094 179480
rect 267150 179424 281630 179480
rect 281686 179424 281691 179480
rect 266353 179422 281691 179424
rect 266353 179419 266419 179422
rect 267089 179419 267155 179422
rect 281625 179419 281691 179422
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 583520 179060 584960 179150
rect 185577 178938 185643 178941
rect 200757 178938 200823 178941
rect 185577 178936 200823 178938
rect 185577 178880 185582 178936
rect 185638 178880 200762 178936
rect 200818 178880 200823 178936
rect 185577 178878 200823 178880
rect 185577 178875 185643 178878
rect 200757 178875 200823 178878
rect 274541 178938 274607 178941
rect 280429 178938 280495 178941
rect 274541 178936 280495 178938
rect 274541 178880 274546 178936
rect 274602 178880 280434 178936
rect 280490 178880 280495 178936
rect 274541 178878 280495 178880
rect 274541 178875 274607 178878
rect 280429 178875 280495 178878
rect 199510 178740 199516 178804
rect 199580 178802 199586 178804
rect 236177 178802 236243 178805
rect 199580 178800 236243 178802
rect 199580 178744 236182 178800
rect 236238 178744 236243 178800
rect 199580 178742 236243 178744
rect 199580 178740 199586 178742
rect 236177 178739 236243 178742
rect 273897 178802 273963 178805
rect 291469 178802 291535 178805
rect 273897 178800 291535 178802
rect 273897 178744 273902 178800
rect 273958 178744 291474 178800
rect 291530 178744 291535 178800
rect 273897 178742 291535 178744
rect 273897 178739 273963 178742
rect 291469 178739 291535 178742
rect 198089 178666 198155 178669
rect 278814 178666 278820 178668
rect 198089 178664 278820 178666
rect 198089 178608 198094 178664
rect 198150 178608 278820 178664
rect 198089 178606 278820 178608
rect 198089 178603 198155 178606
rect 278814 178604 278820 178606
rect 278884 178604 278890 178668
rect 109534 178332 109540 178396
rect 109604 178394 109610 178396
rect 173249 178394 173315 178397
rect 109604 178392 173315 178394
rect 109604 178336 173254 178392
rect 173310 178336 173315 178392
rect 109604 178334 173315 178336
rect 109604 178332 109610 178334
rect 173249 178331 173315 178334
rect 110638 178196 110644 178260
rect 110708 178258 110714 178260
rect 177389 178258 177455 178261
rect 110708 178256 177455 178258
rect 110708 178200 177394 178256
rect 177450 178200 177455 178256
rect 110708 178198 177455 178200
rect 110708 178196 110714 178198
rect 177389 178195 177455 178198
rect 185761 178122 185827 178125
rect 97030 178120 185827 178122
rect 97030 178064 185766 178120
rect 185822 178064 185827 178120
rect 97030 178062 185827 178064
rect 97030 177988 97090 178062
rect 185761 178059 185827 178062
rect 97022 177924 97028 177988
rect 97092 177924 97098 177988
rect 197353 177986 197419 177989
rect 266353 177986 266419 177989
rect 197353 177984 266419 177986
rect 197353 177928 197358 177984
rect 197414 177928 266358 177984
rect 266414 177928 266419 177984
rect 197353 177926 266419 177928
rect 197353 177923 197419 177926
rect 266353 177923 266419 177926
rect 98310 177516 98316 177580
rect 98380 177578 98386 177580
rect 98913 177578 98979 177581
rect 102041 177580 102107 177581
rect 101990 177578 101996 177580
rect 98380 177576 98979 177578
rect 98380 177520 98918 177576
rect 98974 177520 98979 177576
rect 98380 177518 98979 177520
rect 101950 177518 101996 177578
rect 102060 177576 102107 177580
rect 102102 177520 102107 177576
rect 98380 177516 98386 177518
rect 98913 177515 98979 177518
rect 101990 177516 101996 177518
rect 102060 177516 102107 177520
rect 105670 177516 105676 177580
rect 105740 177578 105746 177580
rect 106181 177578 106247 177581
rect 105740 177576 106247 177578
rect 105740 177520 106186 177576
rect 106242 177520 106247 177576
rect 105740 177518 106247 177520
rect 105740 177516 105746 177518
rect 102041 177515 102107 177516
rect 106181 177515 106247 177518
rect 108062 177516 108068 177580
rect 108132 177578 108138 177580
rect 108941 177578 109007 177581
rect 108132 177576 109007 177578
rect 108132 177520 108946 177576
rect 109002 177520 109007 177576
rect 108132 177518 109007 177520
rect 108132 177516 108138 177518
rect 108941 177515 109007 177518
rect 112110 177516 112116 177580
rect 112180 177578 112186 177580
rect 113081 177578 113147 177581
rect 112180 177576 113147 177578
rect 112180 177520 113086 177576
rect 113142 177520 113147 177576
rect 112180 177518 113147 177520
rect 112180 177516 112186 177518
rect 113081 177515 113147 177518
rect 120758 177516 120764 177580
rect 120828 177578 120834 177580
rect 121361 177578 121427 177581
rect 120828 177576 121427 177578
rect 120828 177520 121366 177576
rect 121422 177520 121427 177576
rect 120828 177518 121427 177520
rect 120828 177516 120834 177518
rect 121361 177515 121427 177518
rect 124438 177516 124444 177580
rect 124508 177578 124514 177580
rect 124949 177578 125015 177581
rect 124508 177576 125015 177578
rect 124508 177520 124954 177576
rect 125010 177520 125015 177576
rect 124508 177518 125015 177520
rect 124508 177516 124514 177518
rect 124949 177515 125015 177518
rect 125726 177516 125732 177580
rect 125796 177578 125802 177580
rect 125961 177578 126027 177581
rect 125796 177576 126027 177578
rect 125796 177520 125966 177576
rect 126022 177520 126027 177576
rect 125796 177518 126027 177520
rect 125796 177516 125802 177518
rect 125961 177515 126027 177518
rect 127014 177516 127020 177580
rect 127084 177578 127090 177580
rect 128261 177578 128327 177581
rect 132401 177580 132467 177581
rect 132350 177578 132356 177580
rect 127084 177576 128327 177578
rect 127084 177520 128266 177576
rect 128322 177520 128327 177576
rect 127084 177518 128327 177520
rect 132310 177518 132356 177578
rect 132420 177576 132467 177580
rect 132462 177520 132467 177576
rect 127084 177516 127090 177518
rect 128261 177515 128327 177518
rect 132350 177516 132356 177518
rect 132420 177516 132467 177520
rect 133086 177516 133092 177580
rect 133156 177578 133162 177580
rect 133781 177578 133847 177581
rect 148225 177580 148291 177581
rect 148174 177578 148180 177580
rect 133156 177576 133847 177578
rect 133156 177520 133786 177576
rect 133842 177520 133847 177576
rect 133156 177518 133847 177520
rect 148134 177518 148180 177578
rect 148244 177576 148291 177580
rect 148286 177520 148291 177576
rect 133156 177516 133162 177518
rect 132401 177515 132467 177516
rect 133781 177515 133847 177518
rect 148174 177516 148180 177518
rect 148244 177516 148291 177520
rect 148225 177515 148291 177516
rect 118366 177380 118372 177444
rect 118436 177442 118442 177444
rect 118509 177442 118575 177445
rect 118436 177440 118575 177442
rect 118436 177384 118514 177440
rect 118570 177384 118575 177440
rect 118436 177382 118575 177384
rect 118436 177380 118442 177382
rect 118509 177379 118575 177382
rect 217317 177442 217383 177445
rect 227713 177442 227779 177445
rect 217317 177440 227779 177442
rect 217317 177384 217322 177440
rect 217378 177384 227718 177440
rect 227774 177384 227779 177440
rect 217317 177382 227779 177384
rect 217317 177379 217383 177382
rect 227713 177379 227779 177382
rect 276749 177442 276815 177445
rect 283782 177442 283788 177444
rect 276749 177440 283788 177442
rect 276749 177384 276754 177440
rect 276810 177384 283788 177440
rect 276749 177382 283788 177384
rect 276749 177379 276815 177382
rect 283782 177380 283788 177382
rect 283852 177380 283858 177444
rect 130694 177244 130700 177308
rect 130764 177306 130770 177308
rect 131021 177306 131087 177309
rect 130764 177304 131087 177306
rect 130764 177248 131026 177304
rect 131082 177248 131087 177304
rect 130764 177246 131087 177248
rect 130764 177244 130770 177246
rect 131021 177243 131087 177246
rect 185669 177306 185735 177309
rect 224953 177306 225019 177309
rect 185669 177304 225019 177306
rect 185669 177248 185674 177304
rect 185730 177248 224958 177304
rect 225014 177248 225019 177304
rect 185669 177246 225019 177248
rect 185669 177243 185735 177246
rect 224953 177243 225019 177246
rect 226977 177306 227043 177309
rect 234797 177306 234863 177309
rect 226977 177304 234863 177306
rect 226977 177248 226982 177304
rect 227038 177248 234802 177304
rect 234858 177248 234863 177304
rect 226977 177246 234863 177248
rect 226977 177243 227043 177246
rect 234797 177243 234863 177246
rect 278129 177306 278195 177309
rect 288709 177306 288775 177309
rect 278129 177304 288775 177306
rect 278129 177248 278134 177304
rect 278190 177248 288714 177304
rect 288770 177248 288775 177304
rect 278129 177246 288775 177248
rect 278129 177243 278195 177246
rect 288709 177243 288775 177246
rect 104566 177108 104572 177172
rect 104636 177170 104642 177172
rect 198089 177170 198155 177173
rect 104636 177168 198155 177170
rect 104636 177112 198094 177168
rect 198150 177112 198155 177168
rect 104636 177110 198155 177112
rect 104636 177108 104642 177110
rect 198089 177107 198155 177110
rect 113214 176972 113220 177036
rect 113284 177034 113290 177036
rect 113357 177034 113423 177037
rect 115841 177036 115907 177037
rect 115790 177034 115796 177036
rect 113284 177032 113423 177034
rect 113284 176976 113362 177032
rect 113418 176976 113423 177032
rect 113284 176974 113423 176976
rect 115750 176974 115796 177034
rect 115860 177032 115907 177036
rect 115902 176976 115907 177032
rect 113284 176972 113290 176974
rect 113357 176971 113423 176974
rect 115790 176972 115796 176974
rect 115860 176972 115907 176976
rect 115841 176971 115907 176972
rect 117957 177034 118023 177037
rect 169017 177034 169083 177037
rect 117957 177032 169083 177034
rect 117957 176976 117962 177032
rect 118018 176976 169022 177032
rect 169078 176976 169083 177032
rect 117957 176974 169083 176976
rect 117957 176971 118023 176974
rect 169017 176971 169083 176974
rect 278865 177034 278931 177037
rect 279366 177034 279372 177036
rect 278865 177032 279372 177034
rect 278865 176976 278870 177032
rect 278926 176976 279372 177032
rect 278865 176974 279372 176976
rect 278865 176971 278931 176974
rect 279366 176972 279372 176974
rect 279436 176972 279442 177036
rect 100753 176900 100819 176901
rect 100702 176898 100708 176900
rect 100662 176838 100708 176898
rect 100772 176896 100819 176900
rect 181529 176898 181595 176901
rect 100814 176840 100819 176896
rect 100702 176836 100708 176838
rect 100772 176836 100819 176840
rect 100753 176835 100819 176836
rect 103470 176896 181595 176898
rect 103470 176840 181534 176896
rect 181590 176840 181595 176896
rect 103470 176838 181595 176840
rect 100661 176762 100727 176765
rect 103470 176762 103530 176838
rect 181529 176835 181595 176838
rect 99422 176760 100727 176762
rect 99422 176704 100666 176760
rect 100722 176704 100727 176760
rect 99422 176702 100727 176704
rect 99422 176492 99482 176702
rect 100661 176699 100727 176702
rect 103286 176702 103530 176762
rect 103286 176492 103346 176702
rect 106958 176700 106964 176764
rect 107028 176762 107034 176764
rect 117957 176762 118023 176765
rect 121913 176764 121979 176765
rect 121862 176762 121868 176764
rect 107028 176760 118023 176762
rect 107028 176704 117962 176760
rect 118018 176704 118023 176760
rect 107028 176702 118023 176704
rect 121822 176702 121868 176762
rect 121932 176760 121979 176764
rect 121974 176704 121979 176760
rect 107028 176700 107034 176702
rect 117957 176699 118023 176702
rect 121862 176700 121868 176702
rect 121932 176700 121979 176704
rect 123150 176700 123156 176764
rect 123220 176762 123226 176764
rect 123293 176762 123359 176765
rect 128169 176762 128235 176765
rect 129457 176764 129523 176765
rect 136081 176764 136147 176765
rect 129406 176762 129412 176764
rect 123220 176760 123359 176762
rect 123220 176704 123298 176760
rect 123354 176704 123359 176760
rect 123220 176702 123359 176704
rect 123220 176700 123226 176702
rect 121913 176699 121979 176700
rect 123293 176699 123359 176702
rect 128126 176760 128235 176762
rect 128126 176704 128174 176760
rect 128230 176704 128235 176760
rect 128126 176699 128235 176704
rect 129366 176702 129412 176762
rect 129476 176760 129523 176764
rect 136030 176762 136036 176764
rect 129518 176704 129523 176760
rect 129406 176700 129412 176702
rect 129476 176700 129523 176704
rect 135990 176702 136036 176762
rect 136100 176760 136147 176764
rect 136142 176704 136147 176760
rect 136030 176700 136036 176702
rect 136100 176700 136147 176704
rect 158846 176700 158852 176764
rect 158916 176762 158922 176764
rect 158989 176762 159055 176765
rect 158916 176760 159055 176762
rect 158916 176704 158994 176760
rect 159050 176704 159055 176760
rect 158916 176702 159055 176704
rect 158916 176700 158922 176702
rect 129457 176699 129523 176700
rect 136081 176699 136147 176700
rect 158989 176699 159055 176702
rect 229318 176700 229324 176764
rect 229388 176762 229394 176764
rect 229737 176762 229803 176765
rect 229388 176760 229803 176762
rect 229388 176704 229742 176760
rect 229798 176704 229803 176760
rect 229388 176702 229803 176704
rect 229388 176700 229394 176702
rect 229737 176699 229803 176702
rect 128126 176492 128186 176699
rect 163497 176626 163563 176629
rect 220261 176626 220327 176629
rect 163497 176624 220327 176626
rect 163497 176568 163502 176624
rect 163558 176568 220266 176624
rect 220322 176568 220327 176624
rect 163497 176566 220327 176568
rect 163497 176563 163563 176566
rect 220261 176563 220327 176566
rect 222929 176626 222995 176629
rect 230606 176626 230612 176628
rect 222929 176624 230612 176626
rect 222929 176568 222934 176624
rect 222990 176568 230612 176624
rect 222929 176566 230612 176568
rect 222929 176563 222995 176566
rect 230606 176564 230612 176566
rect 230676 176564 230682 176628
rect 99414 176428 99420 176492
rect 99484 176428 99490 176492
rect 103278 176428 103284 176492
rect 103348 176428 103354 176492
rect 128118 176428 128124 176492
rect 128188 176428 128194 176492
rect 227713 176218 227779 176221
rect 227713 176216 228282 176218
rect 227713 176160 227718 176216
rect 227774 176160 228282 176216
rect 227713 176158 228282 176160
rect 227713 176155 227779 176158
rect -960 175796 480 176036
rect 166993 175948 167059 175949
rect 166942 175884 166948 175948
rect 167012 175946 167059 175948
rect 167012 175944 167104 175946
rect 167054 175888 167104 175944
rect 167012 175886 167104 175888
rect 167012 175884 167059 175886
rect 166993 175883 167059 175884
rect 213913 175674 213979 175677
rect 213913 175672 217028 175674
rect 213913 175616 213918 175672
rect 213974 175616 217028 175672
rect 228222 175644 228282 176158
rect 228449 176082 228515 176085
rect 233509 176082 233575 176085
rect 228449 176080 233575 176082
rect 228449 176024 228454 176080
rect 228510 176024 233514 176080
rect 233570 176024 233575 176080
rect 228449 176022 233575 176024
rect 228449 176019 228515 176022
rect 233509 176019 233575 176022
rect 236637 176082 236703 176085
rect 241646 176082 241652 176084
rect 236637 176080 241652 176082
rect 236637 176024 236642 176080
rect 236698 176024 241652 176080
rect 236637 176022 241652 176024
rect 236637 176019 236703 176022
rect 241646 176020 241652 176022
rect 241716 176020 241722 176084
rect 244457 176082 244523 176085
rect 241838 176080 244523 176082
rect 241838 176024 244462 176080
rect 244518 176024 244523 176080
rect 241838 176022 244523 176024
rect 231761 175946 231827 175949
rect 241838 175946 241898 176022
rect 244457 176019 244523 176022
rect 231761 175944 241898 175946
rect 231761 175888 231766 175944
rect 231822 175888 241898 175944
rect 231761 175886 241898 175888
rect 243721 175946 243787 175949
rect 247217 175946 247283 175949
rect 273345 175948 273411 175949
rect 273294 175946 273300 175948
rect 243721 175944 247283 175946
rect 243721 175888 243726 175944
rect 243782 175888 247222 175944
rect 247278 175888 247283 175944
rect 243721 175886 247283 175888
rect 273254 175886 273300 175946
rect 273364 175944 273411 175948
rect 273406 175888 273411 175944
rect 231761 175883 231827 175886
rect 243721 175883 243787 175886
rect 247217 175883 247283 175886
rect 273294 175884 273300 175886
rect 273364 175884 273411 175888
rect 273345 175883 273411 175884
rect 278773 175946 278839 175949
rect 278773 175944 279434 175946
rect 278773 175888 278778 175944
rect 278834 175888 279434 175944
rect 278773 175886 279434 175888
rect 278773 175883 278839 175886
rect 264973 175674 265039 175677
rect 264973 175672 268180 175674
rect 213913 175614 217028 175616
rect 264973 175616 264978 175672
rect 265034 175616 268180 175672
rect 264973 175614 268180 175616
rect 213913 175611 213979 175614
rect 264973 175611 265039 175614
rect 114318 175476 114324 175540
rect 114388 175538 114394 175540
rect 166533 175538 166599 175541
rect 114388 175536 166599 175538
rect 114388 175480 166538 175536
rect 166594 175480 166599 175536
rect 279374 175508 279434 175886
rect 114388 175478 166599 175480
rect 114388 175476 114394 175478
rect 166533 175475 166599 175478
rect 116894 175340 116900 175404
rect 116964 175402 116970 175404
rect 207749 175402 207815 175405
rect 116964 175400 207815 175402
rect 116964 175344 207754 175400
rect 207810 175344 207815 175400
rect 116964 175342 207815 175344
rect 116964 175340 116970 175342
rect 207749 175339 207815 175342
rect 187141 175266 187207 175269
rect 214557 175266 214623 175269
rect 231761 175266 231827 175269
rect 187141 175264 214623 175266
rect 187141 175208 187146 175264
rect 187202 175208 214562 175264
rect 214618 175208 214623 175264
rect 187141 175206 214623 175208
rect 228988 175264 231827 175266
rect 228988 175208 231766 175264
rect 231822 175208 231827 175264
rect 228988 175206 231827 175208
rect 187141 175203 187207 175206
rect 214557 175203 214623 175206
rect 231761 175203 231827 175206
rect 265065 175266 265131 175269
rect 265065 175264 268180 175266
rect 265065 175208 265070 175264
rect 265126 175208 268180 175264
rect 265065 175206 268180 175208
rect 265065 175203 265131 175206
rect 229093 175132 229159 175133
rect 229093 175128 229140 175132
rect 229204 175130 229210 175132
rect 229093 175072 229098 175128
rect 229093 175068 229140 175072
rect 229204 175070 229250 175130
rect 229204 175068 229210 175070
rect 229686 175068 229692 175132
rect 229756 175130 229762 175132
rect 232037 175130 232103 175133
rect 229756 175128 232103 175130
rect 229756 175072 232042 175128
rect 232098 175072 232103 175128
rect 229756 175070 232103 175072
rect 229756 175068 229762 175070
rect 229093 175067 229159 175068
rect 232037 175067 232103 175070
rect 119429 174996 119495 174997
rect 119392 174994 119398 174996
rect 119338 174934 119398 174994
rect 119462 174992 119495 174996
rect 119490 174936 119495 174992
rect 119392 174932 119398 174934
rect 119462 174932 119495 174936
rect 119429 174931 119495 174932
rect 213913 174994 213979 174997
rect 229277 174994 229343 174997
rect 229502 174994 229508 174996
rect 213913 174992 217028 174994
rect 213913 174936 213918 174992
rect 213974 174936 217028 174992
rect 213913 174934 217028 174936
rect 229277 174992 229508 174994
rect 229277 174936 229282 174992
rect 229338 174936 229508 174992
rect 229277 174934 229508 174936
rect 213913 174931 213979 174934
rect 229277 174931 229343 174934
rect 229502 174932 229508 174934
rect 229572 174932 229578 174996
rect 134352 174796 134358 174860
rect 134422 174858 134428 174860
rect 135253 174858 135319 174861
rect 134422 174856 135319 174858
rect 134422 174800 135258 174856
rect 135314 174800 135319 174856
rect 134422 174798 135319 174800
rect 134422 174796 134428 174798
rect 135253 174795 135319 174798
rect 264973 174858 265039 174861
rect 264973 174856 268180 174858
rect 264973 174800 264978 174856
rect 265034 174800 268180 174856
rect 264973 174798 268180 174800
rect 264973 174795 265039 174798
rect 231117 174722 231183 174725
rect 280337 174722 280403 174725
rect 228988 174720 231183 174722
rect 228988 174664 231122 174720
rect 231178 174664 231183 174720
rect 228988 174662 231183 174664
rect 279956 174720 280403 174722
rect 279956 174664 280342 174720
rect 280398 174664 280403 174720
rect 279956 174662 280403 174664
rect 231117 174659 231183 174662
rect 280337 174659 280403 174662
rect 279417 174450 279483 174453
rect 258030 174390 268180 174450
rect 279374 174448 279483 174450
rect 279374 174392 279422 174448
rect 279478 174392 279483 174448
rect 214005 174314 214071 174317
rect 229134 174314 229140 174316
rect 214005 174312 217028 174314
rect 214005 174256 214010 174312
rect 214066 174256 217028 174312
rect 214005 174254 217028 174256
rect 228988 174254 229140 174314
rect 214005 174251 214071 174254
rect 229134 174252 229140 174254
rect 229204 174252 229210 174316
rect 256141 174314 256207 174317
rect 258030 174314 258090 174390
rect 256141 174312 258090 174314
rect 256141 174256 256146 174312
rect 256202 174256 258090 174312
rect 256141 174254 258090 174256
rect 279374 174387 279483 174392
rect 256141 174251 256207 174254
rect 249149 174042 249215 174045
rect 249149 174040 268180 174042
rect 249149 173984 249154 174040
rect 249210 173984 268180 174040
rect 279374 174012 279434 174387
rect 249149 173982 268180 173984
rect 249149 173979 249215 173982
rect 239029 173906 239095 173909
rect 240358 173906 240364 173908
rect 239029 173904 240364 173906
rect 239029 173848 239034 173904
rect 239090 173848 240364 173904
rect 239029 173846 240364 173848
rect 239029 173843 239095 173846
rect 240358 173844 240364 173846
rect 240428 173844 240434 173908
rect 229093 173770 229159 173773
rect 228988 173768 229159 173770
rect 228988 173712 229098 173768
rect 229154 173712 229159 173768
rect 228988 173710 229159 173712
rect 229093 173707 229159 173710
rect 279366 173708 279372 173772
rect 279436 173708 279442 173772
rect 213913 173634 213979 173637
rect 265065 173634 265131 173637
rect 213913 173632 217028 173634
rect 213913 173576 213918 173632
rect 213974 173576 217028 173632
rect 213913 173574 217028 173576
rect 265065 173632 268180 173634
rect 265065 173576 265070 173632
rect 265126 173576 268180 173632
rect 265065 173574 268180 173576
rect 213913 173571 213979 173574
rect 265065 173571 265131 173574
rect 238518 173362 238524 173364
rect 228988 173302 238524 173362
rect 238518 173300 238524 173302
rect 238588 173300 238594 173364
rect 231761 173226 231827 173229
rect 251357 173226 251423 173229
rect 231761 173224 251423 173226
rect 231761 173168 231766 173224
rect 231822 173168 251362 173224
rect 251418 173168 251423 173224
rect 279374 173196 279434 173708
rect 231761 173166 251423 173168
rect 231761 173163 231827 173166
rect 251357 173163 251423 173166
rect 214005 172954 214071 172957
rect 214005 172952 217028 172954
rect 214005 172896 214010 172952
rect 214066 172896 217028 172952
rect 214005 172894 217028 172896
rect 214005 172891 214071 172894
rect 231577 172818 231643 172821
rect 228988 172816 231643 172818
rect 228988 172760 231582 172816
rect 231638 172760 231643 172816
rect 228988 172758 231643 172760
rect 231577 172755 231643 172758
rect 240869 172818 240935 172821
rect 268150 172818 268210 173060
rect 240869 172816 268210 172818
rect 240869 172760 240874 172816
rect 240930 172760 268210 172816
rect 240869 172758 268210 172760
rect 240869 172755 240935 172758
rect 264973 172682 265039 172685
rect 264973 172680 268180 172682
rect 264973 172624 264978 172680
rect 265034 172624 268180 172680
rect 264973 172622 268180 172624
rect 264973 172619 265039 172622
rect 282453 172546 282519 172549
rect 279956 172544 282519 172546
rect 279956 172488 282458 172544
rect 282514 172488 282519 172544
rect 279956 172486 282519 172488
rect 282453 172483 282519 172486
rect 228988 172350 238770 172410
rect 213913 172274 213979 172277
rect 238710 172274 238770 172350
rect 240358 172348 240364 172412
rect 240428 172410 240434 172412
rect 241421 172410 241487 172413
rect 240428 172408 241487 172410
rect 240428 172352 241426 172408
rect 241482 172352 241487 172408
rect 240428 172350 241487 172352
rect 240428 172348 240434 172350
rect 241421 172347 241487 172350
rect 244273 172274 244339 172277
rect 213913 172272 217028 172274
rect 213913 172216 213918 172272
rect 213974 172216 217028 172272
rect 213913 172214 217028 172216
rect 238710 172272 244339 172274
rect 238710 172216 244278 172272
rect 244334 172216 244339 172272
rect 238710 172214 244339 172216
rect 213913 172211 213979 172214
rect 244273 172211 244339 172214
rect 265065 172274 265131 172277
rect 265065 172272 268180 172274
rect 265065 172216 265070 172272
rect 265126 172216 268180 172272
rect 265065 172214 268180 172216
rect 265065 172211 265131 172214
rect 231761 171866 231827 171869
rect 228988 171864 231827 171866
rect 228988 171808 231766 171864
rect 231822 171808 231827 171864
rect 228988 171806 231827 171808
rect 231761 171803 231827 171806
rect 164724 171594 165354 171600
rect 167637 171594 167703 171597
rect 164724 171592 167703 171594
rect 164724 171540 167642 171592
rect 165294 171536 167642 171540
rect 167698 171536 167703 171592
rect 165294 171534 167703 171536
rect 167637 171531 167703 171534
rect 214097 171594 214163 171597
rect 244917 171594 244983 171597
rect 268150 171594 268210 171836
rect 282085 171730 282151 171733
rect 279956 171728 282151 171730
rect 279956 171672 282090 171728
rect 282146 171672 282151 171728
rect 279956 171670 282151 171672
rect 282085 171667 282151 171670
rect 214097 171592 217028 171594
rect 214097 171536 214102 171592
rect 214158 171536 217028 171592
rect 214097 171534 217028 171536
rect 244917 171592 268210 171594
rect 244917 171536 244922 171592
rect 244978 171536 268210 171592
rect 244917 171534 268210 171536
rect 214097 171531 214163 171534
rect 244917 171531 244983 171534
rect 231577 171458 231643 171461
rect 228988 171456 231643 171458
rect 228988 171400 231582 171456
rect 231638 171400 231643 171456
rect 228988 171398 231643 171400
rect 231577 171395 231643 171398
rect 264973 171458 265039 171461
rect 264973 171456 268180 171458
rect 264973 171400 264978 171456
rect 265034 171400 268180 171456
rect 264973 171398 268180 171400
rect 264973 171395 265039 171398
rect 213913 171050 213979 171053
rect 265065 171050 265131 171053
rect 213913 171048 217028 171050
rect 213913 170992 213918 171048
rect 213974 170992 217028 171048
rect 213913 170990 217028 170992
rect 265065 171048 268180 171050
rect 265065 170992 265070 171048
rect 265126 170992 268180 171048
rect 265065 170990 268180 170992
rect 213913 170987 213979 170990
rect 265065 170987 265131 170990
rect 231117 170914 231183 170917
rect 282821 170914 282887 170917
rect 228988 170912 231183 170914
rect 228988 170856 231122 170912
rect 231178 170856 231183 170912
rect 228988 170854 231183 170856
rect 279956 170912 282887 170914
rect 279956 170856 282826 170912
rect 282882 170856 282887 170912
rect 279956 170854 282887 170856
rect 231117 170851 231183 170854
rect 282821 170851 282887 170854
rect 279325 170642 279391 170645
rect 279325 170640 279434 170642
rect 279325 170584 279330 170640
rect 279386 170584 279434 170640
rect 279325 170579 279434 170584
rect 231945 170506 232011 170509
rect 228988 170504 232011 170506
rect 228988 170448 231950 170504
rect 232006 170448 232011 170504
rect 228988 170446 232011 170448
rect 231945 170443 232011 170446
rect 214005 170370 214071 170373
rect 214005 170368 217028 170370
rect 214005 170312 214010 170368
rect 214066 170312 217028 170368
rect 214005 170310 217028 170312
rect 214005 170307 214071 170310
rect 260281 170234 260347 170237
rect 268150 170234 268210 170476
rect 260281 170232 268210 170234
rect 260281 170176 260286 170232
rect 260342 170176 268210 170232
rect 279374 170204 279434 170579
rect 260281 170174 268210 170176
rect 260281 170171 260347 170174
rect 264973 170098 265039 170101
rect 264973 170096 268180 170098
rect 264973 170040 264978 170096
rect 265034 170040 268180 170096
rect 264973 170038 268180 170040
rect 264973 170035 265039 170038
rect 237465 169962 237531 169965
rect 228988 169960 237531 169962
rect 228988 169904 237470 169960
rect 237526 169904 237531 169960
rect 228988 169902 237531 169904
rect 237465 169899 237531 169902
rect 213913 169690 213979 169693
rect 265065 169690 265131 169693
rect 213913 169688 217028 169690
rect 213913 169632 213918 169688
rect 213974 169632 217028 169688
rect 213913 169630 217028 169632
rect 265065 169688 268180 169690
rect 265065 169632 265070 169688
rect 265126 169632 268180 169688
rect 265065 169630 268180 169632
rect 213913 169627 213979 169630
rect 265065 169627 265131 169630
rect 236085 169554 236151 169557
rect 228988 169552 236151 169554
rect 228988 169496 236090 169552
rect 236146 169496 236151 169552
rect 228988 169494 236151 169496
rect 236085 169491 236151 169494
rect 281533 169418 281599 169421
rect 279956 169416 281599 169418
rect 279956 169360 281538 169416
rect 281594 169360 281599 169416
rect 279956 169358 281599 169360
rect 281533 169355 281599 169358
rect 264973 169282 265039 169285
rect 264973 169280 268180 169282
rect 264973 169224 264978 169280
rect 265034 169224 268180 169280
rect 264973 169222 268180 169224
rect 264973 169219 265039 169222
rect 214005 169010 214071 169013
rect 231761 169010 231827 169013
rect 214005 169008 217028 169010
rect 214005 168952 214010 169008
rect 214066 168952 217028 169008
rect 214005 168950 217028 168952
rect 228988 169008 231827 169010
rect 228988 168952 231766 169008
rect 231822 168952 231827 169008
rect 228988 168950 231827 168952
rect 214005 168947 214071 168950
rect 231761 168947 231827 168950
rect 265157 168874 265223 168877
rect 265157 168872 268180 168874
rect 265157 168816 265162 168872
rect 265218 168816 268180 168872
rect 265157 168814 268180 168816
rect 265157 168811 265223 168814
rect 234889 168738 234955 168741
rect 237414 168738 237420 168740
rect 234889 168736 237420 168738
rect 234889 168680 234894 168736
rect 234950 168680 237420 168736
rect 234889 168678 237420 168680
rect 234889 168675 234955 168678
rect 237414 168676 237420 168678
rect 237484 168676 237490 168740
rect 282821 168738 282887 168741
rect 279956 168736 282887 168738
rect 279956 168680 282826 168736
rect 282882 168680 282887 168736
rect 279956 168678 282887 168680
rect 282821 168675 282887 168678
rect 255313 168602 255379 168605
rect 228988 168600 255379 168602
rect 228988 168544 255318 168600
rect 255374 168544 255379 168600
rect 228988 168542 255379 168544
rect 255313 168539 255379 168542
rect 253289 168466 253355 168469
rect 253289 168464 268180 168466
rect 253289 168408 253294 168464
rect 253350 168408 268180 168464
rect 253289 168406 268180 168408
rect 253289 168403 253355 168406
rect 213913 168330 213979 168333
rect 213913 168328 217028 168330
rect 213913 168272 213918 168328
rect 213974 168272 217028 168328
rect 213913 168270 217028 168272
rect 213913 168267 213979 168270
rect 279366 168268 279372 168332
rect 279436 168268 279442 168332
rect 231761 168058 231827 168061
rect 228988 168056 231827 168058
rect 228988 168000 231766 168056
rect 231822 168000 231827 168056
rect 228988 167998 231827 168000
rect 231761 167995 231827 167998
rect 264973 167922 265039 167925
rect 264973 167920 268180 167922
rect 264973 167864 264978 167920
rect 265034 167864 268180 167920
rect 279374 167892 279434 168268
rect 264973 167862 268180 167864
rect 264973 167859 265039 167862
rect 229369 167650 229435 167653
rect 228988 167648 229435 167650
rect 207657 167106 207723 167109
rect 216998 167106 217058 167620
rect 228988 167592 229374 167648
rect 229430 167592 229435 167648
rect 228988 167590 229435 167592
rect 229369 167587 229435 167590
rect 265065 167514 265131 167517
rect 265065 167512 268180 167514
rect 265065 167456 265070 167512
rect 265126 167456 268180 167512
rect 265065 167454 268180 167456
rect 265065 167451 265131 167454
rect 247125 167242 247191 167245
rect 238710 167240 247191 167242
rect 238710 167184 247130 167240
rect 247186 167184 247191 167240
rect 238710 167182 247191 167184
rect 238710 167106 238770 167182
rect 247125 167179 247191 167182
rect 207657 167104 217058 167106
rect 207657 167048 207662 167104
rect 207718 167048 217058 167104
rect 207657 167046 217058 167048
rect 228988 167046 238770 167106
rect 245101 167106 245167 167109
rect 282821 167106 282887 167109
rect 245101 167104 268180 167106
rect 245101 167048 245106 167104
rect 245162 167048 268180 167104
rect 245101 167046 268180 167048
rect 279956 167104 282887 167106
rect 279956 167048 282826 167104
rect 282882 167048 282887 167104
rect 279956 167046 282887 167048
rect 207657 167043 207723 167046
rect 245101 167043 245167 167046
rect 282821 167043 282887 167046
rect 213913 166970 213979 166973
rect 213913 166968 217028 166970
rect 213913 166912 213918 166968
rect 213974 166912 217028 166968
rect 213913 166910 217028 166912
rect 213913 166907 213979 166910
rect 231761 166698 231827 166701
rect 228988 166696 231827 166698
rect 228988 166640 231766 166696
rect 231822 166640 231827 166696
rect 228988 166638 231827 166640
rect 231761 166635 231827 166638
rect 264973 166698 265039 166701
rect 264973 166696 268180 166698
rect 264973 166640 264978 166696
rect 265034 166640 268180 166696
rect 264973 166638 268180 166640
rect 264973 166635 265039 166638
rect 214005 166426 214071 166429
rect 282821 166426 282887 166429
rect 583661 166426 583727 166429
rect 214005 166424 217028 166426
rect 214005 166368 214010 166424
rect 214066 166368 217028 166424
rect 214005 166366 217028 166368
rect 279956 166424 282887 166426
rect 279956 166368 282826 166424
rect 282882 166368 282887 166424
rect 279956 166366 282887 166368
rect 214005 166363 214071 166366
rect 282821 166363 282887 166366
rect 583526 166424 583727 166426
rect 583526 166368 583666 166424
rect 583722 166368 583727 166424
rect 583526 166366 583727 166368
rect 265341 166290 265407 166293
rect 265341 166288 268180 166290
rect 265341 166232 265346 166288
rect 265402 166232 268180 166288
rect 265341 166230 268180 166232
rect 265341 166227 265407 166230
rect 230749 166154 230815 166157
rect 228988 166152 230815 166154
rect 228988 166096 230754 166152
rect 230810 166096 230815 166152
rect 228988 166094 230815 166096
rect 230749 166091 230815 166094
rect 583526 166018 583586 166366
rect 583661 166363 583727 166366
rect 583342 165972 583586 166018
rect 583342 165958 584960 165972
rect 265709 165882 265775 165885
rect 583342 165882 583402 165958
rect 583520 165882 584960 165958
rect 265709 165880 268180 165882
rect 265709 165824 265714 165880
rect 265770 165824 268180 165880
rect 265709 165822 268180 165824
rect 583342 165822 584960 165882
rect 265709 165819 265775 165822
rect 207749 165746 207815 165749
rect 234705 165746 234771 165749
rect 207749 165744 217028 165746
rect 207749 165688 207754 165744
rect 207810 165688 217028 165744
rect 207749 165686 217028 165688
rect 228988 165744 234771 165746
rect 228988 165688 234710 165744
rect 234766 165688 234771 165744
rect 583520 165732 584960 165822
rect 228988 165686 234771 165688
rect 207749 165683 207815 165686
rect 234705 165683 234771 165686
rect 281993 165610 282059 165613
rect 279956 165608 282059 165610
rect 279956 165552 281998 165608
rect 282054 165552 282059 165608
rect 279956 165550 282059 165552
rect 281993 165547 282059 165550
rect 265065 165338 265131 165341
rect 265065 165336 268180 165338
rect 265065 165280 265070 165336
rect 265126 165280 268180 165336
rect 265065 165278 268180 165280
rect 265065 165275 265131 165278
rect 236494 165202 236500 165204
rect 228988 165142 236500 165202
rect 236494 165140 236500 165142
rect 236564 165140 236570 165204
rect 213913 165066 213979 165069
rect 213913 165064 217028 165066
rect 213913 165008 213918 165064
rect 213974 165008 217028 165064
rect 213913 165006 217028 165008
rect 213913 165003 213979 165006
rect 265617 164930 265683 164933
rect 280061 164930 280127 164933
rect 265617 164928 268180 164930
rect 265617 164872 265622 164928
rect 265678 164872 268180 164928
rect 265617 164870 268180 164872
rect 279956 164928 280127 164930
rect 279956 164872 280066 164928
rect 280122 164872 280127 164928
rect 279956 164870 280127 164872
rect 265617 164867 265683 164870
rect 280061 164867 280127 164870
rect 231485 164794 231551 164797
rect 228988 164792 231551 164794
rect 228988 164736 231490 164792
rect 231546 164736 231551 164792
rect 228988 164734 231551 164736
rect 231485 164731 231551 164734
rect 264973 164522 265039 164525
rect 264973 164520 268180 164522
rect 264973 164464 264978 164520
rect 265034 164464 268180 164520
rect 264973 164462 268180 164464
rect 264973 164459 265039 164462
rect 214005 164386 214071 164389
rect 229185 164386 229251 164389
rect 214005 164384 217028 164386
rect 214005 164328 214010 164384
rect 214066 164328 217028 164384
rect 214005 164326 217028 164328
rect 228988 164384 229251 164386
rect 228988 164328 229190 164384
rect 229246 164328 229251 164384
rect 228988 164326 229251 164328
rect 214005 164323 214071 164326
rect 229185 164323 229251 164326
rect 265065 164114 265131 164117
rect 282821 164114 282887 164117
rect 265065 164112 268180 164114
rect 265065 164056 265070 164112
rect 265126 164056 268180 164112
rect 265065 164054 268180 164056
rect 279956 164112 282887 164114
rect 279956 164056 282826 164112
rect 282882 164056 282887 164112
rect 279956 164054 282887 164056
rect 265065 164051 265131 164054
rect 282821 164051 282887 164054
rect 231761 163842 231827 163845
rect 228988 163840 231827 163842
rect 228988 163784 231766 163840
rect 231822 163784 231827 163840
rect 228988 163782 231827 163784
rect 231761 163779 231827 163782
rect 213913 163706 213979 163709
rect 264973 163706 265039 163709
rect 213913 163704 217028 163706
rect 213913 163648 213918 163704
rect 213974 163648 217028 163704
rect 213913 163646 217028 163648
rect 264973 163704 268180 163706
rect 264973 163648 264978 163704
rect 265034 163648 268180 163704
rect 264973 163646 268180 163648
rect 213913 163643 213979 163646
rect 264973 163643 265039 163646
rect 236177 163434 236243 163437
rect 228988 163432 236243 163434
rect 228988 163376 236182 163432
rect 236238 163376 236243 163432
rect 228988 163374 236243 163376
rect 236177 163371 236243 163374
rect 264513 163298 264579 163301
rect 282453 163298 282519 163301
rect 264513 163296 268180 163298
rect 264513 163240 264518 163296
rect 264574 163240 268180 163296
rect 264513 163238 268180 163240
rect 279956 163296 282519 163298
rect 279956 163240 282458 163296
rect 282514 163240 282519 163296
rect 279956 163238 282519 163240
rect 264513 163235 264579 163238
rect 282453 163235 282519 163238
rect 214005 163026 214071 163029
rect 214005 163024 217028 163026
rect -960 162890 480 162980
rect 214005 162968 214010 163024
rect 214066 162968 217028 163024
rect 214005 162966 217028 162968
rect 214005 162963 214071 162966
rect 3233 162890 3299 162893
rect 231669 162890 231735 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect 228988 162888 231735 162890
rect 228988 162832 231674 162888
rect 231730 162832 231735 162888
rect 228988 162830 231735 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 231669 162827 231735 162830
rect 232589 162890 232655 162893
rect 232589 162888 268180 162890
rect 232589 162832 232594 162888
rect 232650 162832 268180 162888
rect 232589 162830 268180 162832
rect 232589 162827 232655 162830
rect 282821 162618 282887 162621
rect 279956 162616 282887 162618
rect 279956 162560 282826 162616
rect 282882 162560 282887 162616
rect 279956 162558 282887 162560
rect 282821 162555 282887 162558
rect 231117 162482 231183 162485
rect 228988 162480 231183 162482
rect 228988 162424 231122 162480
rect 231178 162424 231183 162480
rect 228988 162422 231183 162424
rect 231117 162419 231183 162422
rect 213913 162346 213979 162349
rect 264973 162346 265039 162349
rect 213913 162344 217028 162346
rect 213913 162288 213918 162344
rect 213974 162288 217028 162344
rect 213913 162286 217028 162288
rect 264973 162344 268180 162346
rect 264973 162288 264978 162344
rect 265034 162288 268180 162344
rect 264973 162286 268180 162288
rect 213913 162283 213979 162286
rect 264973 162283 265039 162286
rect 230105 162210 230171 162213
rect 244406 162210 244412 162212
rect 230105 162208 244412 162210
rect 230105 162152 230110 162208
rect 230166 162152 244412 162208
rect 230105 162150 244412 162152
rect 230105 162147 230171 162150
rect 244406 162148 244412 162150
rect 244476 162148 244482 162212
rect 230749 162074 230815 162077
rect 249977 162074 250043 162077
rect 230749 162072 250043 162074
rect 230749 162016 230754 162072
rect 230810 162016 249982 162072
rect 250038 162016 250043 162072
rect 230749 162014 250043 162016
rect 230749 162011 230815 162014
rect 249977 162011 250043 162014
rect 231301 161938 231367 161941
rect 228988 161936 231367 161938
rect 228988 161880 231306 161936
rect 231362 161880 231367 161936
rect 228988 161878 231367 161880
rect 231301 161875 231367 161878
rect 258030 161878 268180 161938
rect 214005 161802 214071 161805
rect 255957 161802 256023 161805
rect 258030 161802 258090 161878
rect 282821 161802 282887 161805
rect 214005 161800 217028 161802
rect 214005 161744 214010 161800
rect 214066 161744 217028 161800
rect 214005 161742 217028 161744
rect 255957 161800 258090 161802
rect 255957 161744 255962 161800
rect 256018 161744 258090 161800
rect 255957 161742 258090 161744
rect 279956 161800 282887 161802
rect 279956 161744 282826 161800
rect 282882 161744 282887 161800
rect 279956 161742 282887 161744
rect 214005 161739 214071 161742
rect 255957 161739 256023 161742
rect 282821 161739 282887 161742
rect 231894 161530 231900 161532
rect 228988 161470 231900 161530
rect 231894 161468 231900 161470
rect 231964 161468 231970 161532
rect 263225 161530 263291 161533
rect 263225 161528 268180 161530
rect 263225 161472 263230 161528
rect 263286 161472 268180 161528
rect 263225 161470 268180 161472
rect 263225 161467 263291 161470
rect 279325 161394 279391 161397
rect 279325 161392 279434 161394
rect 279325 161336 279330 161392
rect 279386 161336 279434 161392
rect 279325 161331 279434 161336
rect 213913 161122 213979 161125
rect 264973 161122 265039 161125
rect 213913 161120 217028 161122
rect 213913 161064 213918 161120
rect 213974 161064 217028 161120
rect 213913 161062 217028 161064
rect 264973 161120 268180 161122
rect 264973 161064 264978 161120
rect 265034 161064 268180 161120
rect 279374 161092 279434 161331
rect 264973 161062 268180 161064
rect 213913 161059 213979 161062
rect 264973 161059 265039 161062
rect 231761 160986 231827 160989
rect 228988 160984 231827 160986
rect 228988 160928 231766 160984
rect 231822 160928 231827 160984
rect 228988 160926 231827 160928
rect 231761 160923 231827 160926
rect 230933 160578 230999 160581
rect 228988 160576 230999 160578
rect 228988 160520 230938 160576
rect 230994 160520 230999 160576
rect 228988 160518 230999 160520
rect 230933 160515 230999 160518
rect 214005 160442 214071 160445
rect 253197 160442 253263 160445
rect 268150 160442 268210 160684
rect 214005 160440 217028 160442
rect 214005 160384 214010 160440
rect 214066 160384 217028 160440
rect 214005 160382 217028 160384
rect 253197 160440 268210 160442
rect 253197 160384 253202 160440
rect 253258 160384 268210 160440
rect 253197 160382 268210 160384
rect 214005 160379 214071 160382
rect 253197 160379 253263 160382
rect 258717 160306 258783 160309
rect 282821 160306 282887 160309
rect 258717 160304 268180 160306
rect 258717 160248 258722 160304
rect 258778 160248 268180 160304
rect 258717 160246 268180 160248
rect 279956 160304 282887 160306
rect 279956 160248 282826 160304
rect 282882 160248 282887 160304
rect 279956 160246 282887 160248
rect 258717 160243 258783 160246
rect 282821 160243 282887 160246
rect 253933 160034 253999 160037
rect 228988 160032 253999 160034
rect 228988 159976 253938 160032
rect 253994 159976 253999 160032
rect 228988 159974 253999 159976
rect 253933 159971 253999 159974
rect 213913 159762 213979 159765
rect 265065 159762 265131 159765
rect 213913 159760 217028 159762
rect 213913 159704 213918 159760
rect 213974 159704 217028 159760
rect 213913 159702 217028 159704
rect 265065 159760 268180 159762
rect 265065 159704 265070 159760
rect 265126 159704 268180 159760
rect 265065 159702 268180 159704
rect 213913 159699 213979 159702
rect 265065 159699 265131 159702
rect 231761 159626 231827 159629
rect 228988 159624 231827 159626
rect 228988 159568 231766 159624
rect 231822 159568 231827 159624
rect 228988 159566 231827 159568
rect 231761 159563 231827 159566
rect 281901 159490 281967 159493
rect 279956 159488 281967 159490
rect 279956 159432 281906 159488
rect 281962 159432 281967 159488
rect 279956 159430 281967 159432
rect 281901 159427 281967 159430
rect 264973 159354 265039 159357
rect 264973 159352 268180 159354
rect 264973 159296 264978 159352
rect 265034 159296 268180 159352
rect 264973 159294 268180 159296
rect 264973 159291 265039 159294
rect 214005 159082 214071 159085
rect 230749 159082 230815 159085
rect 214005 159080 217028 159082
rect 214005 159024 214010 159080
rect 214066 159024 217028 159080
rect 214005 159022 217028 159024
rect 228988 159080 230815 159082
rect 228988 159024 230754 159080
rect 230810 159024 230815 159080
rect 228988 159022 230815 159024
rect 214005 159019 214071 159022
rect 230749 159019 230815 159022
rect 265157 158946 265223 158949
rect 265157 158944 268180 158946
rect 265157 158888 265162 158944
rect 265218 158888 268180 158944
rect 265157 158886 268180 158888
rect 265157 158883 265223 158886
rect 282361 158810 282427 158813
rect 279956 158808 282427 158810
rect 279956 158752 282366 158808
rect 282422 158752 282427 158808
rect 279956 158750 282427 158752
rect 282361 158747 282427 158750
rect 231761 158674 231827 158677
rect 228988 158672 231827 158674
rect 228988 158616 231766 158672
rect 231822 158616 231827 158672
rect 228988 158614 231827 158616
rect 231761 158611 231827 158614
rect 265249 158538 265315 158541
rect 265249 158536 268180 158538
rect 265249 158480 265254 158536
rect 265310 158480 268180 158536
rect 265249 158478 268180 158480
rect 265249 158475 265315 158478
rect 213913 158402 213979 158405
rect 213913 158400 217028 158402
rect 213913 158344 213918 158400
rect 213974 158344 217028 158400
rect 213913 158342 217028 158344
rect 213913 158339 213979 158342
rect 231209 158130 231275 158133
rect 228988 158128 231275 158130
rect 228988 158072 231214 158128
rect 231270 158072 231275 158128
rect 228988 158070 231275 158072
rect 231209 158067 231275 158070
rect 265065 158130 265131 158133
rect 265065 158128 268180 158130
rect 265065 158072 265070 158128
rect 265126 158072 268180 158128
rect 265065 158070 268180 158072
rect 265065 158067 265131 158070
rect 231485 157994 231551 157997
rect 245837 157994 245903 157997
rect 231485 157992 245903 157994
rect 231485 157936 231490 157992
rect 231546 157936 245842 157992
rect 245898 157936 245903 157992
rect 231485 157934 245903 157936
rect 231485 157931 231551 157934
rect 245837 157931 245903 157934
rect 251909 157994 251975 157997
rect 265157 157994 265223 157997
rect 282085 157994 282151 157997
rect 251909 157992 265223 157994
rect 251909 157936 251914 157992
rect 251970 157936 265162 157992
rect 265218 157936 265223 157992
rect 251909 157934 265223 157936
rect 279956 157992 282151 157994
rect 279956 157936 282090 157992
rect 282146 157936 282151 157992
rect 279956 157934 282151 157936
rect 251909 157931 251975 157934
rect 265157 157931 265223 157934
rect 282085 157931 282151 157934
rect 214005 157722 214071 157725
rect 230841 157722 230907 157725
rect 214005 157720 217028 157722
rect 214005 157664 214010 157720
rect 214066 157664 217028 157720
rect 214005 157662 217028 157664
rect 228988 157720 230907 157722
rect 228988 157664 230846 157720
rect 230902 157664 230907 157720
rect 228988 157662 230907 157664
rect 214005 157659 214071 157662
rect 230841 157659 230907 157662
rect 264973 157722 265039 157725
rect 264973 157720 268180 157722
rect 264973 157664 264978 157720
rect 265034 157664 268180 157720
rect 264973 157662 268180 157664
rect 264973 157659 265039 157662
rect 231669 157450 231735 157453
rect 234797 157450 234863 157453
rect 231669 157448 234863 157450
rect 231669 157392 231674 157448
rect 231730 157392 234802 157448
rect 234858 157392 234863 157448
rect 231669 157390 234863 157392
rect 231669 157387 231735 157390
rect 234797 157387 234863 157390
rect 281574 157314 281580 157316
rect 279956 157254 281580 157314
rect 281574 157252 281580 157254
rect 281644 157252 281650 157316
rect 213913 157178 213979 157181
rect 249793 157178 249859 157181
rect 213913 157176 217028 157178
rect 213913 157120 213918 157176
rect 213974 157120 217028 157176
rect 213913 157118 217028 157120
rect 228988 157176 249859 157178
rect 228988 157120 249798 157176
rect 249854 157120 249859 157176
rect 228988 157118 249859 157120
rect 213913 157115 213979 157118
rect 249793 157115 249859 157118
rect 264973 157178 265039 157181
rect 264973 157176 268180 157178
rect 264973 157120 264978 157176
rect 265034 157120 268180 157176
rect 264973 157118 268180 157120
rect 264973 157115 265039 157118
rect 244222 156770 244228 156772
rect 228988 156710 244228 156770
rect 244222 156708 244228 156710
rect 244292 156708 244298 156772
rect 214005 156498 214071 156501
rect 250437 156498 250503 156501
rect 268150 156498 268210 156740
rect 281809 156498 281875 156501
rect 214005 156496 217028 156498
rect 214005 156440 214010 156496
rect 214066 156440 217028 156496
rect 214005 156438 217028 156440
rect 250437 156496 268210 156498
rect 250437 156440 250442 156496
rect 250498 156440 268210 156496
rect 250437 156438 268210 156440
rect 279956 156496 281875 156498
rect 279956 156440 281814 156496
rect 281870 156440 281875 156496
rect 279956 156438 281875 156440
rect 214005 156435 214071 156438
rect 250437 156435 250503 156438
rect 281809 156435 281875 156438
rect 264329 156362 264395 156365
rect 264329 156360 268180 156362
rect 264329 156304 264334 156360
rect 264390 156304 268180 156360
rect 264329 156302 268180 156304
rect 264329 156299 264395 156302
rect 230933 156226 230999 156229
rect 228988 156224 230999 156226
rect 228988 156168 230938 156224
rect 230994 156168 230999 156224
rect 228988 156166 230999 156168
rect 230933 156163 230999 156166
rect 233325 155954 233391 155957
rect 233550 155954 233556 155956
rect 233325 155952 233556 155954
rect 233325 155896 233330 155952
rect 233386 155896 233556 155952
rect 233325 155894 233556 155896
rect 233325 155891 233391 155894
rect 233550 155892 233556 155894
rect 233620 155892 233626 155956
rect 265065 155954 265131 155957
rect 279325 155954 279391 155957
rect 265065 155952 268180 155954
rect 265065 155896 265070 155952
rect 265126 155896 268180 155952
rect 265065 155894 268180 155896
rect 279325 155952 279434 155954
rect 279325 155896 279330 155952
rect 279386 155896 279434 155952
rect 265065 155891 265131 155894
rect 279325 155891 279434 155896
rect 213913 155818 213979 155821
rect 230606 155818 230612 155820
rect 213913 155816 217028 155818
rect 213913 155760 213918 155816
rect 213974 155760 217028 155816
rect 213913 155758 217028 155760
rect 228988 155758 230612 155818
rect 213913 155755 213979 155758
rect 230606 155756 230612 155758
rect 230676 155756 230682 155820
rect 279374 155652 279434 155891
rect 267089 155546 267155 155549
rect 267089 155544 268180 155546
rect 267089 155488 267094 155544
rect 267150 155488 268180 155544
rect 267089 155486 268180 155488
rect 267089 155483 267155 155486
rect 230841 155274 230907 155277
rect 228988 155272 230907 155274
rect 228988 155216 230846 155272
rect 230902 155216 230907 155272
rect 228988 155214 230907 155216
rect 230841 155211 230907 155214
rect 230974 155212 230980 155276
rect 231044 155274 231050 155276
rect 240869 155274 240935 155277
rect 231044 155272 240935 155274
rect 231044 155216 240874 155272
rect 240930 155216 240935 155272
rect 231044 155214 240935 155216
rect 231044 155212 231050 155214
rect 240869 155211 240935 155214
rect 214005 155138 214071 155141
rect 214005 155136 217028 155138
rect 214005 155080 214010 155136
rect 214066 155080 217028 155136
rect 214005 155078 217028 155080
rect 258030 155078 268180 155138
rect 214005 155075 214071 155078
rect 232681 155002 232747 155005
rect 258030 155002 258090 155078
rect 282269 155002 282335 155005
rect 232681 155000 258090 155002
rect 232681 154944 232686 155000
rect 232742 154944 258090 155000
rect 232681 154942 258090 154944
rect 279956 155000 282335 155002
rect 279956 154944 282274 155000
rect 282330 154944 282335 155000
rect 279956 154942 282335 154944
rect 232681 154939 232747 154942
rect 282269 154939 282335 154942
rect 233182 154866 233188 154868
rect 228988 154806 233188 154866
rect 233182 154804 233188 154806
rect 233252 154804 233258 154868
rect 264973 154594 265039 154597
rect 264973 154592 268180 154594
rect 264973 154536 264978 154592
rect 265034 154536 268180 154592
rect 264973 154534 268180 154536
rect 264973 154531 265039 154534
rect 214005 154458 214071 154461
rect 214005 154456 217028 154458
rect 214005 154400 214010 154456
rect 214066 154400 217028 154456
rect 214005 154398 217028 154400
rect 214005 154395 214071 154398
rect 231669 154322 231735 154325
rect 228988 154320 231735 154322
rect 228988 154264 231674 154320
rect 231730 154264 231735 154320
rect 228988 154262 231735 154264
rect 231669 154259 231735 154262
rect 265341 154186 265407 154189
rect 282821 154186 282887 154189
rect 265341 154184 268180 154186
rect 265341 154128 265346 154184
rect 265402 154128 268180 154184
rect 265341 154126 268180 154128
rect 279956 154184 282887 154186
rect 279956 154128 282826 154184
rect 282882 154128 282887 154184
rect 279956 154126 282887 154128
rect 265341 154123 265407 154126
rect 282821 154123 282887 154126
rect 231301 153914 231367 153917
rect 228988 153912 231367 153914
rect 228988 153856 231306 153912
rect 231362 153856 231367 153912
rect 228988 153854 231367 153856
rect 231301 153851 231367 153854
rect 213913 153778 213979 153781
rect 230841 153778 230907 153781
rect 238845 153778 238911 153781
rect 213913 153776 217028 153778
rect 213913 153720 213918 153776
rect 213974 153720 217028 153776
rect 213913 153718 217028 153720
rect 230841 153776 238911 153778
rect 230841 153720 230846 153776
rect 230902 153720 238850 153776
rect 238906 153720 238911 153776
rect 230841 153718 238911 153720
rect 213913 153715 213979 153718
rect 230841 153715 230907 153718
rect 238845 153715 238911 153718
rect 265157 153778 265223 153781
rect 265157 153776 268180 153778
rect 265157 153720 265162 153776
rect 265218 153720 268180 153776
rect 265157 153718 268180 153720
rect 265157 153715 265223 153718
rect 282269 153506 282335 153509
rect 279956 153504 282335 153506
rect 279956 153448 282274 153504
rect 282330 153448 282335 153504
rect 279956 153446 282335 153448
rect 282269 153443 282335 153446
rect 238753 153370 238819 153373
rect 228988 153368 238819 153370
rect 228988 153312 238758 153368
rect 238814 153312 238819 153368
rect 228988 153310 238819 153312
rect 238753 153307 238819 153310
rect 258030 153310 268180 153370
rect 239581 153234 239647 153237
rect 258030 153234 258090 153310
rect 239581 153232 258090 153234
rect 239581 153176 239586 153232
rect 239642 153176 258090 153232
rect 239581 153174 258090 153176
rect 239581 153171 239647 153174
rect 213177 153098 213243 153101
rect 213177 153096 217028 153098
rect 213177 153040 213182 153096
rect 213238 153040 217028 153096
rect 213177 153038 217028 153040
rect 213177 153035 213243 153038
rect 231485 152962 231551 152965
rect 228988 152960 231551 152962
rect 228988 152904 231490 152960
rect 231546 152904 231551 152960
rect 228988 152902 231551 152904
rect 231485 152899 231551 152902
rect 265065 152962 265131 152965
rect 265065 152960 268180 152962
rect 265065 152904 265070 152960
rect 265126 152904 268180 152960
rect 265065 152902 268180 152904
rect 265065 152899 265131 152902
rect 281717 152690 281783 152693
rect 279956 152688 281783 152690
rect 279956 152632 281722 152688
rect 281778 152632 281783 152688
rect 279956 152630 281783 152632
rect 281717 152627 281783 152630
rect 583293 152690 583359 152693
rect 583520 152690 584960 152780
rect 583293 152688 584960 152690
rect 583293 152632 583298 152688
rect 583354 152632 584960 152688
rect 583293 152630 584960 152632
rect 583293 152627 583359 152630
rect 213913 152554 213979 152557
rect 232078 152554 232084 152556
rect 213913 152552 217028 152554
rect 213913 152496 213918 152552
rect 213974 152496 217028 152552
rect 213913 152494 217028 152496
rect 228988 152494 232084 152554
rect 213913 152491 213979 152494
rect 232078 152492 232084 152494
rect 232148 152492 232154 152556
rect 265249 152554 265315 152557
rect 265249 152552 268180 152554
rect 265249 152496 265254 152552
rect 265310 152496 268180 152552
rect 583520 152540 584960 152630
rect 265249 152494 268180 152496
rect 265249 152491 265315 152494
rect 249926 152010 249932 152012
rect 228988 151950 249932 152010
rect 249926 151948 249932 151950
rect 249996 151948 250002 152012
rect 264973 152010 265039 152013
rect 264973 152008 268180 152010
rect 264973 151952 264978 152008
rect 265034 151952 268180 152008
rect 264973 151950 268180 151952
rect 264973 151947 265039 151950
rect 214649 151874 214715 151877
rect 281533 151874 281599 151877
rect 214649 151872 217028 151874
rect 214649 151816 214654 151872
rect 214710 151816 217028 151872
rect 214649 151814 217028 151816
rect 279956 151872 281599 151874
rect 279956 151816 281538 151872
rect 281594 151816 281599 151872
rect 279956 151814 281599 151816
rect 214649 151811 214715 151814
rect 281533 151811 281599 151814
rect 230473 151602 230539 151605
rect 228988 151600 230539 151602
rect 228988 151544 230478 151600
rect 230534 151544 230539 151600
rect 228988 151542 230539 151544
rect 230473 151539 230539 151542
rect 260189 151330 260255 151333
rect 268150 151330 268210 151572
rect 260189 151328 268210 151330
rect 260189 151272 260194 151328
rect 260250 151272 268210 151328
rect 260189 151270 268210 151272
rect 260189 151267 260255 151270
rect 214097 151194 214163 151197
rect 264973 151194 265039 151197
rect 281901 151194 281967 151197
rect 214097 151192 217028 151194
rect 214097 151136 214102 151192
rect 214158 151136 217028 151192
rect 214097 151134 217028 151136
rect 264973 151192 268180 151194
rect 264973 151136 264978 151192
rect 265034 151136 268180 151192
rect 264973 151134 268180 151136
rect 279956 151192 281967 151194
rect 279956 151136 281906 151192
rect 281962 151136 281967 151192
rect 279956 151134 281967 151136
rect 214097 151131 214163 151134
rect 264973 151131 265039 151134
rect 281901 151131 281967 151134
rect 169201 151058 169267 151061
rect 214649 151058 214715 151061
rect 241462 151058 241468 151060
rect 169201 151056 214715 151058
rect 169201 151000 169206 151056
rect 169262 151000 214654 151056
rect 214710 151000 214715 151056
rect 169201 150998 214715 151000
rect 228988 150998 241468 151058
rect 169201 150995 169267 150998
rect 214649 150995 214715 150998
rect 241462 150996 241468 150998
rect 241532 150996 241538 151060
rect 265341 150786 265407 150789
rect 265341 150784 268180 150786
rect 265341 150728 265346 150784
rect 265402 150728 268180 150784
rect 265341 150726 268180 150728
rect 265341 150723 265407 150726
rect 231761 150650 231827 150653
rect 228988 150648 231827 150650
rect 228988 150592 231766 150648
rect 231822 150592 231827 150648
rect 228988 150590 231827 150592
rect 231761 150587 231827 150590
rect 213913 150514 213979 150517
rect 213913 150512 217028 150514
rect 213913 150456 213918 150512
rect 213974 150456 217028 150512
rect 213913 150454 217028 150456
rect 213913 150451 213979 150454
rect 280245 150378 280311 150381
rect 279956 150376 280311 150378
rect 231577 150106 231643 150109
rect 228988 150104 231643 150106
rect 228988 150048 231582 150104
rect 231638 150048 231643 150104
rect 228988 150046 231643 150048
rect 231577 150043 231643 150046
rect 236913 150106 236979 150109
rect 268150 150106 268210 150348
rect 279956 150320 280250 150376
rect 280306 150320 280311 150376
rect 279956 150318 280311 150320
rect 280245 150315 280311 150318
rect 236913 150104 268210 150106
rect 236913 150048 236918 150104
rect 236974 150048 268210 150104
rect 236913 150046 268210 150048
rect 236913 150043 236979 150046
rect 264973 149970 265039 149973
rect 264973 149968 268180 149970
rect -960 149834 480 149924
rect 264973 149912 264978 149968
rect 265034 149912 268180 149968
rect 264973 149910 268180 149912
rect 264973 149907 265039 149910
rect 2773 149834 2839 149837
rect -960 149832 2839 149834
rect -960 149776 2778 149832
rect 2834 149776 2839 149832
rect -960 149774 2839 149776
rect -960 149684 480 149774
rect 2773 149771 2839 149774
rect 213913 149834 213979 149837
rect 213913 149832 217028 149834
rect 213913 149776 213918 149832
rect 213974 149776 217028 149832
rect 213913 149774 217028 149776
rect 213913 149771 213979 149774
rect 230422 149698 230428 149700
rect 228988 149638 230428 149698
rect 230422 149636 230428 149638
rect 230492 149636 230498 149700
rect 231669 149698 231735 149701
rect 241830 149698 241836 149700
rect 231669 149696 241836 149698
rect 231669 149640 231674 149696
rect 231730 149640 241836 149696
rect 231669 149638 241836 149640
rect 231669 149635 231735 149638
rect 241830 149636 241836 149638
rect 241900 149636 241906 149700
rect 265893 149562 265959 149565
rect 265893 149560 268180 149562
rect 265893 149504 265898 149560
rect 265954 149504 268180 149560
rect 265893 149502 268180 149504
rect 265893 149499 265959 149502
rect 230289 149290 230355 149293
rect 237598 149290 237604 149292
rect 230289 149288 237604 149290
rect 230289 149232 230294 149288
rect 230350 149232 237604 149288
rect 230289 149230 237604 149232
rect 230289 149227 230355 149230
rect 237598 149228 237604 149230
rect 237668 149228 237674 149292
rect 214005 149154 214071 149157
rect 230565 149154 230631 149157
rect 214005 149152 217028 149154
rect 214005 149096 214010 149152
rect 214066 149096 217028 149152
rect 214005 149094 217028 149096
rect 228988 149152 230631 149154
rect 228988 149096 230570 149152
rect 230626 149096 230631 149152
rect 228988 149094 230631 149096
rect 279926 149154 279986 149668
rect 291326 149154 291332 149156
rect 279926 149094 291332 149154
rect 214005 149091 214071 149094
rect 230565 149091 230631 149094
rect 291326 149092 291332 149094
rect 291396 149092 291402 149156
rect 264973 149018 265039 149021
rect 264973 149016 268180 149018
rect 264973 148960 264978 149016
rect 265034 148960 268180 149016
rect 264973 148958 268180 148960
rect 264973 148955 265039 148958
rect 282637 148882 282703 148885
rect 279956 148880 282703 148882
rect 279956 148824 282642 148880
rect 282698 148824 282703 148880
rect 279956 148822 282703 148824
rect 282637 148819 282703 148822
rect 231761 148746 231827 148749
rect 228988 148744 231827 148746
rect 228988 148688 231766 148744
rect 231822 148688 231827 148744
rect 228988 148686 231827 148688
rect 231761 148683 231827 148686
rect 265065 148610 265131 148613
rect 265065 148608 268180 148610
rect 265065 148552 265070 148608
rect 265126 148552 268180 148608
rect 265065 148550 268180 148552
rect 265065 148547 265131 148550
rect 214557 148474 214623 148477
rect 214557 148472 217028 148474
rect 214557 148416 214562 148472
rect 214618 148416 217028 148472
rect 214557 148414 217028 148416
rect 214557 148411 214623 148414
rect 229737 148202 229803 148205
rect 228988 148200 229803 148202
rect 228988 148144 229742 148200
rect 229798 148144 229803 148200
rect 228988 148142 229803 148144
rect 229737 148139 229803 148142
rect 258030 148142 268180 148202
rect 230381 148066 230447 148069
rect 258030 148066 258090 148142
rect 282821 148066 282887 148069
rect 230381 148064 258090 148066
rect 230381 148008 230386 148064
rect 230442 148008 258090 148064
rect 230381 148006 258090 148008
rect 279956 148064 282887 148066
rect 279956 148008 282826 148064
rect 282882 148008 282887 148064
rect 279956 148006 282887 148008
rect 230381 148003 230447 148006
rect 282821 148003 282887 148006
rect 213913 147930 213979 147933
rect 213913 147928 217028 147930
rect 213913 147872 213918 147928
rect 213974 147872 217028 147928
rect 213913 147870 217028 147872
rect 213913 147867 213979 147870
rect 230657 147794 230723 147797
rect 228988 147792 230723 147794
rect 228988 147736 230662 147792
rect 230718 147736 230723 147792
rect 228988 147734 230723 147736
rect 230657 147731 230723 147734
rect 262857 147794 262923 147797
rect 262857 147792 268180 147794
rect 262857 147736 262862 147792
rect 262918 147736 268180 147792
rect 262857 147734 268180 147736
rect 262857 147731 262923 147734
rect 264973 147386 265039 147389
rect 282821 147386 282887 147389
rect 264973 147384 268180 147386
rect 264973 147328 264978 147384
rect 265034 147328 268180 147384
rect 264973 147326 268180 147328
rect 279956 147384 282887 147386
rect 279956 147328 282826 147384
rect 282882 147328 282887 147384
rect 279956 147326 282887 147328
rect 264973 147323 265039 147326
rect 282821 147323 282887 147326
rect 213913 147250 213979 147253
rect 240542 147250 240548 147252
rect 213913 147248 217028 147250
rect 213913 147192 213918 147248
rect 213974 147192 217028 147248
rect 213913 147190 217028 147192
rect 228988 147190 240548 147250
rect 213913 147187 213979 147190
rect 240542 147188 240548 147190
rect 240612 147188 240618 147252
rect 264421 146978 264487 146981
rect 264421 146976 268180 146978
rect 264421 146920 264426 146976
rect 264482 146920 268180 146976
rect 264421 146918 268180 146920
rect 264421 146915 264487 146918
rect 229093 146842 229159 146845
rect 228988 146840 229159 146842
rect 228988 146784 229098 146840
rect 229154 146784 229159 146840
rect 228988 146782 229159 146784
rect 229093 146779 229159 146782
rect 216121 146570 216187 146573
rect 282269 146570 282335 146573
rect 216121 146568 217028 146570
rect 216121 146512 216126 146568
rect 216182 146512 217028 146568
rect 216121 146510 217028 146512
rect 279956 146568 282335 146570
rect 279956 146512 282274 146568
rect 282330 146512 282335 146568
rect 279956 146510 282335 146512
rect 216121 146507 216187 146510
rect 282269 146507 282335 146510
rect 238293 146434 238359 146437
rect 238293 146432 268180 146434
rect 238293 146376 238298 146432
rect 238354 146376 268180 146432
rect 238293 146374 268180 146376
rect 238293 146371 238359 146374
rect 229318 146298 229324 146300
rect 228988 146238 229324 146298
rect 229318 146236 229324 146238
rect 229388 146236 229394 146300
rect 265065 146026 265131 146029
rect 265065 146024 268180 146026
rect 265065 145968 265070 146024
rect 265126 145968 268180 146024
rect 265065 145966 268180 145968
rect 265065 145963 265131 145966
rect 214005 145890 214071 145893
rect 230841 145890 230907 145893
rect 282821 145890 282887 145893
rect 214005 145888 217028 145890
rect 214005 145832 214010 145888
rect 214066 145832 217028 145888
rect 214005 145830 217028 145832
rect 228988 145888 230907 145890
rect 228988 145832 230846 145888
rect 230902 145832 230907 145888
rect 228988 145830 230907 145832
rect 279956 145888 282887 145890
rect 279956 145832 282826 145888
rect 282882 145832 282887 145888
rect 279956 145830 282887 145832
rect 214005 145827 214071 145830
rect 230841 145827 230907 145830
rect 282821 145827 282887 145830
rect 189717 145618 189783 145621
rect 207749 145618 207815 145621
rect 189717 145616 207815 145618
rect 189717 145560 189722 145616
rect 189778 145560 207754 145616
rect 207810 145560 207815 145616
rect 189717 145558 207815 145560
rect 189717 145555 189783 145558
rect 207749 145555 207815 145558
rect 233550 145346 233556 145348
rect 228988 145286 233556 145346
rect 233550 145284 233556 145286
rect 233620 145284 233626 145348
rect 233734 145284 233740 145348
rect 233804 145346 233810 145348
rect 268150 145346 268210 145588
rect 233804 145286 268210 145346
rect 233804 145284 233810 145286
rect 213913 145210 213979 145213
rect 264973 145210 265039 145213
rect 213913 145208 217028 145210
rect 213913 145152 213918 145208
rect 213974 145152 217028 145208
rect 213913 145150 217028 145152
rect 264973 145208 268180 145210
rect 264973 145152 264978 145208
rect 265034 145152 268180 145208
rect 264973 145150 268180 145152
rect 213913 145147 213979 145150
rect 264973 145147 265039 145150
rect 282729 145074 282795 145077
rect 279956 145072 282795 145074
rect 279956 145016 282734 145072
rect 282790 145016 282795 145072
rect 279956 145014 282795 145016
rect 282729 145011 282795 145014
rect 231669 144938 231735 144941
rect 228988 144936 231735 144938
rect 228988 144880 231674 144936
rect 231730 144880 231735 144936
rect 228988 144878 231735 144880
rect 231669 144875 231735 144878
rect 251173 144802 251239 144805
rect 238710 144800 251239 144802
rect 238710 144744 251178 144800
rect 251234 144744 251239 144800
rect 238710 144742 251239 144744
rect 214005 144530 214071 144533
rect 214005 144528 217028 144530
rect 214005 144472 214010 144528
rect 214066 144472 217028 144528
rect 214005 144470 217028 144472
rect 214005 144467 214071 144470
rect 238710 144394 238770 144742
rect 251173 144739 251239 144742
rect 265065 144802 265131 144805
rect 265065 144800 268180 144802
rect 265065 144744 265070 144800
rect 265126 144744 268180 144800
rect 265065 144742 268180 144744
rect 265065 144739 265131 144742
rect 228988 144334 238770 144394
rect 264973 144394 265039 144397
rect 264973 144392 268180 144394
rect 264973 144336 264978 144392
rect 265034 144336 268180 144392
rect 264973 144334 268180 144336
rect 264973 144331 265039 144334
rect 282821 144258 282887 144261
rect 279956 144256 282887 144258
rect 279956 144200 282826 144256
rect 282882 144200 282887 144256
rect 279956 144198 282887 144200
rect 282821 144195 282887 144198
rect 252093 144122 252159 144125
rect 265341 144122 265407 144125
rect 252093 144120 265407 144122
rect 252093 144064 252098 144120
rect 252154 144064 265346 144120
rect 265402 144064 265407 144120
rect 252093 144062 265407 144064
rect 252093 144059 252159 144062
rect 265341 144059 265407 144062
rect 231761 143986 231827 143989
rect 228988 143984 231827 143986
rect 228988 143928 231766 143984
rect 231822 143928 231827 143984
rect 228988 143926 231827 143928
rect 231761 143923 231827 143926
rect 213913 143850 213979 143853
rect 265157 143850 265223 143853
rect 213913 143848 217028 143850
rect 213913 143792 213918 143848
rect 213974 143792 217028 143848
rect 213913 143790 217028 143792
rect 265157 143848 268180 143850
rect 265157 143792 265162 143848
rect 265218 143792 268180 143848
rect 265157 143790 268180 143792
rect 213913 143787 213979 143790
rect 265157 143787 265223 143790
rect 283782 143578 283788 143580
rect 279956 143518 283788 143578
rect 283782 143516 283788 143518
rect 283852 143516 283858 143580
rect 231761 143442 231827 143445
rect 228988 143440 231827 143442
rect 228988 143384 231766 143440
rect 231822 143384 231827 143440
rect 228988 143382 231827 143384
rect 231761 143379 231827 143382
rect 265065 143442 265131 143445
rect 265065 143440 268180 143442
rect 265065 143384 265070 143440
rect 265126 143384 268180 143440
rect 265065 143382 268180 143384
rect 265065 143379 265131 143382
rect 214005 143306 214071 143309
rect 231761 143306 231827 143309
rect 240358 143306 240364 143308
rect 214005 143304 217028 143306
rect 214005 143248 214010 143304
rect 214066 143248 217028 143304
rect 214005 143246 217028 143248
rect 231761 143304 240364 143306
rect 231761 143248 231766 143304
rect 231822 143248 240364 143304
rect 231761 143246 240364 143248
rect 214005 143243 214071 143246
rect 231761 143243 231827 143246
rect 240358 143244 240364 143246
rect 240428 143244 240434 143308
rect 252829 143034 252895 143037
rect 228988 143032 252895 143034
rect 228988 142976 252834 143032
rect 252890 142976 252895 143032
rect 228988 142974 252895 142976
rect 252829 142971 252895 142974
rect 265249 143034 265315 143037
rect 265249 143032 268180 143034
rect 265249 142976 265254 143032
rect 265310 142976 268180 143032
rect 265249 142974 268180 142976
rect 265249 142971 265315 142974
rect 282821 142762 282887 142765
rect 279956 142760 282887 142762
rect 279956 142704 282826 142760
rect 282882 142704 282887 142760
rect 279956 142702 282887 142704
rect 282821 142699 282887 142702
rect 213913 142626 213979 142629
rect 213913 142624 217028 142626
rect 213913 142568 213918 142624
rect 213974 142568 217028 142624
rect 213913 142566 217028 142568
rect 258030 142566 268180 142626
rect 213913 142563 213979 142566
rect 231761 142490 231827 142493
rect 228988 142488 231827 142490
rect 228988 142432 231766 142488
rect 231822 142432 231827 142488
rect 228988 142430 231827 142432
rect 231761 142427 231827 142430
rect 249333 142490 249399 142493
rect 258030 142490 258090 142566
rect 249333 142488 258090 142490
rect 249333 142432 249338 142488
rect 249394 142432 258090 142488
rect 249333 142430 258090 142432
rect 249333 142427 249399 142430
rect 264973 142218 265039 142221
rect 264973 142216 268180 142218
rect 264973 142160 264978 142216
rect 265034 142160 268180 142216
rect 264973 142158 268180 142160
rect 264973 142155 265039 142158
rect 230565 142082 230631 142085
rect 282545 142082 282611 142085
rect 228988 142080 230631 142082
rect 228988 142024 230570 142080
rect 230626 142024 230631 142080
rect 228988 142022 230631 142024
rect 279956 142080 282611 142082
rect 279956 142024 282550 142080
rect 282606 142024 282611 142080
rect 279956 142022 282611 142024
rect 230565 142019 230631 142022
rect 282545 142019 282611 142022
rect 213913 141946 213979 141949
rect 213913 141944 217028 141946
rect 213913 141888 213918 141944
rect 213974 141888 217028 141944
rect 213913 141886 217028 141888
rect 213913 141883 213979 141886
rect 264973 141810 265039 141813
rect 264973 141808 268180 141810
rect 264973 141752 264978 141808
rect 265034 141752 268180 141808
rect 264973 141750 268180 141752
rect 264973 141747 265039 141750
rect 245653 141674 245719 141677
rect 228988 141672 245719 141674
rect 228988 141616 245658 141672
rect 245714 141616 245719 141672
rect 228988 141614 245719 141616
rect 245653 141611 245719 141614
rect 244774 141340 244780 141404
rect 244844 141402 244850 141404
rect 265157 141402 265223 141405
rect 244844 141400 265223 141402
rect 244844 141344 265162 141400
rect 265218 141344 265223 141400
rect 244844 141342 265223 141344
rect 244844 141340 244850 141342
rect 265157 141339 265223 141342
rect 214005 141266 214071 141269
rect 265065 141266 265131 141269
rect 282821 141266 282887 141269
rect 214005 141264 217028 141266
rect 214005 141208 214010 141264
rect 214066 141208 217028 141264
rect 214005 141206 217028 141208
rect 265065 141264 268180 141266
rect 265065 141208 265070 141264
rect 265126 141208 268180 141264
rect 265065 141206 268180 141208
rect 279956 141264 282887 141266
rect 279956 141208 282826 141264
rect 282882 141208 282887 141264
rect 279956 141206 282887 141208
rect 214005 141203 214071 141206
rect 265065 141203 265131 141206
rect 282821 141203 282887 141206
rect 238937 141130 239003 141133
rect 228988 141128 239003 141130
rect 228988 141072 238942 141128
rect 238998 141072 239003 141128
rect 228988 141070 239003 141072
rect 238937 141067 239003 141070
rect 265157 140858 265223 140861
rect 265157 140856 268180 140858
rect 265157 140800 265162 140856
rect 265218 140800 268180 140856
rect 265157 140798 268180 140800
rect 265157 140795 265223 140798
rect 231761 140722 231827 140725
rect 228988 140720 231827 140722
rect 228988 140664 231766 140720
rect 231822 140664 231827 140720
rect 228988 140662 231827 140664
rect 231761 140659 231827 140662
rect 213913 140586 213979 140589
rect 213913 140584 217028 140586
rect 213913 140528 213918 140584
rect 213974 140528 217028 140584
rect 213913 140526 217028 140528
rect 213913 140523 213979 140526
rect 284334 140450 284340 140452
rect 251214 140178 251220 140180
rect 228988 140118 251220 140178
rect 251214 140116 251220 140118
rect 251284 140116 251290 140180
rect 260046 140116 260052 140180
rect 260116 140178 260122 140180
rect 268150 140178 268210 140420
rect 279956 140390 284340 140450
rect 284334 140388 284340 140390
rect 284404 140388 284410 140452
rect 260116 140118 268210 140178
rect 260116 140116 260122 140118
rect 231158 139980 231164 140044
rect 231228 140042 231234 140044
rect 258809 140042 258875 140045
rect 231228 140040 258875 140042
rect 231228 139984 258814 140040
rect 258870 139984 258875 140040
rect 231228 139982 258875 139984
rect 231228 139980 231234 139982
rect 258809 139979 258875 139982
rect 214097 139906 214163 139909
rect 214097 139904 217028 139906
rect 214097 139848 214102 139904
rect 214158 139848 217028 139904
rect 214097 139846 217028 139848
rect 214097 139843 214163 139846
rect 233366 139770 233372 139772
rect 228988 139710 233372 139770
rect 233366 139708 233372 139710
rect 233436 139708 233442 139772
rect 246389 139770 246455 139773
rect 268150 139770 268210 140012
rect 282821 139770 282887 139773
rect 246389 139768 268210 139770
rect 246389 139712 246394 139768
rect 246450 139712 268210 139768
rect 246389 139710 268210 139712
rect 279956 139768 282887 139770
rect 279956 139712 282826 139768
rect 282882 139712 282887 139768
rect 279956 139710 282887 139712
rect 246389 139707 246455 139710
rect 282821 139707 282887 139710
rect 264973 139634 265039 139637
rect 264973 139632 268180 139634
rect 264973 139576 264978 139632
rect 265034 139576 268180 139632
rect 264973 139574 268180 139576
rect 264973 139571 265039 139574
rect 583201 139362 583267 139365
rect 583520 139362 584960 139452
rect 583201 139360 584960 139362
rect 583201 139304 583206 139360
rect 583262 139304 584960 139360
rect 583201 139302 584960 139304
rect 583201 139299 583267 139302
rect 213913 139226 213979 139229
rect 234654 139226 234660 139228
rect 213913 139224 217028 139226
rect 213913 139168 213918 139224
rect 213974 139168 217028 139224
rect 213913 139166 217028 139168
rect 228988 139166 234660 139226
rect 213913 139163 213979 139166
rect 234654 139164 234660 139166
rect 234724 139164 234730 139228
rect 583520 139212 584960 139302
rect 265065 138954 265131 138957
rect 258030 138952 265131 138954
rect 258030 138896 265070 138952
rect 265126 138896 265131 138952
rect 258030 138894 265131 138896
rect 230289 138818 230355 138821
rect 228988 138816 230355 138818
rect 228988 138760 230294 138816
rect 230350 138760 230355 138816
rect 228988 138758 230355 138760
rect 230289 138755 230355 138758
rect 214649 138682 214715 138685
rect 214649 138680 217028 138682
rect 214649 138624 214654 138680
rect 214710 138624 217028 138680
rect 214649 138622 217028 138624
rect 214649 138619 214715 138622
rect 232446 138620 232452 138684
rect 232516 138682 232522 138684
rect 258030 138682 258090 138894
rect 265065 138891 265131 138894
rect 268150 138818 268210 139196
rect 281533 138954 281599 138957
rect 279956 138952 281599 138954
rect 279956 138896 281538 138952
rect 281594 138896 281599 138952
rect 279956 138894 281599 138896
rect 281533 138891 281599 138894
rect 232516 138622 258090 138682
rect 262814 138758 268210 138818
rect 232516 138620 232522 138622
rect 229737 138410 229803 138413
rect 262814 138410 262874 138758
rect 265801 138682 265867 138685
rect 265801 138680 268180 138682
rect 265801 138624 265806 138680
rect 265862 138624 268180 138680
rect 265801 138622 268180 138624
rect 265801 138619 265867 138622
rect 229737 138408 262874 138410
rect 229737 138352 229742 138408
rect 229798 138352 262874 138408
rect 229737 138350 262874 138352
rect 229737 138347 229803 138350
rect 230105 138274 230171 138277
rect 228988 138272 230171 138274
rect 228988 138216 230110 138272
rect 230166 138216 230171 138272
rect 228988 138214 230171 138216
rect 230105 138211 230171 138214
rect 264973 138274 265039 138277
rect 281533 138274 281599 138277
rect 264973 138272 268180 138274
rect 264973 138216 264978 138272
rect 265034 138216 268180 138272
rect 264973 138214 268180 138216
rect 279956 138272 281599 138274
rect 279956 138216 281538 138272
rect 281594 138216 281599 138272
rect 279956 138214 281599 138216
rect 264973 138211 265039 138214
rect 281533 138211 281599 138214
rect 216029 138002 216095 138005
rect 216029 138000 217028 138002
rect 216029 137944 216034 138000
rect 216090 137944 217028 138000
rect 216029 137942 217028 137944
rect 216029 137939 216095 137942
rect 231761 137866 231827 137869
rect 228988 137864 231827 137866
rect 228988 137808 231766 137864
rect 231822 137808 231827 137864
rect 228988 137806 231827 137808
rect 231761 137803 231827 137806
rect 265065 137866 265131 137869
rect 265065 137864 268180 137866
rect 265065 137808 265070 137864
rect 265126 137808 268180 137864
rect 265065 137806 268180 137808
rect 265065 137803 265131 137806
rect 282821 137458 282887 137461
rect 279956 137456 282887 137458
rect 213913 137322 213979 137325
rect 229134 137322 229140 137324
rect 213913 137320 217028 137322
rect 213913 137264 213918 137320
rect 213974 137264 217028 137320
rect 213913 137262 217028 137264
rect 228988 137262 229140 137322
rect 213913 137259 213979 137262
rect 229134 137260 229140 137262
rect 229204 137260 229210 137324
rect 239397 137186 239463 137189
rect 268150 137186 268210 137428
rect 279956 137400 282826 137456
rect 282882 137400 282887 137456
rect 279956 137398 282887 137400
rect 282821 137395 282887 137398
rect 239397 137184 268210 137186
rect 239397 137128 239402 137184
rect 239458 137128 268210 137184
rect 239397 137126 268210 137128
rect 239397 137123 239463 137126
rect 264973 137050 265039 137053
rect 264973 137048 268180 137050
rect 264973 136992 264978 137048
rect 265034 136992 268180 137048
rect 264973 136990 268180 136992
rect 264973 136987 265039 136990
rect 231485 136914 231551 136917
rect 228988 136912 231551 136914
rect -960 136778 480 136868
rect 228988 136856 231490 136912
rect 231546 136856 231551 136912
rect 228988 136854 231551 136856
rect 231485 136851 231551 136854
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 181437 136642 181503 136645
rect 188521 136642 188587 136645
rect 181437 136640 188587 136642
rect 181437 136584 181442 136640
rect 181498 136584 188526 136640
rect 188582 136584 188587 136640
rect 181437 136582 188587 136584
rect 181437 136579 181503 136582
rect 188521 136579 188587 136582
rect 215937 136642 216003 136645
rect 282821 136642 282887 136645
rect 215937 136640 217028 136642
rect 215937 136584 215942 136640
rect 215998 136584 217028 136640
rect 279956 136640 282887 136642
rect 215937 136582 217028 136584
rect 215937 136579 216003 136582
rect 231761 136370 231827 136373
rect 268150 136370 268210 136612
rect 279956 136584 282826 136640
rect 282882 136584 282887 136640
rect 279956 136582 282887 136584
rect 282821 136579 282887 136582
rect 228988 136368 231827 136370
rect 228988 136312 231766 136368
rect 231822 136312 231827 136368
rect 228988 136310 231827 136312
rect 231761 136307 231827 136310
rect 258030 136310 268210 136370
rect 214005 135962 214071 135965
rect 231669 135962 231735 135965
rect 214005 135960 217028 135962
rect 214005 135904 214010 135960
rect 214066 135904 217028 135960
rect 214005 135902 217028 135904
rect 228988 135960 231735 135962
rect 228988 135904 231674 135960
rect 231730 135904 231735 135960
rect 228988 135902 231735 135904
rect 214005 135899 214071 135902
rect 231669 135899 231735 135902
rect 242198 135764 242204 135828
rect 242268 135826 242274 135828
rect 258030 135826 258090 136310
rect 264973 136234 265039 136237
rect 264973 136232 268180 136234
rect 264973 136176 264978 136232
rect 265034 136176 268180 136232
rect 264973 136174 268180 136176
rect 264973 136171 265039 136174
rect 280470 135962 280476 135964
rect 279956 135902 280476 135962
rect 280470 135900 280476 135902
rect 280540 135900 280546 135964
rect 242268 135766 258090 135826
rect 242268 135764 242274 135766
rect 267774 135628 267780 135692
rect 267844 135690 267850 135692
rect 267844 135630 268180 135690
rect 267844 135628 267850 135630
rect 230933 135418 230999 135421
rect 228988 135416 230999 135418
rect 228988 135360 230938 135416
rect 230994 135360 230999 135416
rect 228988 135358 230999 135360
rect 230933 135355 230999 135358
rect 247677 135418 247743 135421
rect 247677 135416 268210 135418
rect 247677 135360 247682 135416
rect 247738 135360 268210 135416
rect 247677 135358 268210 135360
rect 247677 135355 247743 135358
rect 213913 135282 213979 135285
rect 213913 135280 217028 135282
rect 213913 135224 213918 135280
rect 213974 135224 217028 135280
rect 268150 135252 268210 135358
rect 213913 135222 217028 135224
rect 213913 135219 213979 135222
rect 283097 135146 283163 135149
rect 279956 135144 283163 135146
rect 279956 135088 283102 135144
rect 283158 135088 283163 135144
rect 279956 135086 283163 135088
rect 283097 135083 283163 135086
rect 231761 135010 231827 135013
rect 228988 135008 231827 135010
rect 228988 134952 231766 135008
rect 231822 134952 231827 135008
rect 228988 134950 231827 134952
rect 231761 134947 231827 134950
rect 265065 134874 265131 134877
rect 265065 134872 268180 134874
rect 265065 134816 265070 134872
rect 265126 134816 268180 134872
rect 265065 134814 268180 134816
rect 265065 134811 265131 134814
rect 214557 134602 214623 134605
rect 214557 134600 217028 134602
rect 214557 134544 214562 134600
rect 214618 134544 217028 134600
rect 214557 134542 217028 134544
rect 214557 134539 214623 134542
rect 231669 134466 231735 134469
rect 228988 134464 231735 134466
rect 228988 134408 231674 134464
rect 231730 134408 231735 134464
rect 228988 134406 231735 134408
rect 231669 134403 231735 134406
rect 250294 134404 250300 134468
rect 250364 134466 250370 134468
rect 265893 134466 265959 134469
rect 250364 134464 265959 134466
rect 250364 134408 265898 134464
rect 265954 134408 265959 134464
rect 250364 134406 265959 134408
rect 250364 134404 250370 134406
rect 265893 134403 265959 134406
rect 265617 134194 265683 134197
rect 268150 134194 268210 134436
rect 265617 134192 268210 134194
rect 265617 134136 265622 134192
rect 265678 134136 268210 134192
rect 265617 134134 268210 134136
rect 265617 134131 265683 134134
rect 231301 134058 231367 134061
rect 228988 134056 231367 134058
rect 228988 134000 231306 134056
rect 231362 134000 231367 134056
rect 228988 133998 231367 134000
rect 231301 133995 231367 133998
rect 264973 134058 265039 134061
rect 264973 134056 268180 134058
rect 264973 134000 264978 134056
rect 265034 134000 268180 134056
rect 264973 133998 268180 134000
rect 264973 133995 265039 133998
rect 213913 133922 213979 133925
rect 279926 133922 279986 134436
rect 290590 133922 290596 133924
rect 213913 133920 217028 133922
rect 213913 133864 213918 133920
rect 213974 133864 217028 133920
rect 213913 133862 217028 133864
rect 279926 133862 290596 133922
rect 213913 133859 213979 133862
rect 290590 133860 290596 133862
rect 290660 133860 290666 133924
rect 230974 133514 230980 133516
rect 228988 133454 230980 133514
rect 230974 133452 230980 133454
rect 231044 133452 231050 133516
rect 214005 133378 214071 133381
rect 214005 133376 217028 133378
rect 214005 133320 214010 133376
rect 214066 133320 217028 133376
rect 214005 133318 217028 133320
rect 214005 133315 214071 133318
rect 262765 133242 262831 133245
rect 268150 133242 268210 133620
rect 262765 133240 268210 133242
rect 262765 133184 262770 133240
rect 262826 133184 268210 133240
rect 262765 133182 268210 133184
rect 262765 133179 262831 133182
rect 191097 133106 191163 133109
rect 213269 133106 213335 133109
rect 231485 133106 231551 133109
rect 191097 133104 213335 133106
rect 191097 133048 191102 133104
rect 191158 133048 213274 133104
rect 213330 133048 213335 133104
rect 191097 133046 213335 133048
rect 228988 133104 231551 133106
rect 228988 133048 231490 133104
rect 231546 133048 231551 133104
rect 228988 133046 231551 133048
rect 191097 133043 191163 133046
rect 213269 133043 213335 133046
rect 231485 133043 231551 133046
rect 258030 133046 268180 133106
rect 242014 132908 242020 132972
rect 242084 132970 242090 132972
rect 258030 132970 258090 133046
rect 242084 132910 258090 132970
rect 279926 132970 279986 133620
rect 279926 132910 287070 132970
rect 242084 132908 242090 132910
rect 229686 132772 229692 132836
rect 229756 132834 229762 132836
rect 262765 132834 262831 132837
rect 282821 132834 282887 132837
rect 229756 132832 262831 132834
rect 229756 132776 262770 132832
rect 262826 132776 262831 132832
rect 229756 132774 262831 132776
rect 279956 132832 282887 132834
rect 279956 132776 282826 132832
rect 282882 132776 282887 132832
rect 279956 132774 282887 132776
rect 229756 132772 229762 132774
rect 262765 132771 262831 132774
rect 282821 132771 282887 132774
rect 213913 132698 213979 132701
rect 265709 132698 265775 132701
rect 213913 132696 217028 132698
rect 213913 132640 213918 132696
rect 213974 132640 217028 132696
rect 213913 132638 217028 132640
rect 265709 132696 268180 132698
rect 265709 132640 265714 132696
rect 265770 132640 268180 132696
rect 265709 132638 268180 132640
rect 213913 132635 213979 132638
rect 265709 132635 265775 132638
rect 231209 132562 231275 132565
rect 228988 132560 231275 132562
rect 228988 132504 231214 132560
rect 231270 132504 231275 132560
rect 228988 132502 231275 132504
rect 287010 132562 287070 132910
rect 295374 132562 295380 132564
rect 287010 132502 295380 132562
rect 231209 132499 231275 132502
rect 295374 132500 295380 132502
rect 295444 132500 295450 132564
rect 265065 132290 265131 132293
rect 265065 132288 268180 132290
rect 265065 132232 265070 132288
rect 265126 132232 268180 132288
rect 265065 132230 268180 132232
rect 265065 132227 265131 132230
rect 230933 132154 230999 132157
rect 282821 132154 282887 132157
rect 228988 132152 230999 132154
rect 228988 132096 230938 132152
rect 230994 132096 230999 132152
rect 228988 132094 230999 132096
rect 279956 132152 282887 132154
rect 279956 132096 282826 132152
rect 282882 132096 282887 132152
rect 279956 132094 282887 132096
rect 230933 132091 230999 132094
rect 282821 132091 282887 132094
rect 214005 132018 214071 132021
rect 214005 132016 217028 132018
rect 214005 131960 214010 132016
rect 214066 131960 217028 132016
rect 214005 131958 217028 131960
rect 214005 131955 214071 131958
rect 264973 131882 265039 131885
rect 264973 131880 268180 131882
rect 264973 131824 264978 131880
rect 265034 131824 268180 131880
rect 264973 131822 268180 131824
rect 264973 131819 265039 131822
rect 231158 131610 231164 131612
rect 228988 131550 231164 131610
rect 231158 131548 231164 131550
rect 231228 131548 231234 131612
rect 245009 131474 245075 131477
rect 245009 131472 268180 131474
rect 245009 131416 245014 131472
rect 245070 131416 268180 131472
rect 245009 131414 268180 131416
rect 245009 131411 245075 131414
rect 213913 131338 213979 131341
rect 280286 131338 280292 131340
rect 213913 131336 217028 131338
rect 213913 131280 213918 131336
rect 213974 131280 217028 131336
rect 213913 131278 217028 131280
rect 279956 131278 280292 131338
rect 213913 131275 213979 131278
rect 280286 131276 280292 131278
rect 280356 131276 280362 131340
rect 230473 131202 230539 131205
rect 228988 131200 230539 131202
rect 228988 131144 230478 131200
rect 230534 131144 230539 131200
rect 228988 131142 230539 131144
rect 230473 131139 230539 131142
rect 266854 131004 266860 131068
rect 266924 131066 266930 131068
rect 266924 131006 268180 131066
rect 266924 131004 266930 131006
rect 214005 130658 214071 130661
rect 231761 130658 231827 130661
rect 282269 130658 282335 130661
rect 214005 130656 217028 130658
rect 214005 130600 214010 130656
rect 214066 130600 217028 130656
rect 214005 130598 217028 130600
rect 228988 130656 231827 130658
rect 228988 130600 231766 130656
rect 231822 130600 231827 130656
rect 228988 130598 231827 130600
rect 279956 130656 282335 130658
rect 279956 130600 282274 130656
rect 282330 130600 282335 130656
rect 279956 130598 282335 130600
rect 214005 130595 214071 130598
rect 231761 130595 231827 130598
rect 282269 130595 282335 130598
rect 264973 130522 265039 130525
rect 264973 130520 268180 130522
rect 264973 130464 264978 130520
rect 265034 130464 268180 130520
rect 264973 130462 268180 130464
rect 264973 130459 265039 130462
rect 231301 130386 231367 130389
rect 257613 130386 257679 130389
rect 231301 130384 257679 130386
rect 231301 130328 231306 130384
rect 231362 130328 257618 130384
rect 257674 130328 257679 130384
rect 231301 130326 257679 130328
rect 231301 130323 231367 130326
rect 257613 130323 257679 130326
rect 231117 130250 231183 130253
rect 228988 130248 231183 130250
rect 228988 130192 231122 130248
rect 231178 130192 231183 130248
rect 228988 130190 231183 130192
rect 231117 130187 231183 130190
rect 258030 130054 268180 130114
rect 213913 129978 213979 129981
rect 254853 129978 254919 129981
rect 258030 129978 258090 130054
rect 213913 129976 217028 129978
rect 213913 129920 213918 129976
rect 213974 129920 217028 129976
rect 213913 129918 217028 129920
rect 254853 129976 258090 129978
rect 254853 129920 254858 129976
rect 254914 129920 258090 129976
rect 254853 129918 258090 129920
rect 213913 129915 213979 129918
rect 254853 129915 254919 129918
rect 231485 129842 231551 129845
rect 280153 129842 280219 129845
rect 228988 129840 231551 129842
rect 228988 129784 231490 129840
rect 231546 129784 231551 129840
rect 228988 129782 231551 129784
rect 279956 129840 280219 129842
rect 279956 129784 280158 129840
rect 280214 129784 280219 129840
rect 279956 129782 280219 129784
rect 231485 129779 231551 129782
rect 280153 129779 280219 129782
rect 268150 129434 268210 129676
rect 258030 129374 268210 129434
rect 66161 129298 66227 129301
rect 68142 129298 68816 129304
rect 66161 129296 68816 129298
rect 66161 129240 66166 129296
rect 66222 129244 68816 129296
rect 213913 129298 213979 129301
rect 231761 129298 231827 129301
rect 213913 129296 217028 129298
rect 66222 129240 68202 129244
rect 66161 129238 68202 129240
rect 213913 129240 213918 129296
rect 213974 129240 217028 129296
rect 213913 129238 217028 129240
rect 228988 129296 231827 129298
rect 228988 129240 231766 129296
rect 231822 129240 231827 129296
rect 228988 129238 231827 129240
rect 66161 129235 66227 129238
rect 213913 129235 213979 129238
rect 231761 129235 231827 129238
rect 230749 129026 230815 129029
rect 245101 129026 245167 129029
rect 230749 129024 245167 129026
rect 230749 128968 230754 129024
rect 230810 128968 245106 129024
rect 245162 128968 245167 129024
rect 230749 128966 245167 128968
rect 230749 128963 230815 128966
rect 245101 128963 245167 128966
rect 251766 128964 251772 129028
rect 251836 129026 251842 129028
rect 258030 129026 258090 129374
rect 264973 129298 265039 129301
rect 264973 129296 268180 129298
rect 264973 129240 264978 129296
rect 265034 129240 268180 129296
rect 264973 129238 268180 129240
rect 264973 129235 265039 129238
rect 282085 129026 282151 129029
rect 251836 128966 258090 129026
rect 279956 129024 282151 129026
rect 279956 128968 282090 129024
rect 282146 128968 282151 129024
rect 279956 128966 282151 128968
rect 251836 128964 251842 128966
rect 282085 128963 282151 128966
rect 231485 128890 231551 128893
rect 228988 128888 231551 128890
rect 228988 128832 231490 128888
rect 231546 128832 231551 128888
rect 228988 128830 231551 128832
rect 231485 128827 231551 128830
rect 265157 128890 265223 128893
rect 265157 128888 268180 128890
rect 265157 128832 265162 128888
rect 265218 128832 268180 128888
rect 265157 128830 268180 128832
rect 265157 128827 265223 128830
rect 214005 128754 214071 128757
rect 214005 128752 217028 128754
rect 214005 128696 214010 128752
rect 214066 128696 217028 128752
rect 214005 128694 217028 128696
rect 214005 128691 214071 128694
rect 264237 128482 264303 128485
rect 264237 128480 268180 128482
rect 264237 128424 264242 128480
rect 264298 128424 268180 128480
rect 264237 128422 268180 128424
rect 264237 128419 264303 128422
rect 231761 128346 231827 128349
rect 282821 128346 282887 128349
rect 228988 128344 231827 128346
rect 228988 128288 231766 128344
rect 231822 128288 231827 128344
rect 228988 128286 231827 128288
rect 279956 128344 282887 128346
rect 279956 128288 282826 128344
rect 282882 128288 282887 128344
rect 279956 128286 282887 128288
rect 231761 128283 231827 128286
rect 282821 128283 282887 128286
rect 65517 128074 65583 128077
rect 68142 128074 68816 128080
rect 65517 128072 68816 128074
rect 65517 128016 65522 128072
rect 65578 128020 68816 128072
rect 214005 128074 214071 128077
rect 214005 128072 217028 128074
rect 65578 128016 68202 128020
rect 65517 128014 68202 128016
rect 214005 128016 214010 128072
rect 214066 128016 217028 128072
rect 214005 128014 217028 128016
rect 65517 128011 65583 128014
rect 214005 128011 214071 128014
rect 231669 127938 231735 127941
rect 228988 127936 231735 127938
rect 228988 127880 231674 127936
rect 231730 127880 231735 127936
rect 228988 127878 231735 127880
rect 231669 127875 231735 127878
rect 262765 127666 262831 127669
rect 268150 127666 268210 127908
rect 262765 127664 268210 127666
rect 262765 127608 262770 127664
rect 262826 127608 268210 127664
rect 262765 127606 268210 127608
rect 262765 127603 262831 127606
rect 281993 127530 282059 127533
rect 258030 127470 268180 127530
rect 279956 127528 282059 127530
rect 279956 127472 281998 127528
rect 282054 127472 282059 127528
rect 279956 127470 282059 127472
rect 213913 127394 213979 127397
rect 230657 127394 230723 127397
rect 213913 127392 217028 127394
rect 213913 127336 213918 127392
rect 213974 127336 217028 127392
rect 213913 127334 217028 127336
rect 228988 127392 230723 127394
rect 228988 127336 230662 127392
rect 230718 127336 230723 127392
rect 228988 127334 230723 127336
rect 213913 127331 213979 127334
rect 230657 127331 230723 127334
rect 246481 127394 246547 127397
rect 258030 127394 258090 127470
rect 281993 127467 282059 127470
rect 246481 127392 258090 127394
rect 246481 127336 246486 127392
rect 246542 127336 258090 127392
rect 246481 127334 258090 127336
rect 246481 127331 246547 127334
rect 255814 127196 255820 127260
rect 255884 127258 255890 127260
rect 262765 127258 262831 127261
rect 255884 127256 262831 127258
rect 255884 127200 262770 127256
rect 262826 127200 262831 127256
rect 255884 127198 262831 127200
rect 255884 127196 255890 127198
rect 262765 127195 262831 127198
rect 264094 127060 264100 127124
rect 264164 127122 264170 127124
rect 264164 127062 268180 127122
rect 264164 127060 264170 127062
rect 230749 126986 230815 126989
rect 228988 126984 230815 126986
rect 228988 126928 230754 126984
rect 230810 126928 230815 126984
rect 228988 126926 230815 126928
rect 230749 126923 230815 126926
rect 214741 126714 214807 126717
rect 214741 126712 217028 126714
rect 214741 126656 214746 126712
rect 214802 126656 217028 126712
rect 214741 126654 217028 126656
rect 214741 126651 214807 126654
rect 232773 126442 232839 126445
rect 268150 126442 268210 126684
rect 228988 126440 232839 126442
rect 228988 126384 232778 126440
rect 232834 126384 232839 126440
rect 228988 126382 232839 126384
rect 232773 126379 232839 126382
rect 258030 126382 268210 126442
rect 67633 126306 67699 126309
rect 68142 126306 68816 126312
rect 67633 126304 68816 126306
rect 67633 126248 67638 126304
rect 67694 126252 68816 126304
rect 174813 126306 174879 126309
rect 214005 126306 214071 126309
rect 174813 126304 214071 126306
rect 67694 126248 68202 126252
rect 67633 126246 68202 126248
rect 174813 126248 174818 126304
rect 174874 126248 214010 126304
rect 214066 126248 214071 126304
rect 174813 126246 214071 126248
rect 67633 126243 67699 126246
rect 174813 126243 174879 126246
rect 214005 126243 214071 126246
rect 231209 126306 231275 126309
rect 240777 126306 240843 126309
rect 231209 126304 240843 126306
rect 231209 126248 231214 126304
rect 231270 126248 240782 126304
rect 240838 126248 240843 126304
rect 231209 126246 240843 126248
rect 231209 126243 231275 126246
rect 240777 126243 240843 126246
rect 213913 126034 213979 126037
rect 231761 126034 231827 126037
rect 213913 126032 217028 126034
rect 213913 125976 213918 126032
rect 213974 125976 217028 126032
rect 213913 125974 217028 125976
rect 228988 126032 231827 126034
rect 228988 125976 231766 126032
rect 231822 125976 231827 126032
rect 228988 125974 231827 125976
rect 213913 125971 213979 125974
rect 231761 125971 231827 125974
rect 232497 126034 232563 126037
rect 258030 126034 258090 126382
rect 279374 126309 279434 126820
rect 265065 126306 265131 126309
rect 265065 126304 268180 126306
rect 265065 126248 265070 126304
rect 265126 126248 268180 126304
rect 265065 126246 268180 126248
rect 279325 126304 279434 126309
rect 279325 126248 279330 126304
rect 279386 126248 279434 126304
rect 279325 126246 279434 126248
rect 265065 126243 265131 126246
rect 279325 126243 279391 126246
rect 282269 126034 282335 126037
rect 232497 126032 258090 126034
rect 232497 125976 232502 126032
rect 232558 125976 258090 126032
rect 232497 125974 258090 125976
rect 279956 126032 282335 126034
rect 279956 125976 282274 126032
rect 282330 125976 282335 126032
rect 279956 125974 282335 125976
rect 232497 125971 232563 125974
rect 282269 125971 282335 125974
rect 580901 126034 580967 126037
rect 583520 126034 584960 126124
rect 580901 126032 584960 126034
rect 580901 125976 580906 126032
rect 580962 125976 584960 126032
rect 580901 125974 584960 125976
rect 580901 125971 580967 125974
rect 264973 125898 265039 125901
rect 264973 125896 268180 125898
rect 264973 125840 264978 125896
rect 265034 125840 268180 125896
rect 583520 125884 584960 125974
rect 264973 125838 268180 125840
rect 264973 125835 265039 125838
rect 234153 125490 234219 125493
rect 228988 125488 234219 125490
rect 228988 125432 234158 125488
rect 234214 125432 234219 125488
rect 228988 125430 234219 125432
rect 234153 125427 234219 125430
rect 214557 125354 214623 125357
rect 265065 125354 265131 125357
rect 214557 125352 217028 125354
rect 214557 125296 214562 125352
rect 214618 125296 217028 125352
rect 214557 125294 217028 125296
rect 265065 125352 268180 125354
rect 265065 125296 265070 125352
rect 265126 125296 268180 125352
rect 265065 125294 268180 125296
rect 214557 125291 214623 125294
rect 265065 125291 265131 125294
rect 65977 125218 66043 125221
rect 68142 125218 68816 125224
rect 282821 125218 282887 125221
rect 65977 125216 68816 125218
rect 65977 125160 65982 125216
rect 66038 125164 68816 125216
rect 279956 125216 282887 125218
rect 66038 125160 68202 125164
rect 65977 125158 68202 125160
rect 279956 125160 282826 125216
rect 282882 125160 282887 125216
rect 279956 125158 282887 125160
rect 65977 125155 66043 125158
rect 282821 125155 282887 125158
rect 231301 125082 231367 125085
rect 228988 125080 231367 125082
rect 228988 125024 231306 125080
rect 231362 125024 231367 125080
rect 228988 125022 231367 125024
rect 231301 125019 231367 125022
rect 213913 124674 213979 124677
rect 235441 124674 235507 124677
rect 268150 124674 268210 124916
rect 213913 124672 217028 124674
rect 213913 124616 213918 124672
rect 213974 124616 217028 124672
rect 213913 124614 217028 124616
rect 235441 124672 268210 124674
rect 235441 124616 235446 124672
rect 235502 124616 268210 124672
rect 235441 124614 268210 124616
rect 213913 124611 213979 124614
rect 235441 124611 235507 124614
rect 232865 124538 232931 124541
rect 228988 124536 232931 124538
rect 228988 124480 232870 124536
rect 232926 124480 232931 124536
rect 228988 124478 232931 124480
rect 232865 124475 232931 124478
rect 264973 124538 265039 124541
rect 282729 124538 282795 124541
rect 264973 124536 268180 124538
rect 264973 124480 264978 124536
rect 265034 124480 268180 124536
rect 264973 124478 268180 124480
rect 279956 124536 282795 124538
rect 279956 124480 282734 124536
rect 282790 124480 282795 124536
rect 279956 124478 282795 124480
rect 264973 124475 265039 124478
rect 282729 124475 282795 124478
rect 214005 124130 214071 124133
rect 251817 124130 251883 124133
rect 214005 124128 217028 124130
rect 214005 124072 214010 124128
rect 214066 124072 217028 124128
rect 214005 124070 217028 124072
rect 228988 124128 251883 124130
rect 228988 124072 251822 124128
rect 251878 124072 251883 124128
rect 228988 124070 251883 124072
rect 214005 124067 214071 124070
rect 251817 124067 251883 124070
rect 264973 124130 265039 124133
rect 264973 124128 268180 124130
rect 264973 124072 264978 124128
rect 265034 124072 268180 124128
rect 264973 124070 268180 124072
rect 264973 124067 265039 124070
rect -960 123572 480 123812
rect 267641 123722 267707 123725
rect 282821 123722 282887 123725
rect 267641 123720 268180 123722
rect 267641 123664 267646 123720
rect 267702 123664 268180 123720
rect 267641 123662 268180 123664
rect 279956 123720 282887 123722
rect 279956 123664 282826 123720
rect 282882 123664 282887 123720
rect 279956 123662 282887 123664
rect 267641 123659 267707 123662
rect 282821 123659 282887 123662
rect 67449 123586 67515 123589
rect 68142 123586 68816 123592
rect 231761 123586 231827 123589
rect 67449 123584 68816 123586
rect 67449 123528 67454 123584
rect 67510 123532 68816 123584
rect 228988 123584 231827 123586
rect 67510 123528 68202 123532
rect 67449 123526 68202 123528
rect 228988 123528 231766 123584
rect 231822 123528 231827 123584
rect 228988 123526 231827 123528
rect 67449 123523 67515 123526
rect 231761 123523 231827 123526
rect 213913 123450 213979 123453
rect 213913 123448 217028 123450
rect 213913 123392 213918 123448
rect 213974 123392 217028 123448
rect 213913 123390 217028 123392
rect 213913 123387 213979 123390
rect 258030 123254 268180 123314
rect 230933 123178 230999 123181
rect 228988 123176 230999 123178
rect 228988 123120 230938 123176
rect 230994 123120 230999 123176
rect 228988 123118 230999 123120
rect 230933 123115 230999 123118
rect 243813 123178 243879 123181
rect 258030 123178 258090 123254
rect 243813 123176 258090 123178
rect 243813 123120 243818 123176
rect 243874 123120 258090 123176
rect 243813 123118 258090 123120
rect 243813 123115 243879 123118
rect 258809 123042 258875 123045
rect 282269 123042 282335 123045
rect 258809 123040 268210 123042
rect 258809 122984 258814 123040
rect 258870 122984 268210 123040
rect 258809 122982 268210 122984
rect 279956 123040 282335 123042
rect 279956 122984 282274 123040
rect 282330 122984 282335 123040
rect 279956 122982 282335 122984
rect 258809 122979 258875 122982
rect 268150 122876 268210 122982
rect 282269 122979 282335 122982
rect 213913 122770 213979 122773
rect 264513 122770 264579 122773
rect 213913 122768 217028 122770
rect 213913 122712 213918 122768
rect 213974 122712 217028 122768
rect 213913 122710 217028 122712
rect 238710 122768 264579 122770
rect 238710 122712 264518 122768
rect 264574 122712 264579 122768
rect 238710 122710 264579 122712
rect 213913 122707 213979 122710
rect 66069 122634 66135 122637
rect 68142 122634 68816 122640
rect 238710 122634 238770 122710
rect 264513 122707 264579 122710
rect 66069 122632 68816 122634
rect 66069 122576 66074 122632
rect 66130 122580 68816 122632
rect 66130 122576 68202 122580
rect 66069 122574 68202 122576
rect 228988 122574 238770 122634
rect 66069 122571 66135 122574
rect 264973 122362 265039 122365
rect 264973 122360 268180 122362
rect 264973 122304 264978 122360
rect 265034 122304 268180 122360
rect 264973 122302 268180 122304
rect 264973 122299 265039 122302
rect 230749 122226 230815 122229
rect 282821 122226 282887 122229
rect 228988 122224 230815 122226
rect 228988 122168 230754 122224
rect 230810 122168 230815 122224
rect 228988 122166 230815 122168
rect 279956 122224 282887 122226
rect 279956 122168 282826 122224
rect 282882 122168 282887 122224
rect 279956 122166 282887 122168
rect 230749 122163 230815 122166
rect 282821 122163 282887 122166
rect 213361 122090 213427 122093
rect 213361 122088 217028 122090
rect 213361 122032 213366 122088
rect 213422 122032 217028 122088
rect 213361 122030 217028 122032
rect 213361 122027 213427 122030
rect 258030 121894 268180 121954
rect 232773 121818 232839 121821
rect 258030 121818 258090 121894
rect 232773 121816 258090 121818
rect 232773 121760 232778 121816
rect 232834 121760 258090 121816
rect 232773 121758 258090 121760
rect 232773 121755 232839 121758
rect 231577 121682 231643 121685
rect 228988 121680 231643 121682
rect 228988 121624 231582 121680
rect 231638 121624 231643 121680
rect 228988 121622 231643 121624
rect 231577 121619 231643 121622
rect 264605 121546 264671 121549
rect 264605 121544 268180 121546
rect 264605 121488 264610 121544
rect 264666 121488 268180 121544
rect 264605 121486 268180 121488
rect 264605 121483 264671 121486
rect 214005 121410 214071 121413
rect 282821 121410 282887 121413
rect 214005 121408 217028 121410
rect 214005 121352 214010 121408
rect 214066 121352 217028 121408
rect 214005 121350 217028 121352
rect 279956 121408 282887 121410
rect 279956 121352 282826 121408
rect 282882 121352 282887 121408
rect 279956 121350 282887 121352
rect 214005 121347 214071 121350
rect 282821 121347 282887 121350
rect 231761 121274 231827 121277
rect 228988 121272 231827 121274
rect 228988 121216 231766 121272
rect 231822 121216 231827 121272
rect 228988 121214 231827 121216
rect 231761 121211 231827 121214
rect 67725 120866 67791 120869
rect 68142 120866 68816 120872
rect 67725 120864 68816 120866
rect 67725 120808 67730 120864
rect 67786 120812 68816 120864
rect 67786 120808 68202 120812
rect 67725 120806 68202 120808
rect 67725 120803 67791 120806
rect 240726 120804 240732 120868
rect 240796 120866 240802 120868
rect 268150 120866 268210 121108
rect 240796 120806 268210 120866
rect 240796 120804 240802 120806
rect 213913 120730 213979 120733
rect 231209 120730 231275 120733
rect 282821 120730 282887 120733
rect 213913 120728 217028 120730
rect 213913 120672 213918 120728
rect 213974 120672 217028 120728
rect 213913 120670 217028 120672
rect 228988 120728 231275 120730
rect 228988 120672 231214 120728
rect 231270 120672 231275 120728
rect 279956 120728 282887 120730
rect 228988 120670 231275 120672
rect 213913 120667 213979 120670
rect 231209 120667 231275 120670
rect 229829 120458 229895 120461
rect 268150 120458 268210 120700
rect 279956 120672 282826 120728
rect 282882 120672 282887 120728
rect 279956 120670 282887 120672
rect 282821 120667 282887 120670
rect 229829 120456 268210 120458
rect 229829 120400 229834 120456
rect 229890 120400 268210 120456
rect 229829 120398 268210 120400
rect 229829 120395 229895 120398
rect 231669 120322 231735 120325
rect 228988 120320 231735 120322
rect 228988 120264 231674 120320
rect 231730 120264 231735 120320
rect 228988 120262 231735 120264
rect 231669 120259 231735 120262
rect 264973 120322 265039 120325
rect 264973 120320 268180 120322
rect 264973 120264 264978 120320
rect 265034 120264 268180 120320
rect 264973 120262 268180 120264
rect 264973 120259 265039 120262
rect 214005 120050 214071 120053
rect 253197 120050 253263 120053
rect 214005 120048 217028 120050
rect 214005 119992 214010 120048
rect 214066 119992 217028 120048
rect 214005 119990 217028 119992
rect 238710 120048 253263 120050
rect 238710 119992 253202 120048
rect 253258 119992 253263 120048
rect 238710 119990 253263 119992
rect 214005 119987 214071 119990
rect 238710 119778 238770 119990
rect 253197 119987 253263 119990
rect 282821 119914 282887 119917
rect 279956 119912 282887 119914
rect 279956 119856 282826 119912
rect 282882 119856 282887 119912
rect 279956 119854 282887 119856
rect 282821 119851 282887 119854
rect 228988 119718 238770 119778
rect 264973 119778 265039 119781
rect 264973 119776 268180 119778
rect 264973 119720 264978 119776
rect 265034 119720 268180 119776
rect 264973 119718 268180 119720
rect 264973 119715 265039 119718
rect 213913 119506 213979 119509
rect 213913 119504 217028 119506
rect 213913 119448 213918 119504
rect 213974 119448 217028 119504
rect 213913 119446 217028 119448
rect 213913 119443 213979 119446
rect 231761 119370 231827 119373
rect 228988 119368 231827 119370
rect 228988 119312 231766 119368
rect 231822 119312 231827 119368
rect 228988 119310 231827 119312
rect 231761 119307 231827 119310
rect 238017 119098 238083 119101
rect 268150 119098 268210 119340
rect 282729 119234 282795 119237
rect 279956 119232 282795 119234
rect 279956 119176 282734 119232
rect 282790 119176 282795 119232
rect 279956 119174 282795 119176
rect 282729 119171 282795 119174
rect 238017 119096 268210 119098
rect 238017 119040 238022 119096
rect 238078 119040 268210 119096
rect 238017 119038 268210 119040
rect 238017 119035 238083 119038
rect 230657 118962 230723 118965
rect 228988 118960 230723 118962
rect 228988 118904 230662 118960
rect 230718 118904 230723 118960
rect 228988 118902 230723 118904
rect 230657 118899 230723 118902
rect 265433 118962 265499 118965
rect 265433 118960 268180 118962
rect 265433 118904 265438 118960
rect 265494 118904 268180 118960
rect 265433 118902 268180 118904
rect 265433 118899 265499 118902
rect 189901 118826 189967 118829
rect 189901 118824 217028 118826
rect 189901 118768 189906 118824
rect 189962 118768 217028 118824
rect 189901 118766 217028 118768
rect 189901 118763 189967 118766
rect 233877 118418 233943 118421
rect 228988 118416 233943 118418
rect 228988 118360 233882 118416
rect 233938 118360 233943 118416
rect 228988 118358 233943 118360
rect 233877 118355 233943 118358
rect 268150 118282 268210 118524
rect 282821 118418 282887 118421
rect 279956 118416 282887 118418
rect 279956 118360 282826 118416
rect 282882 118360 282887 118416
rect 279956 118358 282887 118360
rect 282821 118355 282887 118358
rect 258030 118222 268210 118282
rect 214005 118146 214071 118149
rect 214005 118144 217028 118146
rect 214005 118088 214010 118144
rect 214066 118088 217028 118144
rect 214005 118086 217028 118088
rect 214005 118083 214071 118086
rect 231393 118010 231459 118013
rect 228988 118008 231459 118010
rect 228988 117952 231398 118008
rect 231454 117952 231459 118008
rect 228988 117950 231459 117952
rect 231393 117947 231459 117950
rect 234153 117874 234219 117877
rect 258030 117874 258090 118222
rect 265065 118146 265131 118149
rect 265065 118144 268180 118146
rect 265065 118088 265070 118144
rect 265126 118088 268180 118144
rect 265065 118086 268180 118088
rect 265065 118083 265131 118086
rect 234153 117872 258090 117874
rect 234153 117816 234158 117872
rect 234214 117816 258090 117872
rect 234153 117814 258090 117816
rect 234153 117811 234219 117814
rect 264973 117738 265039 117741
rect 264973 117736 268180 117738
rect 264973 117680 264978 117736
rect 265034 117680 268180 117736
rect 264973 117678 268180 117680
rect 264973 117675 265039 117678
rect 282269 117602 282335 117605
rect 279956 117600 282335 117602
rect 279956 117544 282274 117600
rect 282330 117544 282335 117600
rect 279956 117542 282335 117544
rect 282269 117539 282335 117542
rect 213913 117466 213979 117469
rect 231485 117466 231551 117469
rect 213913 117464 217028 117466
rect 213913 117408 213918 117464
rect 213974 117408 217028 117464
rect 213913 117406 217028 117408
rect 228988 117464 231551 117466
rect 228988 117408 231490 117464
rect 231546 117408 231551 117464
rect 228988 117406 231551 117408
rect 213913 117403 213979 117406
rect 231485 117403 231551 117406
rect 266997 117194 267063 117197
rect 266997 117192 268180 117194
rect 266997 117136 267002 117192
rect 267058 117136 268180 117192
rect 266997 117134 268180 117136
rect 266997 117131 267063 117134
rect 231761 117058 231827 117061
rect 228988 117056 231827 117058
rect 228988 117000 231766 117056
rect 231822 117000 231827 117056
rect 228988 116998 231827 117000
rect 231761 116995 231827 116998
rect 284518 116922 284524 116924
rect 279956 116862 284524 116922
rect 284518 116860 284524 116862
rect 284588 116860 284594 116924
rect 214005 116786 214071 116789
rect 265065 116786 265131 116789
rect 214005 116784 217028 116786
rect 214005 116728 214010 116784
rect 214066 116728 217028 116784
rect 214005 116726 217028 116728
rect 265065 116784 268180 116786
rect 265065 116728 265070 116784
rect 265126 116728 268180 116784
rect 265065 116726 268180 116728
rect 214005 116723 214071 116726
rect 265065 116723 265131 116726
rect 176009 116514 176075 116517
rect 214557 116514 214623 116517
rect 231669 116514 231735 116517
rect 176009 116512 214623 116514
rect 176009 116456 176014 116512
rect 176070 116456 214562 116512
rect 214618 116456 214623 116512
rect 176009 116454 214623 116456
rect 228988 116512 231735 116514
rect 228988 116456 231674 116512
rect 231730 116456 231735 116512
rect 228988 116454 231735 116456
rect 176009 116451 176075 116454
rect 214557 116451 214623 116454
rect 231669 116451 231735 116454
rect 258030 116318 268180 116378
rect 233877 116242 233943 116245
rect 258030 116242 258090 116318
rect 233877 116240 258090 116242
rect 233877 116184 233882 116240
rect 233938 116184 258090 116240
rect 233877 116182 258090 116184
rect 233877 116179 233943 116182
rect 213913 116106 213979 116109
rect 230841 116106 230907 116109
rect 282821 116106 282887 116109
rect 213913 116104 217028 116106
rect 213913 116048 213918 116104
rect 213974 116048 217028 116104
rect 213913 116046 217028 116048
rect 228988 116104 230907 116106
rect 228988 116048 230846 116104
rect 230902 116048 230907 116104
rect 228988 116046 230907 116048
rect 279956 116104 282887 116106
rect 279956 116048 282826 116104
rect 282882 116048 282887 116104
rect 279956 116046 282887 116048
rect 213913 116043 213979 116046
rect 230841 116043 230907 116046
rect 282821 116043 282887 116046
rect 264973 115970 265039 115973
rect 264973 115968 268180 115970
rect 264973 115912 264978 115968
rect 265034 115912 268180 115968
rect 264973 115910 268180 115912
rect 264973 115907 265039 115910
rect 250437 115834 250503 115837
rect 238710 115832 250503 115834
rect 238710 115776 250442 115832
rect 250498 115776 250503 115832
rect 238710 115774 250503 115776
rect 238710 115562 238770 115774
rect 250437 115771 250503 115774
rect 228988 115502 238770 115562
rect 264973 115562 265039 115565
rect 264973 115560 268180 115562
rect 264973 115504 264978 115560
rect 265034 115504 268180 115560
rect 264973 115502 268180 115504
rect 264973 115499 265039 115502
rect 214005 115426 214071 115429
rect 282821 115426 282887 115429
rect 214005 115424 217028 115426
rect 214005 115368 214010 115424
rect 214066 115368 217028 115424
rect 214005 115366 217028 115368
rect 279956 115424 282887 115426
rect 279956 115368 282826 115424
rect 282882 115368 282887 115424
rect 279956 115366 282887 115368
rect 214005 115363 214071 115366
rect 282821 115363 282887 115366
rect 182909 115154 182975 115157
rect 205081 115154 205147 115157
rect 231485 115154 231551 115157
rect 182909 115152 205147 115154
rect 182909 115096 182914 115152
rect 182970 115096 205086 115152
rect 205142 115096 205147 115152
rect 182909 115094 205147 115096
rect 228988 115152 231551 115154
rect 228988 115096 231490 115152
rect 231546 115096 231551 115152
rect 228988 115094 231551 115096
rect 182909 115091 182975 115094
rect 205081 115091 205147 115094
rect 231485 115091 231551 115094
rect 213913 114882 213979 114885
rect 235257 114882 235323 114885
rect 268150 114882 268210 115124
rect 213913 114880 217028 114882
rect 213913 114824 213918 114880
rect 213974 114824 217028 114880
rect 213913 114822 217028 114824
rect 235257 114880 268210 114882
rect 235257 114824 235262 114880
rect 235318 114824 268210 114880
rect 235257 114822 268210 114824
rect 213913 114819 213979 114822
rect 235257 114819 235323 114822
rect 258073 114746 258139 114749
rect 258073 114744 268210 114746
rect 258073 114688 258078 114744
rect 258134 114688 268210 114744
rect 258073 114686 268210 114688
rect 258073 114683 258139 114686
rect 231117 114610 231183 114613
rect 228988 114608 231183 114610
rect 228988 114552 231122 114608
rect 231178 114552 231183 114608
rect 268150 114580 268210 114686
rect 282361 114610 282427 114613
rect 279956 114608 282427 114610
rect 228988 114550 231183 114552
rect 279956 114552 282366 114608
rect 282422 114552 282427 114608
rect 279956 114550 282427 114552
rect 231117 114547 231183 114550
rect 282361 114547 282427 114550
rect 213913 114202 213979 114205
rect 231761 114202 231827 114205
rect 213913 114200 217028 114202
rect 213913 114144 213918 114200
rect 213974 114144 217028 114200
rect 213913 114142 217028 114144
rect 228988 114200 231827 114202
rect 228988 114144 231766 114200
rect 231822 114144 231827 114200
rect 228988 114142 231827 114144
rect 213913 114139 213979 114142
rect 231761 114139 231827 114142
rect 264973 114202 265039 114205
rect 264973 114200 268180 114202
rect 264973 114144 264978 114200
rect 265034 114144 268180 114200
rect 264973 114142 268180 114144
rect 264973 114139 265039 114142
rect 189717 113794 189783 113797
rect 215937 113794 216003 113797
rect 189717 113792 216003 113794
rect 189717 113736 189722 113792
rect 189778 113736 215942 113792
rect 215998 113736 216003 113792
rect 189717 113734 216003 113736
rect 189717 113731 189783 113734
rect 215937 113731 216003 113734
rect 230841 113794 230907 113797
rect 261477 113794 261543 113797
rect 230841 113792 261543 113794
rect 230841 113736 230846 113792
rect 230902 113736 261482 113792
rect 261538 113736 261543 113792
rect 230841 113734 261543 113736
rect 230841 113731 230907 113734
rect 261477 113731 261543 113734
rect 262806 113732 262812 113796
rect 262876 113794 262882 113796
rect 282085 113794 282151 113797
rect 262876 113734 268180 113794
rect 279956 113792 282151 113794
rect 279956 113736 282090 113792
rect 282146 113736 282151 113792
rect 279956 113734 282151 113736
rect 262876 113732 262882 113734
rect 282085 113731 282151 113734
rect 230565 113658 230631 113661
rect 228988 113656 230631 113658
rect 228988 113600 230570 113656
rect 230626 113600 230631 113656
rect 228988 113598 230631 113600
rect 230565 113595 230631 113598
rect 214281 113522 214347 113525
rect 214281 113520 217028 113522
rect 214281 113464 214286 113520
rect 214342 113464 217028 113520
rect 214281 113462 217028 113464
rect 214281 113459 214347 113462
rect 258030 113326 268180 113386
rect 231485 113250 231551 113253
rect 228988 113248 231551 113250
rect 228988 113192 231490 113248
rect 231546 113192 231551 113248
rect 228988 113190 231551 113192
rect 231485 113187 231551 113190
rect 250437 113250 250503 113253
rect 258030 113250 258090 113326
rect 250437 113248 258090 113250
rect 250437 113192 250442 113248
rect 250498 113192 258090 113248
rect 250437 113190 258090 113192
rect 250437 113187 250503 113190
rect 282453 113114 282519 113117
rect 279956 113112 282519 113114
rect 279956 113056 282458 113112
rect 282514 113056 282519 113112
rect 279956 113054 282519 113056
rect 282453 113051 282519 113054
rect 213913 112842 213979 112845
rect 213913 112840 217028 112842
rect 213913 112784 213918 112840
rect 213974 112784 217028 112840
rect 213913 112782 217028 112784
rect 213913 112779 213979 112782
rect 231761 112706 231827 112709
rect 268150 112706 268210 112948
rect 582925 112842 582991 112845
rect 583520 112842 584960 112932
rect 582925 112840 584960 112842
rect 582925 112784 582930 112840
rect 582986 112784 584960 112840
rect 582925 112782 584960 112784
rect 582925 112779 582991 112782
rect 228988 112704 231827 112706
rect 228988 112648 231766 112704
rect 231822 112648 231827 112704
rect 228988 112646 231827 112648
rect 231761 112643 231827 112646
rect 258030 112646 268210 112706
rect 583520 112692 584960 112782
rect 231393 112298 231459 112301
rect 228988 112296 231459 112298
rect 228988 112240 231398 112296
rect 231454 112240 231459 112296
rect 228988 112238 231459 112240
rect 231393 112235 231459 112238
rect 239489 112162 239555 112165
rect 258030 112162 258090 112646
rect 264973 112570 265039 112573
rect 264973 112568 268180 112570
rect 264973 112512 264978 112568
rect 265034 112512 268180 112568
rect 264973 112510 268180 112512
rect 264973 112507 265039 112510
rect 282821 112298 282887 112301
rect 279956 112296 282887 112298
rect 279956 112240 282826 112296
rect 282882 112240 282887 112296
rect 279956 112238 282887 112240
rect 282821 112235 282887 112238
rect 239489 112160 258090 112162
rect 166441 112026 166507 112029
rect 216998 112026 217058 112132
rect 239489 112104 239494 112160
rect 239550 112104 258090 112160
rect 239489 112102 258090 112104
rect 239489 112099 239555 112102
rect 166441 112024 217058 112026
rect 166441 111968 166446 112024
rect 166502 111968 217058 112024
rect 166441 111966 217058 111968
rect 250621 112026 250687 112029
rect 250621 112024 268180 112026
rect 250621 111968 250626 112024
rect 250682 111968 268180 112024
rect 250621 111966 268180 111968
rect 166441 111963 166507 111966
rect 250621 111963 250687 111966
rect 164724 111754 165354 111760
rect 167821 111754 167887 111757
rect 239581 111754 239647 111757
rect 164724 111752 167887 111754
rect 164724 111700 167826 111752
rect 165294 111696 167826 111700
rect 167882 111696 167887 111752
rect 165294 111694 167887 111696
rect 228988 111752 239647 111754
rect 228988 111696 239586 111752
rect 239642 111696 239647 111752
rect 228988 111694 239647 111696
rect 167821 111691 167887 111694
rect 239581 111691 239647 111694
rect 264973 111618 265039 111621
rect 281717 111618 281783 111621
rect 264973 111616 268180 111618
rect 264973 111560 264978 111616
rect 265034 111560 268180 111616
rect 264973 111558 268180 111560
rect 279956 111616 281783 111618
rect 279956 111560 281722 111616
rect 281778 111560 281783 111616
rect 279956 111558 281783 111560
rect 264973 111555 265039 111558
rect 281717 111555 281783 111558
rect 214005 111482 214071 111485
rect 214005 111480 217028 111482
rect 214005 111424 214010 111480
rect 214066 111424 217028 111480
rect 214005 111422 217028 111424
rect 214005 111419 214071 111422
rect 231209 111346 231275 111349
rect 228988 111344 231275 111346
rect 228988 111288 231214 111344
rect 231270 111288 231275 111344
rect 228988 111286 231275 111288
rect 231209 111283 231275 111286
rect 230974 111148 230980 111212
rect 231044 111210 231050 111212
rect 243629 111210 243695 111213
rect 231044 111208 243695 111210
rect 231044 111152 243634 111208
rect 243690 111152 243695 111208
rect 231044 111150 243695 111152
rect 231044 111148 231050 111150
rect 243629 111147 243695 111150
rect 265065 111210 265131 111213
rect 265065 111208 268180 111210
rect 265065 111152 265070 111208
rect 265126 111152 268180 111208
rect 265065 111150 268180 111152
rect 265065 111147 265131 111150
rect 231485 111074 231551 111077
rect 260189 111074 260255 111077
rect 231485 111072 260255 111074
rect 231485 111016 231490 111072
rect 231546 111016 260194 111072
rect 260250 111016 260255 111072
rect 231485 111014 260255 111016
rect 231485 111011 231551 111014
rect 260189 111011 260255 111014
rect 213913 110802 213979 110805
rect 230749 110802 230815 110805
rect 213913 110800 217028 110802
rect -960 110666 480 110756
rect 213913 110744 213918 110800
rect 213974 110744 217028 110800
rect 213913 110742 217028 110744
rect 228988 110800 230815 110802
rect 228988 110744 230754 110800
rect 230810 110744 230815 110800
rect 228988 110742 230815 110744
rect 213913 110739 213979 110742
rect 230749 110739 230815 110742
rect 264329 110802 264395 110805
rect 282821 110802 282887 110805
rect 264329 110800 268180 110802
rect 264329 110744 264334 110800
rect 264390 110744 268180 110800
rect 264329 110742 268180 110744
rect 279956 110800 282887 110802
rect 279956 110744 282826 110800
rect 282882 110744 282887 110800
rect 279956 110742 282887 110744
rect 264329 110739 264395 110742
rect 282821 110739 282887 110742
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 231761 110394 231827 110397
rect 228988 110392 231827 110394
rect 228988 110336 231766 110392
rect 231822 110336 231827 110392
rect 228988 110334 231827 110336
rect 231761 110331 231827 110334
rect 254669 110394 254735 110397
rect 258073 110394 258139 110397
rect 254669 110392 258139 110394
rect 254669 110336 254674 110392
rect 254730 110336 258078 110392
rect 258134 110336 258139 110392
rect 254669 110334 258139 110336
rect 254669 110331 254735 110334
rect 258073 110331 258139 110334
rect 265065 110394 265131 110397
rect 265065 110392 268180 110394
rect 265065 110336 265070 110392
rect 265126 110336 268180 110392
rect 265065 110334 268180 110336
rect 265065 110331 265131 110334
rect 214005 110258 214071 110261
rect 214005 110256 217028 110258
rect 214005 110200 214010 110256
rect 214066 110200 217028 110256
rect 214005 110198 217028 110200
rect 214005 110195 214071 110198
rect 164724 110122 165354 110128
rect 168281 110122 168347 110125
rect 164724 110120 168347 110122
rect 164724 110068 168286 110120
rect 165294 110064 168286 110068
rect 168342 110064 168347 110120
rect 165294 110062 168347 110064
rect 168281 110059 168347 110062
rect 267733 109986 267799 109989
rect 282821 109986 282887 109989
rect 267733 109984 268180 109986
rect 267733 109928 267738 109984
rect 267794 109928 268180 109984
rect 267733 109926 268180 109928
rect 279956 109984 282887 109986
rect 279956 109928 282826 109984
rect 282882 109928 282887 109984
rect 279956 109926 282887 109928
rect 267733 109923 267799 109926
rect 282821 109923 282887 109926
rect 231485 109850 231551 109853
rect 228988 109848 231551 109850
rect 228988 109792 231490 109848
rect 231546 109792 231551 109848
rect 228988 109790 231551 109792
rect 231485 109787 231551 109790
rect 249241 109850 249307 109853
rect 261753 109850 261819 109853
rect 249241 109848 261819 109850
rect 249241 109792 249246 109848
rect 249302 109792 261758 109848
rect 261814 109792 261819 109848
rect 249241 109790 261819 109792
rect 249241 109787 249307 109790
rect 261753 109787 261819 109790
rect 232681 109714 232747 109717
rect 253381 109714 253447 109717
rect 232681 109712 253447 109714
rect 232681 109656 232686 109712
rect 232742 109656 253386 109712
rect 253442 109656 253447 109712
rect 232681 109654 253447 109656
rect 232681 109651 232747 109654
rect 253381 109651 253447 109654
rect 213913 109578 213979 109581
rect 264973 109578 265039 109581
rect 213913 109576 217028 109578
rect 213913 109520 213918 109576
rect 213974 109520 217028 109576
rect 213913 109518 217028 109520
rect 264973 109576 268180 109578
rect 264973 109520 264978 109576
rect 265034 109520 268180 109576
rect 264973 109518 268180 109520
rect 213913 109515 213979 109518
rect 264973 109515 265039 109518
rect 230841 109442 230907 109445
rect 228988 109440 230907 109442
rect 228988 109384 230846 109440
rect 230902 109384 230907 109440
rect 228988 109382 230907 109384
rect 230841 109379 230907 109382
rect 282269 109306 282335 109309
rect 279956 109304 282335 109306
rect 279956 109248 282274 109304
rect 282330 109248 282335 109304
rect 279956 109246 282335 109248
rect 282269 109243 282335 109246
rect 252093 109034 252159 109037
rect 238710 109032 252159 109034
rect 238710 108976 252098 109032
rect 252154 108976 252159 109032
rect 238710 108974 252159 108976
rect 214005 108898 214071 108901
rect 238710 108898 238770 108974
rect 252093 108971 252159 108974
rect 265065 109034 265131 109037
rect 265065 109032 268180 109034
rect 265065 108976 265070 109032
rect 265126 108976 268180 109032
rect 265065 108974 268180 108976
rect 265065 108971 265131 108974
rect 214005 108896 217028 108898
rect 214005 108840 214010 108896
rect 214066 108840 217028 108896
rect 214005 108838 217028 108840
rect 228988 108838 238770 108898
rect 214005 108835 214071 108838
rect 164724 108762 165354 108768
rect 168005 108762 168071 108765
rect 164724 108760 168071 108762
rect 164724 108708 168010 108760
rect 165294 108704 168010 108708
rect 168066 108704 168071 108760
rect 165294 108702 168071 108704
rect 168005 108699 168071 108702
rect 264973 108626 265039 108629
rect 264973 108624 268180 108626
rect 264973 108568 264978 108624
rect 265034 108568 268180 108624
rect 264973 108566 268180 108568
rect 264973 108563 265039 108566
rect 231761 108490 231827 108493
rect 282821 108490 282887 108493
rect 228988 108488 231827 108490
rect 228988 108432 231766 108488
rect 231822 108432 231827 108488
rect 228988 108430 231827 108432
rect 279956 108488 282887 108490
rect 279956 108432 282826 108488
rect 282882 108432 282887 108488
rect 279956 108430 282887 108432
rect 231761 108427 231827 108430
rect 282821 108427 282887 108430
rect 213913 108218 213979 108221
rect 213913 108216 217028 108218
rect 213913 108160 213918 108216
rect 213974 108160 217028 108216
rect 213913 108158 217028 108160
rect 213913 108155 213979 108158
rect 231577 107946 231643 107949
rect 228988 107944 231643 107946
rect 228988 107888 231582 107944
rect 231638 107888 231643 107944
rect 228988 107886 231643 107888
rect 231577 107883 231643 107886
rect 251909 107946 251975 107949
rect 268150 107946 268210 108188
rect 251909 107944 268210 107946
rect 251909 107888 251914 107944
rect 251970 107888 268210 107944
rect 251909 107886 268210 107888
rect 251909 107883 251975 107886
rect 256325 107810 256391 107813
rect 282361 107810 282427 107813
rect 256325 107808 268180 107810
rect 256325 107752 256330 107808
rect 256386 107752 268180 107808
rect 256325 107750 268180 107752
rect 279956 107808 282427 107810
rect 279956 107752 282366 107808
rect 282422 107752 282427 107808
rect 279956 107750 282427 107752
rect 256325 107747 256391 107750
rect 282361 107747 282427 107750
rect 214005 107538 214071 107541
rect 250294 107538 250300 107540
rect 214005 107536 217028 107538
rect 214005 107480 214010 107536
rect 214066 107480 217028 107536
rect 214005 107478 217028 107480
rect 228988 107478 250300 107538
rect 214005 107475 214071 107478
rect 250294 107476 250300 107478
rect 250364 107476 250370 107540
rect 264973 107402 265039 107405
rect 264973 107400 268180 107402
rect 264973 107344 264978 107400
rect 265034 107344 268180 107400
rect 264973 107342 268180 107344
rect 264973 107339 265039 107342
rect 231301 107130 231367 107133
rect 228988 107128 231367 107130
rect 228988 107072 231306 107128
rect 231362 107072 231367 107128
rect 228988 107070 231367 107072
rect 231301 107067 231367 107070
rect 265065 106994 265131 106997
rect 265065 106992 268180 106994
rect 265065 106936 265070 106992
rect 265126 106936 268180 106992
rect 265065 106934 268180 106936
rect 265065 106931 265131 106934
rect 170581 106858 170647 106861
rect 210601 106858 210667 106861
rect 170581 106856 210667 106858
rect 170581 106800 170586 106856
rect 170642 106800 210606 106856
rect 210662 106800 210667 106856
rect 170581 106798 210667 106800
rect 170581 106795 170647 106798
rect 210601 106795 210667 106798
rect 213913 106858 213979 106861
rect 239581 106858 239647 106861
rect 251766 106858 251772 106860
rect 213913 106856 217028 106858
rect 213913 106800 213918 106856
rect 213974 106800 217028 106856
rect 213913 106798 217028 106800
rect 239581 106856 251772 106858
rect 239581 106800 239586 106856
rect 239642 106800 251772 106856
rect 239581 106798 251772 106800
rect 213913 106795 213979 106798
rect 239581 106795 239647 106798
rect 251766 106796 251772 106798
rect 251836 106796 251842 106860
rect 231761 106586 231827 106589
rect 228988 106584 231827 106586
rect 228988 106528 231766 106584
rect 231822 106528 231827 106584
rect 228988 106526 231827 106528
rect 231761 106523 231827 106526
rect 258030 106390 268180 106450
rect 256049 106314 256115 106317
rect 258030 106314 258090 106390
rect 256049 106312 258090 106314
rect 256049 106256 256054 106312
rect 256110 106256 258090 106312
rect 256049 106254 258090 106256
rect 279926 106314 279986 106964
rect 288566 106314 288572 106316
rect 279926 106254 288572 106314
rect 256049 106251 256115 106254
rect 288566 106252 288572 106254
rect 288636 106252 288642 106316
rect 214005 106178 214071 106181
rect 230473 106178 230539 106181
rect 285806 106178 285812 106180
rect 214005 106176 217028 106178
rect 214005 106120 214010 106176
rect 214066 106120 217028 106176
rect 214005 106118 217028 106120
rect 228988 106176 230539 106178
rect 228988 106120 230478 106176
rect 230534 106120 230539 106176
rect 228988 106118 230539 106120
rect 279956 106118 285812 106178
rect 214005 106115 214071 106118
rect 230473 106115 230539 106118
rect 285806 106116 285812 106118
rect 285876 106116 285882 106180
rect 264973 106042 265039 106045
rect 264973 106040 268180 106042
rect 264973 105984 264978 106040
rect 265034 105984 268180 106040
rect 264973 105982 268180 105984
rect 264973 105979 265039 105982
rect 231393 105634 231459 105637
rect 228988 105632 231459 105634
rect 167913 105498 167979 105501
rect 181529 105498 181595 105501
rect 167913 105496 181595 105498
rect 167913 105440 167918 105496
rect 167974 105440 181534 105496
rect 181590 105440 181595 105496
rect 167913 105438 181595 105440
rect 167913 105435 167979 105438
rect 181529 105435 181595 105438
rect 198089 105226 198155 105229
rect 216998 105226 217058 105604
rect 228988 105576 231398 105632
rect 231454 105576 231459 105632
rect 228988 105574 231459 105576
rect 231393 105571 231459 105574
rect 265065 105634 265131 105637
rect 265065 105632 268180 105634
rect 265065 105576 265070 105632
rect 265126 105576 268180 105632
rect 265065 105574 268180 105576
rect 265065 105571 265131 105574
rect 231209 105498 231275 105501
rect 256233 105498 256299 105501
rect 282821 105498 282887 105501
rect 231209 105496 256299 105498
rect 231209 105440 231214 105496
rect 231270 105440 256238 105496
rect 256294 105440 256299 105496
rect 231209 105438 256299 105440
rect 279956 105496 282887 105498
rect 279956 105440 282826 105496
rect 282882 105440 282887 105496
rect 279956 105438 282887 105440
rect 231209 105435 231275 105438
rect 256233 105435 256299 105438
rect 282821 105435 282887 105438
rect 231761 105226 231827 105229
rect 198089 105224 217058 105226
rect 198089 105168 198094 105224
rect 198150 105168 217058 105224
rect 198089 105166 217058 105168
rect 228988 105224 231827 105226
rect 228988 105168 231766 105224
rect 231822 105168 231827 105224
rect 228988 105166 231827 105168
rect 198089 105163 198155 105166
rect 231761 105163 231827 105166
rect 260189 105226 260255 105229
rect 260189 105224 268180 105226
rect 260189 105168 260194 105224
rect 260250 105168 268180 105224
rect 260189 105166 268180 105168
rect 260189 105163 260255 105166
rect 213913 104954 213979 104957
rect 213913 104952 217028 104954
rect 213913 104896 213918 104952
rect 213974 104896 217028 104952
rect 213913 104894 217028 104896
rect 213913 104891 213979 104894
rect 264421 104818 264487 104821
rect 238710 104816 264487 104818
rect 238710 104760 264426 104816
rect 264482 104760 264487 104816
rect 238710 104758 264487 104760
rect 238710 104682 238770 104758
rect 264421 104755 264487 104758
rect 267089 104818 267155 104821
rect 267089 104816 268180 104818
rect 267089 104760 267094 104816
rect 267150 104760 268180 104816
rect 267089 104758 268180 104760
rect 267089 104755 267155 104758
rect 281533 104682 281599 104685
rect 228988 104622 238770 104682
rect 279956 104680 281599 104682
rect 279956 104624 281538 104680
rect 281594 104624 281599 104680
rect 279956 104622 281599 104624
rect 281533 104619 281599 104622
rect 214005 104274 214071 104277
rect 231761 104274 231827 104277
rect 214005 104272 217028 104274
rect 214005 104216 214010 104272
rect 214066 104216 217028 104272
rect 214005 104214 217028 104216
rect 228988 104272 231827 104274
rect 228988 104216 231766 104272
rect 231822 104216 231827 104272
rect 228988 104214 231827 104216
rect 214005 104211 214071 104214
rect 231761 104211 231827 104214
rect 233969 104002 234035 104005
rect 268150 104002 268210 104380
rect 282821 104002 282887 104005
rect 233969 104000 268210 104002
rect 233969 103944 233974 104000
rect 234030 103944 268210 104000
rect 233969 103942 268210 103944
rect 279956 104000 282887 104002
rect 279956 103944 282826 104000
rect 282882 103944 282887 104000
rect 279956 103942 282887 103944
rect 233969 103939 234035 103942
rect 282821 103939 282887 103942
rect 264973 103866 265039 103869
rect 264973 103864 268180 103866
rect 264973 103808 264978 103864
rect 265034 103808 268180 103864
rect 264973 103806 268180 103808
rect 264973 103803 265039 103806
rect 231117 103730 231183 103733
rect 228988 103728 231183 103730
rect 228988 103672 231122 103728
rect 231178 103672 231183 103728
rect 228988 103670 231183 103672
rect 231117 103667 231183 103670
rect 213913 103594 213979 103597
rect 213913 103592 217028 103594
rect 213913 103536 213918 103592
rect 213974 103536 217028 103592
rect 213913 103534 217028 103536
rect 213913 103531 213979 103534
rect 264973 103458 265039 103461
rect 264973 103456 268180 103458
rect 264973 103400 264978 103456
rect 265034 103400 268180 103456
rect 264973 103398 268180 103400
rect 264973 103395 265039 103398
rect 233734 103322 233740 103324
rect 228988 103262 233740 103322
rect 233734 103260 233740 103262
rect 233804 103260 233810 103324
rect 282821 103186 282887 103189
rect 279956 103184 282887 103186
rect 279956 103128 282826 103184
rect 282882 103128 282887 103184
rect 279956 103126 282887 103128
rect 282821 103123 282887 103126
rect 265157 103050 265223 103053
rect 265157 103048 268180 103050
rect 265157 102992 265162 103048
rect 265218 102992 268180 103048
rect 265157 102990 268180 102992
rect 265157 102987 265223 102990
rect 166206 102444 166212 102508
rect 166276 102506 166282 102508
rect 216998 102506 217058 102884
rect 231761 102778 231827 102781
rect 228988 102776 231827 102778
rect 228988 102720 231766 102776
rect 231822 102720 231827 102776
rect 228988 102718 231827 102720
rect 231761 102715 231827 102718
rect 264421 102642 264487 102645
rect 264421 102640 268180 102642
rect 264421 102584 264426 102640
rect 264482 102584 268180 102640
rect 264421 102582 268180 102584
rect 264421 102579 264487 102582
rect 166276 102446 217058 102506
rect 166276 102444 166282 102446
rect 67357 102370 67423 102373
rect 68142 102370 68816 102376
rect 231393 102370 231459 102373
rect 67357 102368 68816 102370
rect 67357 102312 67362 102368
rect 67418 102316 68816 102368
rect 228988 102368 231459 102370
rect 67418 102312 68202 102316
rect 67357 102310 68202 102312
rect 228988 102312 231398 102368
rect 231454 102312 231459 102368
rect 228988 102310 231459 102312
rect 279956 102310 287070 102370
rect 67357 102307 67423 102310
rect 231393 102307 231459 102310
rect 213453 102234 213519 102237
rect 245101 102234 245167 102237
rect 287010 102234 287070 102310
rect 287278 102234 287284 102236
rect 213453 102232 217028 102234
rect 213453 102176 213458 102232
rect 213514 102176 217028 102232
rect 213453 102174 217028 102176
rect 245101 102232 268180 102234
rect 245101 102176 245106 102232
rect 245162 102176 268180 102232
rect 245101 102174 268180 102176
rect 287010 102174 287284 102234
rect 213453 102171 213519 102174
rect 245101 102171 245167 102174
rect 287278 102172 287284 102174
rect 287348 102172 287354 102236
rect 231761 102098 231827 102101
rect 244774 102098 244780 102100
rect 231761 102096 244780 102098
rect 231761 102040 231766 102096
rect 231822 102040 244780 102096
rect 231761 102038 244780 102040
rect 231761 102035 231827 102038
rect 244774 102036 244780 102038
rect 244844 102036 244850 102100
rect 230565 101826 230631 101829
rect 228988 101824 230631 101826
rect 228988 101768 230570 101824
rect 230626 101768 230631 101824
rect 228988 101766 230631 101768
rect 230565 101763 230631 101766
rect 264973 101826 265039 101829
rect 264973 101824 268180 101826
rect 264973 101768 264978 101824
rect 265034 101768 268180 101824
rect 264973 101766 268180 101768
rect 264973 101763 265039 101766
rect 281717 101690 281783 101693
rect 279956 101688 281783 101690
rect 279956 101632 281722 101688
rect 281778 101632 281783 101688
rect 279956 101630 281783 101632
rect 281717 101627 281783 101630
rect 214189 101554 214255 101557
rect 214189 101552 217028 101554
rect 214189 101496 214194 101552
rect 214250 101496 217028 101552
rect 214189 101494 217028 101496
rect 214189 101491 214255 101494
rect 231761 101418 231827 101421
rect 228988 101416 231827 101418
rect 228988 101360 231766 101416
rect 231822 101360 231827 101416
rect 228988 101358 231827 101360
rect 231761 101355 231827 101358
rect 258030 101222 268180 101282
rect 242157 101146 242223 101149
rect 258030 101146 258090 101222
rect 242157 101144 258090 101146
rect 242157 101088 242162 101144
rect 242218 101088 258090 101144
rect 242157 101086 258090 101088
rect 242157 101083 242223 101086
rect 213913 101010 213979 101013
rect 213913 101008 217028 101010
rect 213913 100952 213918 101008
rect 213974 100952 217028 101008
rect 213913 100950 217028 100952
rect 213913 100947 213979 100950
rect 231669 100874 231735 100877
rect 228988 100872 231735 100874
rect 228988 100816 231674 100872
rect 231730 100816 231735 100872
rect 228988 100814 231735 100816
rect 231669 100811 231735 100814
rect 267038 100812 267044 100876
rect 267108 100874 267114 100876
rect 281625 100874 281691 100877
rect 267108 100814 268180 100874
rect 279956 100872 281691 100874
rect 279956 100816 281630 100872
rect 281686 100816 281691 100872
rect 279956 100814 281691 100816
rect 267108 100812 267114 100814
rect 281625 100811 281691 100814
rect 67265 100738 67331 100741
rect 68142 100738 68816 100744
rect 67265 100736 68816 100738
rect 67265 100680 67270 100736
rect 67326 100684 68816 100736
rect 67326 100680 68202 100684
rect 67265 100678 68202 100680
rect 67265 100675 67331 100678
rect 230565 100466 230631 100469
rect 228988 100464 230631 100466
rect 228988 100408 230570 100464
rect 230626 100408 230631 100464
rect 228988 100406 230631 100408
rect 230565 100403 230631 100406
rect 264973 100466 265039 100469
rect 264973 100464 268180 100466
rect 264973 100408 264978 100464
rect 265034 100408 268180 100464
rect 264973 100406 268180 100408
rect 264973 100403 265039 100406
rect 214005 100330 214071 100333
rect 214005 100328 217028 100330
rect 214005 100272 214010 100328
rect 214066 100272 217028 100328
rect 214005 100270 217028 100272
rect 214005 100267 214071 100270
rect 281717 100194 281783 100197
rect 279956 100192 281783 100194
rect 279956 100136 281722 100192
rect 281778 100136 281783 100192
rect 279956 100134 281783 100136
rect 281717 100131 281783 100134
rect 236913 100058 236979 100061
rect 257521 100058 257587 100061
rect 236913 100056 257587 100058
rect 236913 100000 236918 100056
rect 236974 100000 257526 100056
rect 257582 100000 257587 100056
rect 236913 99998 257587 100000
rect 236913 99995 236979 99998
rect 257521 99995 257587 99998
rect 265065 100058 265131 100061
rect 265065 100056 268180 100058
rect 265065 100000 265070 100056
rect 265126 100000 268180 100056
rect 265065 99998 268180 100000
rect 265065 99995 265131 99998
rect 231301 99922 231367 99925
rect 228988 99920 231367 99922
rect 228988 99864 231306 99920
rect 231362 99864 231367 99920
rect 228988 99862 231367 99864
rect 231301 99859 231367 99862
rect 213913 99650 213979 99653
rect 262857 99650 262923 99653
rect 213913 99648 217028 99650
rect 213913 99592 213918 99648
rect 213974 99592 217028 99648
rect 213913 99590 217028 99592
rect 262857 99648 268180 99650
rect 262857 99592 262862 99648
rect 262918 99592 268180 99648
rect 262857 99590 268180 99592
rect 213913 99587 213979 99590
rect 262857 99587 262923 99590
rect 231117 99514 231183 99517
rect 228988 99512 231183 99514
rect 228988 99456 231122 99512
rect 231178 99456 231183 99512
rect 228988 99454 231183 99456
rect 231117 99451 231183 99454
rect 583017 99514 583083 99517
rect 583520 99514 584960 99604
rect 583017 99512 584960 99514
rect 583017 99456 583022 99512
rect 583078 99456 584960 99512
rect 583017 99454 584960 99456
rect 583017 99451 583083 99454
rect 282821 99378 282887 99381
rect 279956 99376 282887 99378
rect 279956 99320 282826 99376
rect 282882 99320 282887 99376
rect 583520 99364 584960 99454
rect 279956 99318 282887 99320
rect 282821 99315 282887 99318
rect 265065 99242 265131 99245
rect 265065 99240 268180 99242
rect 265065 99184 265070 99240
rect 265126 99184 268180 99240
rect 265065 99182 268180 99184
rect 265065 99179 265131 99182
rect 214097 98970 214163 98973
rect 230974 98970 230980 98972
rect 214097 98968 217028 98970
rect 214097 98912 214102 98968
rect 214158 98912 217028 98968
rect 214097 98910 217028 98912
rect 228988 98910 230980 98970
rect 214097 98907 214163 98910
rect 230974 98908 230980 98910
rect 231044 98908 231050 98972
rect 235349 98698 235415 98701
rect 262806 98698 262812 98700
rect 235349 98696 262812 98698
rect 235349 98640 235354 98696
rect 235410 98640 262812 98696
rect 235349 98638 262812 98640
rect 235349 98635 235415 98638
rect 262806 98636 262812 98638
rect 262876 98636 262882 98700
rect 264973 98698 265039 98701
rect 264973 98696 268180 98698
rect 264973 98640 264978 98696
rect 265034 98640 268180 98696
rect 264973 98638 268180 98640
rect 264973 98635 265039 98638
rect 231117 98562 231183 98565
rect 228988 98560 231183 98562
rect 228988 98504 231122 98560
rect 231178 98504 231183 98560
rect 228988 98502 231183 98504
rect 231117 98499 231183 98502
rect 213913 98290 213979 98293
rect 213913 98288 217028 98290
rect 213913 98232 213918 98288
rect 213974 98232 217028 98288
rect 213913 98230 217028 98232
rect 213913 98227 213979 98230
rect 232446 98018 232452 98020
rect 228988 97958 232452 98018
rect 232446 97956 232452 97958
rect 232516 97956 232522 98020
rect 267958 97956 267964 98020
rect 268028 98018 268034 98020
rect 268150 98018 268210 98260
rect 279374 98157 279434 98532
rect 279325 98152 279434 98157
rect 279325 98096 279330 98152
rect 279386 98096 279434 98152
rect 279325 98094 279434 98096
rect 279325 98091 279391 98094
rect 268028 97958 268210 98018
rect 268028 97956 268034 97958
rect 204897 97882 204963 97885
rect 214465 97882 214531 97885
rect 204897 97880 214531 97882
rect 204897 97824 204902 97880
rect 204958 97824 214470 97880
rect 214526 97824 214531 97880
rect 204897 97822 214531 97824
rect 204897 97819 204963 97822
rect 214465 97819 214531 97822
rect 264973 97882 265039 97885
rect 282821 97882 282887 97885
rect 264973 97880 268180 97882
rect 264973 97824 264978 97880
rect 265034 97824 268180 97880
rect 264973 97822 268180 97824
rect 279956 97880 282887 97882
rect 279956 97824 282826 97880
rect 282882 97824 282887 97880
rect 279956 97822 282887 97824
rect 264973 97819 265039 97822
rect 282821 97819 282887 97822
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 213913 97610 213979 97613
rect 231761 97610 231827 97613
rect 213913 97608 217028 97610
rect 213913 97552 213918 97608
rect 213974 97552 217028 97608
rect 213913 97550 217028 97552
rect 228988 97608 231827 97610
rect 228988 97552 231766 97608
rect 231822 97552 231827 97608
rect 228988 97550 231827 97552
rect 213913 97547 213979 97550
rect 231761 97547 231827 97550
rect 265065 97474 265131 97477
rect 265065 97472 268180 97474
rect 265065 97416 265070 97472
rect 265126 97416 268180 97472
rect 265065 97414 268180 97416
rect 265065 97411 265131 97414
rect 229134 97140 229140 97204
rect 229204 97202 229210 97204
rect 229204 97142 258090 97202
rect 229204 97140 229210 97142
rect 230473 97066 230539 97069
rect 228988 97064 230539 97066
rect 228988 97008 230478 97064
rect 230534 97008 230539 97064
rect 228988 97006 230539 97008
rect 230473 97003 230539 97006
rect 214741 96930 214807 96933
rect 214741 96928 217028 96930
rect 214741 96872 214746 96928
rect 214802 96872 217028 96928
rect 214741 96870 217028 96872
rect 214741 96867 214807 96870
rect 258030 96794 258090 97142
rect 265893 97066 265959 97069
rect 282177 97066 282243 97069
rect 265893 97064 268180 97066
rect 265893 97008 265898 97064
rect 265954 97008 268180 97064
rect 265893 97006 268180 97008
rect 279956 97064 282243 97066
rect 279956 97008 282182 97064
rect 282238 97008 282243 97064
rect 279956 97006 282243 97008
rect 265893 97003 265959 97006
rect 282177 97003 282243 97006
rect 258030 96734 268210 96794
rect 229134 96658 229140 96660
rect 228988 96598 229140 96658
rect 229134 96596 229140 96598
rect 229204 96658 229210 96660
rect 231669 96658 231735 96661
rect 229204 96656 231735 96658
rect 229204 96600 231674 96656
rect 231730 96600 231735 96656
rect 268150 96628 268210 96734
rect 229204 96598 231735 96600
rect 229204 96596 229210 96598
rect 231669 96595 231735 96598
rect 214005 96386 214071 96389
rect 214005 96384 217028 96386
rect 214005 96328 214010 96384
rect 214066 96328 217028 96384
rect 214005 96326 217028 96328
rect 214005 96323 214071 96326
rect 230565 96250 230631 96253
rect 228988 96248 230631 96250
rect 228988 96192 230570 96248
rect 230626 96192 230631 96248
rect 228988 96190 230631 96192
rect 230565 96187 230631 96190
rect 219249 95980 219315 95981
rect 219198 95978 219204 95980
rect 219158 95918 219204 95978
rect 219268 95976 219315 95980
rect 219310 95920 219315 95976
rect 219198 95916 219204 95918
rect 219268 95916 219315 95920
rect 219249 95915 219315 95916
rect 226977 95978 227043 95981
rect 262857 95978 262923 95981
rect 226977 95976 262923 95978
rect 226977 95920 226982 95976
rect 227038 95920 262862 95976
rect 262918 95920 262923 95976
rect 226977 95918 262923 95920
rect 226977 95915 227043 95918
rect 262857 95915 262923 95918
rect 166390 95780 166396 95844
rect 166460 95842 166466 95844
rect 214189 95842 214255 95845
rect 219157 95844 219223 95845
rect 219157 95842 219204 95844
rect 166460 95840 214255 95842
rect 166460 95784 214194 95840
rect 214250 95784 214255 95840
rect 166460 95782 214255 95784
rect 219112 95840 219204 95842
rect 219112 95784 219162 95840
rect 219112 95782 219204 95784
rect 166460 95780 166466 95782
rect 214189 95779 214255 95782
rect 219157 95780 219204 95782
rect 219268 95780 219274 95844
rect 219157 95779 219223 95780
rect 224902 95508 224908 95572
rect 224972 95570 224978 95572
rect 228582 95570 228588 95572
rect 224972 95510 228588 95570
rect 224972 95508 224978 95510
rect 228582 95508 228588 95510
rect 228652 95508 228658 95572
rect 227713 95298 227779 95301
rect 268150 95298 268210 96220
rect 278773 95842 278839 95845
rect 279374 95842 279434 96356
rect 278773 95840 279434 95842
rect 278773 95784 278778 95840
rect 278834 95784 279434 95840
rect 278773 95782 279434 95784
rect 278773 95779 278839 95782
rect 227713 95296 268210 95298
rect 227713 95240 227718 95296
rect 227774 95240 268210 95296
rect 227713 95238 268210 95240
rect 227713 95235 227779 95238
rect 205398 95100 205404 95164
rect 205468 95162 205474 95164
rect 279325 95162 279391 95165
rect 205468 95160 279391 95162
rect 205468 95104 279330 95160
rect 279386 95104 279391 95160
rect 205468 95102 279391 95104
rect 205468 95100 205474 95102
rect 279325 95099 279391 95102
rect 100661 94756 100727 94757
rect 100624 94692 100630 94756
rect 100694 94754 100727 94756
rect 100694 94752 100786 94754
rect 100722 94696 100786 94752
rect 100694 94694 100786 94696
rect 100694 94692 100727 94694
rect 151302 94692 151308 94756
rect 151372 94754 151378 94756
rect 151760 94754 151766 94756
rect 151372 94694 151766 94754
rect 151372 94692 151378 94694
rect 151760 94692 151766 94694
rect 151830 94692 151836 94756
rect 100661 94691 100727 94692
rect 133873 94482 133939 94485
rect 173249 94482 173315 94485
rect 133873 94480 173315 94482
rect 133873 94424 133878 94480
rect 133934 94424 173254 94480
rect 173310 94424 173315 94480
rect 133873 94422 173315 94424
rect 133873 94419 133939 94422
rect 173249 94419 173315 94422
rect 216213 94482 216279 94485
rect 245193 94482 245259 94485
rect 216213 94480 245259 94482
rect 216213 94424 216218 94480
rect 216274 94424 245198 94480
rect 245254 94424 245259 94480
rect 216213 94422 245259 94424
rect 216213 94419 216279 94422
rect 245193 94419 245259 94422
rect 126646 94012 126652 94076
rect 126716 94074 126722 94076
rect 180333 94074 180399 94077
rect 126716 94072 180399 94074
rect 126716 94016 180338 94072
rect 180394 94016 180399 94072
rect 126716 94014 180399 94016
rect 126716 94012 126722 94014
rect 180333 94011 180399 94014
rect 111926 93876 111932 93940
rect 111996 93938 112002 93940
rect 187049 93938 187115 93941
rect 111996 93936 187115 93938
rect 111996 93880 187054 93936
rect 187110 93880 187115 93936
rect 111996 93878 187115 93880
rect 111996 93876 112002 93878
rect 187049 93875 187115 93878
rect 114870 93740 114876 93804
rect 114940 93802 114946 93804
rect 211797 93802 211863 93805
rect 114940 93800 211863 93802
rect 114940 93744 211802 93800
rect 211858 93744 211863 93800
rect 114940 93742 211863 93744
rect 114940 93740 114946 93742
rect 211797 93739 211863 93742
rect 134374 93604 134380 93668
rect 134444 93666 134450 93668
rect 135805 93666 135871 93669
rect 134444 93664 135871 93666
rect 134444 93608 135810 93664
rect 135866 93608 135871 93664
rect 134444 93606 135871 93608
rect 134444 93604 134450 93606
rect 135805 93603 135871 93606
rect 135989 93666 136055 93669
rect 216121 93666 216187 93669
rect 135989 93664 216187 93666
rect 135989 93608 135994 93664
rect 136050 93608 216126 93664
rect 216182 93608 216187 93664
rect 135989 93606 216187 93608
rect 135989 93603 136055 93606
rect 216121 93603 216187 93606
rect 117129 93532 117195 93533
rect 121729 93532 121795 93533
rect 117078 93530 117084 93532
rect 117038 93470 117084 93530
rect 117148 93528 117195 93532
rect 121678 93530 121684 93532
rect 117190 93472 117195 93528
rect 117078 93468 117084 93470
rect 117148 93468 117195 93472
rect 121638 93470 121684 93530
rect 121748 93528 121795 93532
rect 121790 93472 121795 93528
rect 121678 93468 121684 93470
rect 121748 93468 121795 93472
rect 123150 93468 123156 93532
rect 123220 93530 123226 93532
rect 167913 93530 167979 93533
rect 123220 93528 167979 93530
rect 123220 93472 167918 93528
rect 167974 93472 167979 93528
rect 123220 93470 167979 93472
rect 123220 93468 123226 93470
rect 117129 93467 117195 93468
rect 121729 93467 121795 93468
rect 167913 93467 167979 93470
rect 133086 93332 133092 93396
rect 133156 93394 133162 93396
rect 135989 93394 136055 93397
rect 133156 93392 136055 93394
rect 133156 93336 135994 93392
rect 136050 93336 136055 93392
rect 133156 93334 136055 93336
rect 133156 93332 133162 93334
rect 135989 93331 136055 93334
rect 110137 93260 110203 93261
rect 113817 93260 113883 93261
rect 110086 93258 110092 93260
rect 110046 93198 110092 93258
rect 110156 93256 110203 93260
rect 113766 93258 113772 93260
rect 110198 93200 110203 93256
rect 110086 93196 110092 93198
rect 110156 93196 110203 93200
rect 113726 93198 113772 93258
rect 113836 93256 113883 93260
rect 113878 93200 113883 93256
rect 113766 93196 113772 93198
rect 113836 93196 113883 93200
rect 110137 93195 110203 93196
rect 113817 93195 113883 93196
rect 215937 93258 216003 93261
rect 241053 93258 241119 93261
rect 215937 93256 241119 93258
rect 215937 93200 215942 93256
rect 215998 93200 241058 93256
rect 241114 93200 241119 93256
rect 215937 93198 241119 93200
rect 215937 93195 216003 93198
rect 241053 93195 241119 93198
rect 207749 93122 207815 93125
rect 270493 93122 270559 93125
rect 207749 93120 270559 93122
rect 207749 93064 207754 93120
rect 207810 93064 270498 93120
rect 270554 93064 270559 93120
rect 207749 93062 270559 93064
rect 207749 93059 207815 93062
rect 270493 93059 270559 93062
rect 253197 92578 253263 92581
rect 254853 92578 254919 92581
rect 253197 92576 254919 92578
rect 253197 92520 253202 92576
rect 253258 92520 254858 92576
rect 254914 92520 254919 92576
rect 253197 92518 254919 92520
rect 253197 92515 253263 92518
rect 254853 92515 254919 92518
rect 84377 92444 84443 92445
rect 84326 92442 84332 92444
rect 84286 92382 84332 92442
rect 84396 92440 84443 92444
rect 84438 92384 84443 92440
rect 84326 92380 84332 92382
rect 84396 92380 84443 92384
rect 88926 92380 88932 92444
rect 88996 92442 89002 92444
rect 89069 92442 89135 92445
rect 99097 92444 99163 92445
rect 106825 92444 106891 92445
rect 99046 92442 99052 92444
rect 88996 92440 89135 92442
rect 88996 92384 89074 92440
rect 89130 92384 89135 92440
rect 88996 92382 89135 92384
rect 99006 92382 99052 92442
rect 99116 92440 99163 92444
rect 106774 92442 106780 92444
rect 99158 92384 99163 92440
rect 88996 92380 89002 92382
rect 84377 92379 84443 92380
rect 89069 92379 89135 92382
rect 99046 92380 99052 92382
rect 99116 92380 99163 92384
rect 106734 92382 106780 92442
rect 106844 92440 106891 92444
rect 106886 92384 106891 92440
rect 106774 92380 106780 92382
rect 106844 92380 106891 92384
rect 109166 92380 109172 92444
rect 109236 92442 109242 92444
rect 109677 92442 109743 92445
rect 110689 92444 110755 92445
rect 110638 92442 110644 92444
rect 109236 92440 109743 92442
rect 109236 92384 109682 92440
rect 109738 92384 109743 92440
rect 109236 92382 109743 92384
rect 110598 92382 110644 92442
rect 110708 92440 110755 92444
rect 110750 92384 110755 92440
rect 109236 92380 109242 92382
rect 99097 92379 99163 92380
rect 106825 92379 106891 92380
rect 109677 92379 109743 92382
rect 110638 92380 110644 92382
rect 110708 92380 110755 92384
rect 111190 92380 111196 92444
rect 111260 92442 111266 92444
rect 111517 92442 111583 92445
rect 124121 92444 124187 92445
rect 136081 92444 136147 92445
rect 124070 92442 124076 92444
rect 111260 92440 111583 92442
rect 111260 92384 111522 92440
rect 111578 92384 111583 92440
rect 111260 92382 111583 92384
rect 124030 92382 124076 92442
rect 124140 92440 124187 92444
rect 136030 92442 136036 92444
rect 124182 92384 124187 92440
rect 111260 92380 111266 92382
rect 110689 92379 110755 92380
rect 111517 92379 111583 92382
rect 124070 92380 124076 92382
rect 124140 92380 124187 92384
rect 135990 92382 136036 92442
rect 136100 92440 136147 92444
rect 136142 92384 136147 92440
rect 136030 92380 136036 92382
rect 136100 92380 136147 92384
rect 151302 92380 151308 92444
rect 151372 92442 151378 92444
rect 151445 92442 151511 92445
rect 151372 92440 151511 92442
rect 151372 92384 151450 92440
rect 151506 92384 151511 92440
rect 151372 92382 151511 92384
rect 151372 92380 151378 92382
rect 124121 92379 124187 92380
rect 136081 92379 136147 92380
rect 151445 92379 151511 92382
rect 116710 92244 116716 92308
rect 116780 92306 116786 92308
rect 216029 92306 216095 92309
rect 116780 92304 216095 92306
rect 116780 92248 216034 92304
rect 216090 92248 216095 92304
rect 116780 92246 216095 92248
rect 116780 92244 116786 92246
rect 216029 92243 216095 92246
rect 130694 92108 130700 92172
rect 130764 92170 130770 92172
rect 169017 92170 169083 92173
rect 130764 92168 169083 92170
rect 130764 92112 169022 92168
rect 169078 92112 169083 92168
rect 130764 92110 169083 92112
rect 130764 92108 130770 92110
rect 169017 92107 169083 92110
rect 96337 91900 96403 91901
rect 96286 91898 96292 91900
rect 96246 91838 96292 91898
rect 96356 91896 96403 91900
rect 96398 91840 96403 91896
rect 96286 91836 96292 91838
rect 96356 91836 96403 91840
rect 96337 91835 96403 91836
rect 224217 91898 224283 91901
rect 242198 91898 242204 91900
rect 224217 91896 242204 91898
rect 224217 91840 224222 91896
rect 224278 91840 242204 91896
rect 224217 91838 242204 91840
rect 224217 91835 224283 91838
rect 242198 91836 242204 91838
rect 242268 91836 242274 91900
rect 92606 91700 92612 91764
rect 92676 91762 92682 91764
rect 93209 91762 93275 91765
rect 92676 91760 93275 91762
rect 92676 91704 93214 91760
rect 93270 91704 93275 91760
rect 92676 91702 93275 91704
rect 92676 91700 92682 91702
rect 93209 91699 93275 91702
rect 98126 91700 98132 91764
rect 98196 91762 98202 91764
rect 99281 91762 99347 91765
rect 98196 91760 99347 91762
rect 98196 91704 99286 91760
rect 99342 91704 99347 91760
rect 98196 91702 99347 91704
rect 98196 91700 98202 91702
rect 99281 91699 99347 91702
rect 119654 91700 119660 91764
rect 119724 91762 119730 91764
rect 119797 91762 119863 91765
rect 119724 91760 119863 91762
rect 119724 91704 119802 91760
rect 119858 91704 119863 91760
rect 119724 91702 119863 91704
rect 119724 91700 119730 91702
rect 119797 91699 119863 91702
rect 209129 91762 209195 91765
rect 229686 91762 229692 91764
rect 209129 91760 229692 91762
rect 209129 91704 209134 91760
rect 209190 91704 229692 91760
rect 209129 91702 229692 91704
rect 209129 91699 209195 91702
rect 229686 91700 229692 91702
rect 229756 91700 229762 91764
rect 104566 91564 104572 91628
rect 104636 91626 104642 91628
rect 209313 91626 209379 91629
rect 104636 91624 209379 91626
rect 104636 91568 209318 91624
rect 209374 91568 209379 91624
rect 104636 91566 209379 91568
rect 104636 91564 104642 91566
rect 209313 91563 209379 91566
rect 122782 91428 122788 91492
rect 122852 91490 122858 91492
rect 124029 91490 124095 91493
rect 122852 91488 124095 91490
rect 122852 91432 124034 91488
rect 124090 91432 124095 91488
rect 122852 91430 124095 91432
rect 122852 91428 122858 91430
rect 124029 91427 124095 91430
rect 96654 91292 96660 91356
rect 96724 91354 96730 91356
rect 97901 91354 97967 91357
rect 96724 91352 97967 91354
rect 96724 91296 97906 91352
rect 97962 91296 97967 91352
rect 96724 91294 97967 91296
rect 96724 91292 96730 91294
rect 97901 91291 97967 91294
rect 101806 91292 101812 91356
rect 101876 91354 101882 91356
rect 102041 91354 102107 91357
rect 101876 91352 102107 91354
rect 101876 91296 102046 91352
rect 102102 91296 102107 91352
rect 101876 91294 102107 91296
rect 101876 91292 101882 91294
rect 102041 91291 102107 91294
rect 113214 91292 113220 91356
rect 113284 91354 113290 91356
rect 114277 91354 114343 91357
rect 113284 91352 114343 91354
rect 113284 91296 114282 91352
rect 114338 91296 114343 91352
rect 113284 91294 114343 91296
rect 113284 91292 113290 91294
rect 114277 91291 114343 91294
rect 115749 91356 115815 91357
rect 115749 91352 115796 91356
rect 115860 91354 115866 91356
rect 115749 91296 115754 91352
rect 115749 91292 115796 91296
rect 115860 91294 115906 91354
rect 115860 91292 115866 91294
rect 117998 91292 118004 91356
rect 118068 91354 118074 91356
rect 118601 91354 118667 91357
rect 118068 91352 118667 91354
rect 118068 91296 118606 91352
rect 118662 91296 118667 91352
rect 118068 91294 118667 91296
rect 118068 91292 118074 91294
rect 115749 91291 115815 91292
rect 118601 91291 118667 91294
rect 124438 91292 124444 91356
rect 124508 91354 124514 91356
rect 125409 91354 125475 91357
rect 124508 91352 125475 91354
rect 124508 91296 125414 91352
rect 125470 91296 125475 91352
rect 124508 91294 125475 91296
rect 124508 91292 124514 91294
rect 125409 91291 125475 91294
rect 125726 91292 125732 91356
rect 125796 91354 125802 91356
rect 126881 91354 126947 91357
rect 125796 91352 126947 91354
rect 125796 91296 126886 91352
rect 126942 91296 126947 91352
rect 125796 91294 126947 91296
rect 125796 91292 125802 91294
rect 126881 91291 126947 91294
rect 151537 91354 151603 91357
rect 151670 91354 151676 91356
rect 151537 91352 151676 91354
rect 151537 91296 151542 91352
rect 151598 91296 151676 91352
rect 151537 91294 151676 91296
rect 151537 91291 151603 91294
rect 151670 91292 151676 91294
rect 151740 91292 151746 91356
rect 74758 91156 74764 91220
rect 74828 91218 74834 91220
rect 75361 91218 75427 91221
rect 74828 91216 75427 91218
rect 74828 91160 75366 91216
rect 75422 91160 75427 91216
rect 74828 91158 75427 91160
rect 74828 91156 74834 91158
rect 75361 91155 75427 91158
rect 85798 91156 85804 91220
rect 85868 91218 85874 91220
rect 86217 91218 86283 91221
rect 85868 91216 86283 91218
rect 85868 91160 86222 91216
rect 86278 91160 86283 91216
rect 85868 91158 86283 91160
rect 85868 91156 85874 91158
rect 86217 91155 86283 91158
rect 86718 91156 86724 91220
rect 86788 91218 86794 91220
rect 86861 91218 86927 91221
rect 86788 91216 86927 91218
rect 86788 91160 86866 91216
rect 86922 91160 86927 91216
rect 86788 91158 86927 91160
rect 86788 91156 86794 91158
rect 86861 91155 86927 91158
rect 88006 91156 88012 91220
rect 88076 91218 88082 91220
rect 88241 91218 88307 91221
rect 88076 91216 88307 91218
rect 88076 91160 88246 91216
rect 88302 91160 88307 91216
rect 88076 91158 88307 91160
rect 88076 91156 88082 91158
rect 88241 91155 88307 91158
rect 90214 91156 90220 91220
rect 90284 91218 90290 91220
rect 91001 91218 91067 91221
rect 90284 91216 91067 91218
rect 90284 91160 91006 91216
rect 91062 91160 91067 91216
rect 90284 91158 91067 91160
rect 90284 91156 90290 91158
rect 91001 91155 91067 91158
rect 91318 91156 91324 91220
rect 91388 91218 91394 91220
rect 91921 91218 91987 91221
rect 91388 91216 91987 91218
rect 91388 91160 91926 91216
rect 91982 91160 91987 91216
rect 91388 91158 91987 91160
rect 91388 91156 91394 91158
rect 91921 91155 91987 91158
rect 93894 91156 93900 91220
rect 93964 91218 93970 91220
rect 95141 91218 95207 91221
rect 93964 91216 95207 91218
rect 93964 91160 95146 91216
rect 95202 91160 95207 91216
rect 93964 91158 95207 91160
rect 93964 91156 93970 91158
rect 95141 91155 95207 91158
rect 97206 91156 97212 91220
rect 97276 91218 97282 91220
rect 97809 91218 97875 91221
rect 97276 91216 97875 91218
rect 97276 91160 97814 91216
rect 97870 91160 97875 91216
rect 97276 91158 97875 91160
rect 97276 91156 97282 91158
rect 97809 91155 97875 91158
rect 98494 91156 98500 91220
rect 98564 91218 98570 91220
rect 99189 91218 99255 91221
rect 100017 91220 100083 91221
rect 99966 91218 99972 91220
rect 98564 91216 99255 91218
rect 98564 91160 99194 91216
rect 99250 91160 99255 91216
rect 98564 91158 99255 91160
rect 99926 91158 99972 91218
rect 100036 91216 100083 91220
rect 100078 91160 100083 91216
rect 98564 91156 98570 91158
rect 99189 91155 99255 91158
rect 99966 91156 99972 91158
rect 100036 91156 100083 91160
rect 100886 91156 100892 91220
rect 100956 91218 100962 91220
rect 101213 91218 101279 91221
rect 101949 91220 102015 91221
rect 101949 91218 101996 91220
rect 100956 91216 101279 91218
rect 100956 91160 101218 91216
rect 101274 91160 101279 91216
rect 100956 91158 101279 91160
rect 101904 91216 101996 91218
rect 101904 91160 101954 91216
rect 101904 91158 101996 91160
rect 100956 91156 100962 91158
rect 100017 91155 100083 91156
rect 101213 91155 101279 91158
rect 101949 91156 101996 91158
rect 102060 91156 102066 91220
rect 102542 91156 102548 91220
rect 102612 91156 102618 91220
rect 102726 91156 102732 91220
rect 102796 91218 102802 91220
rect 103421 91218 103487 91221
rect 102796 91216 103487 91218
rect 102796 91160 103426 91216
rect 103482 91160 103487 91216
rect 102796 91158 103487 91160
rect 102796 91156 102802 91158
rect 101949 91155 102015 91156
rect 102550 91082 102610 91156
rect 103421 91155 103487 91158
rect 104198 91156 104204 91220
rect 104268 91218 104274 91220
rect 104433 91218 104499 91221
rect 105537 91220 105603 91221
rect 105486 91218 105492 91220
rect 104268 91216 104499 91218
rect 104268 91160 104438 91216
rect 104494 91160 104499 91216
rect 104268 91158 104499 91160
rect 105446 91158 105492 91218
rect 105556 91216 105603 91220
rect 105598 91160 105603 91216
rect 104268 91156 104274 91158
rect 104433 91155 104499 91158
rect 105486 91156 105492 91158
rect 105556 91156 105603 91160
rect 105670 91156 105676 91220
rect 105740 91218 105746 91220
rect 106089 91218 106155 91221
rect 105740 91216 106155 91218
rect 105740 91160 106094 91216
rect 106150 91160 106155 91216
rect 105740 91158 106155 91160
rect 105740 91156 105746 91158
rect 105537 91155 105603 91156
rect 106089 91155 106155 91158
rect 106406 91156 106412 91220
rect 106476 91218 106482 91220
rect 107561 91218 107627 91221
rect 106476 91216 107627 91218
rect 106476 91160 107566 91216
rect 107622 91160 107627 91216
rect 106476 91158 107627 91160
rect 106476 91156 106482 91158
rect 107561 91155 107627 91158
rect 108062 91156 108068 91220
rect 108132 91218 108138 91220
rect 108481 91218 108547 91221
rect 108132 91216 108547 91218
rect 108132 91160 108486 91216
rect 108542 91160 108547 91216
rect 108132 91158 108547 91160
rect 108132 91156 108138 91158
rect 108481 91155 108547 91158
rect 109534 91156 109540 91220
rect 109604 91218 109610 91220
rect 110229 91218 110295 91221
rect 109604 91216 110295 91218
rect 109604 91160 110234 91216
rect 110290 91160 110295 91216
rect 109604 91158 110295 91160
rect 109604 91156 109610 91158
rect 110229 91155 110295 91158
rect 112294 91156 112300 91220
rect 112364 91218 112370 91220
rect 112713 91218 112779 91221
rect 114369 91220 114435 91221
rect 114318 91218 114324 91220
rect 112364 91216 112779 91218
rect 112364 91160 112718 91216
rect 112774 91160 112779 91216
rect 112364 91158 112779 91160
rect 114278 91158 114324 91218
rect 114388 91216 114435 91220
rect 114430 91160 114435 91216
rect 112364 91156 112370 91158
rect 112713 91155 112779 91158
rect 114318 91156 114324 91158
rect 114388 91156 114435 91160
rect 115422 91156 115428 91220
rect 115492 91218 115498 91220
rect 115841 91218 115907 91221
rect 115492 91216 115907 91218
rect 115492 91160 115846 91216
rect 115902 91160 115907 91216
rect 115492 91158 115907 91160
rect 115492 91156 115498 91158
rect 114369 91155 114435 91156
rect 115841 91155 115907 91158
rect 118182 91156 118188 91220
rect 118252 91218 118258 91220
rect 118509 91218 118575 91221
rect 118252 91216 118575 91218
rect 118252 91160 118514 91216
rect 118570 91160 118575 91216
rect 118252 91158 118575 91160
rect 118252 91156 118258 91158
rect 118509 91155 118575 91158
rect 119286 91156 119292 91220
rect 119356 91218 119362 91220
rect 119889 91218 119955 91221
rect 119356 91216 119955 91218
rect 119356 91160 119894 91216
rect 119950 91160 119955 91216
rect 119356 91158 119955 91160
rect 119356 91156 119362 91158
rect 119889 91155 119955 91158
rect 120206 91156 120212 91220
rect 120276 91218 120282 91220
rect 120441 91218 120507 91221
rect 120276 91216 120507 91218
rect 120276 91160 120446 91216
rect 120502 91160 120507 91216
rect 120276 91158 120507 91160
rect 120276 91156 120282 91158
rect 120441 91155 120507 91158
rect 120574 91156 120580 91220
rect 120644 91218 120650 91220
rect 120717 91218 120783 91221
rect 120644 91216 120783 91218
rect 120644 91160 120722 91216
rect 120778 91160 120783 91216
rect 120644 91158 120783 91160
rect 120644 91156 120650 91158
rect 120717 91155 120783 91158
rect 122046 91156 122052 91220
rect 122116 91218 122122 91220
rect 122741 91218 122807 91221
rect 122116 91216 122807 91218
rect 122116 91160 122746 91216
rect 122802 91160 122807 91216
rect 122116 91158 122807 91160
rect 122116 91156 122122 91158
rect 122741 91155 122807 91158
rect 125358 91156 125364 91220
rect 125428 91218 125434 91220
rect 125501 91218 125567 91221
rect 125428 91216 125567 91218
rect 125428 91160 125506 91216
rect 125562 91160 125567 91216
rect 125428 91158 125567 91160
rect 125428 91156 125434 91158
rect 125501 91155 125567 91158
rect 126462 91156 126468 91220
rect 126532 91218 126538 91220
rect 126789 91218 126855 91221
rect 126532 91216 126855 91218
rect 126532 91160 126794 91216
rect 126850 91160 126855 91216
rect 126532 91158 126855 91160
rect 126532 91156 126538 91158
rect 126789 91155 126855 91158
rect 127566 91156 127572 91220
rect 127636 91218 127642 91220
rect 128261 91218 128327 91221
rect 127636 91216 128327 91218
rect 127636 91160 128266 91216
rect 128322 91160 128327 91216
rect 127636 91158 128327 91160
rect 127636 91156 127642 91158
rect 128261 91155 128327 91158
rect 129406 91156 129412 91220
rect 129476 91218 129482 91220
rect 129641 91218 129707 91221
rect 132401 91220 132467 91221
rect 132350 91218 132356 91220
rect 129476 91216 129707 91218
rect 129476 91160 129646 91216
rect 129702 91160 129707 91216
rect 129476 91158 129707 91160
rect 132310 91158 132356 91218
rect 132420 91216 132467 91220
rect 132462 91160 132467 91216
rect 129476 91156 129482 91158
rect 129641 91155 129707 91158
rect 132350 91156 132356 91158
rect 132420 91156 132467 91160
rect 151486 91156 151492 91220
rect 151556 91218 151562 91220
rect 151629 91218 151695 91221
rect 151556 91216 151695 91218
rect 151556 91160 151634 91216
rect 151690 91160 151695 91216
rect 151556 91158 151695 91160
rect 151556 91156 151562 91158
rect 132401 91155 132467 91156
rect 151629 91155 151695 91158
rect 152038 91156 152044 91220
rect 152108 91218 152114 91220
rect 152457 91218 152523 91221
rect 152108 91216 152523 91218
rect 152108 91160 152462 91216
rect 152518 91160 152523 91216
rect 152108 91158 152523 91160
rect 152108 91156 152114 91158
rect 152457 91155 152523 91158
rect 211981 91082 212047 91085
rect 102550 91080 212047 91082
rect 102550 91024 211986 91080
rect 212042 91024 212047 91080
rect 102550 91022 212047 91024
rect 211981 91019 212047 91022
rect 107694 90884 107700 90948
rect 107764 90946 107770 90948
rect 199469 90946 199535 90949
rect 107764 90944 199535 90946
rect 107764 90888 199474 90944
rect 199530 90888 199535 90944
rect 107764 90886 199535 90888
rect 107764 90884 107770 90886
rect 199469 90883 199535 90886
rect 94998 90748 95004 90812
rect 95068 90810 95074 90812
rect 165061 90810 165127 90813
rect 95068 90808 165127 90810
rect 95068 90752 165066 90808
rect 165122 90752 165127 90808
rect 95068 90750 165127 90752
rect 95068 90748 95074 90750
rect 165061 90747 165127 90750
rect 197118 90340 197124 90404
rect 197188 90402 197194 90404
rect 580165 90402 580231 90405
rect 197188 90400 580231 90402
rect 197188 90344 580170 90400
rect 580226 90344 580231 90400
rect 197188 90342 580231 90344
rect 197188 90340 197194 90342
rect 580165 90339 580231 90342
rect 93209 89722 93275 89725
rect 209221 89722 209287 89725
rect 93209 89720 209287 89722
rect 93209 89664 93214 89720
rect 93270 89664 209226 89720
rect 209282 89664 209287 89720
rect 93209 89662 209287 89664
rect 93209 89659 93275 89662
rect 209221 89659 209287 89662
rect 99281 89586 99347 89589
rect 174813 89586 174879 89589
rect 99281 89584 174879 89586
rect 99281 89528 99286 89584
rect 99342 89528 174818 89584
rect 174874 89528 174879 89584
rect 99281 89526 174879 89528
rect 99281 89523 99347 89526
rect 174813 89523 174879 89526
rect 113817 89450 113883 89453
rect 176101 89450 176167 89453
rect 113817 89448 176167 89450
rect 113817 89392 113822 89448
rect 113878 89392 176106 89448
rect 176162 89392 176167 89448
rect 113817 89390 176167 89392
rect 113817 89387 113883 89390
rect 176101 89387 176167 89390
rect 191189 89042 191255 89045
rect 280153 89042 280219 89045
rect 191189 89040 280219 89042
rect 191189 88984 191194 89040
rect 191250 88984 280158 89040
rect 280214 88984 280219 89040
rect 191189 88982 280219 88984
rect 191189 88979 191255 88982
rect 280153 88979 280219 88982
rect 75361 88226 75427 88229
rect 214005 88226 214071 88229
rect 75361 88224 214071 88226
rect 75361 88168 75366 88224
rect 75422 88168 214010 88224
rect 214066 88168 214071 88224
rect 75361 88166 214071 88168
rect 75361 88163 75427 88166
rect 214005 88163 214071 88166
rect 91921 88090 91987 88093
rect 181621 88090 181687 88093
rect 91921 88088 181687 88090
rect 91921 88032 91926 88088
rect 91982 88032 181626 88088
rect 181682 88032 181687 88088
rect 91921 88030 181687 88032
rect 91921 88027 91987 88030
rect 181621 88027 181687 88030
rect 108481 87954 108547 87957
rect 173157 87954 173223 87957
rect 108481 87952 173223 87954
rect 108481 87896 108486 87952
rect 108542 87896 173162 87952
rect 173218 87896 173223 87952
rect 108481 87894 173223 87896
rect 108481 87891 108547 87894
rect 173157 87891 173223 87894
rect 213269 87546 213335 87549
rect 246481 87546 246547 87549
rect 213269 87544 246547 87546
rect 213269 87488 213274 87544
rect 213330 87488 246486 87544
rect 246542 87488 246547 87544
rect 213269 87486 246547 87488
rect 213269 87483 213335 87486
rect 246481 87483 246547 87486
rect 101213 86866 101279 86869
rect 196801 86866 196867 86869
rect 101213 86864 196867 86866
rect 101213 86808 101218 86864
rect 101274 86808 196806 86864
rect 196862 86808 196867 86864
rect 101213 86806 196867 86808
rect 101213 86803 101279 86806
rect 196801 86803 196867 86806
rect 219198 86804 219204 86868
rect 219268 86866 219274 86868
rect 279049 86866 279115 86869
rect 219268 86864 279115 86866
rect 219268 86808 279054 86864
rect 279110 86808 279115 86864
rect 219268 86806 279115 86808
rect 219268 86804 219274 86806
rect 279049 86803 279115 86806
rect 100017 86730 100083 86733
rect 167637 86730 167703 86733
rect 100017 86728 167703 86730
rect 100017 86672 100022 86728
rect 100078 86672 167642 86728
rect 167698 86672 167703 86728
rect 100017 86670 167703 86672
rect 100017 86667 100083 86670
rect 167637 86667 167703 86670
rect 220169 86186 220235 86189
rect 267038 86186 267044 86188
rect 220169 86184 267044 86186
rect 220169 86128 220174 86184
rect 220230 86128 267044 86184
rect 220169 86126 267044 86128
rect 220169 86123 220235 86126
rect 267038 86124 267044 86126
rect 267108 86124 267114 86188
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect 86217 85506 86283 85509
rect 167821 85506 167887 85509
rect 86217 85504 167887 85506
rect 86217 85448 86222 85504
rect 86278 85448 167826 85504
rect 167882 85448 167887 85504
rect 86217 85446 167887 85448
rect 86217 85443 86283 85446
rect 167821 85443 167887 85446
rect 96337 85370 96403 85373
rect 173341 85370 173407 85373
rect 96337 85368 173407 85370
rect 96337 85312 96342 85368
rect 96398 85312 173346 85368
rect 173402 85312 173407 85368
rect 96337 85310 173407 85312
rect 96337 85307 96403 85310
rect 173341 85307 173407 85310
rect 120441 85234 120507 85237
rect 170581 85234 170647 85237
rect 120441 85232 170647 85234
rect 120441 85176 120446 85232
rect 120502 85176 170586 85232
rect 170642 85176 170647 85232
rect 120441 85174 170647 85176
rect 120441 85171 120507 85174
rect 170581 85171 170647 85174
rect 171869 84962 171935 84965
rect 205173 84962 205239 84965
rect 171869 84960 205239 84962
rect 171869 84904 171874 84960
rect 171930 84904 205178 84960
rect 205234 84904 205239 84960
rect 171869 84902 205239 84904
rect 171869 84899 171935 84902
rect 205173 84899 205239 84902
rect 181437 84826 181503 84829
rect 264605 84826 264671 84829
rect 181437 84824 264671 84826
rect -960 84690 480 84780
rect 181437 84768 181442 84824
rect 181498 84768 264610 84824
rect 264666 84768 264671 84824
rect 181437 84766 264671 84768
rect 181437 84763 181503 84766
rect 264605 84763 264671 84766
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 110229 84146 110295 84149
rect 204989 84146 205055 84149
rect 110229 84144 205055 84146
rect 110229 84088 110234 84144
rect 110290 84088 204994 84144
rect 205050 84088 205055 84144
rect 110229 84086 205055 84088
rect 110229 84083 110295 84086
rect 204989 84083 205055 84086
rect 124121 83466 124187 83469
rect 253289 83466 253355 83469
rect 124121 83464 253355 83466
rect 124121 83408 124126 83464
rect 124182 83408 253294 83464
rect 253350 83408 253355 83464
rect 124121 83406 253355 83408
rect 124121 83403 124187 83406
rect 253289 83403 253355 83406
rect 66069 82786 66135 82789
rect 213453 82786 213519 82789
rect 66069 82784 213519 82786
rect 66069 82728 66074 82784
rect 66130 82728 213458 82784
rect 213514 82728 213519 82784
rect 66069 82726 213519 82728
rect 66069 82723 66135 82726
rect 213453 82723 213519 82726
rect 99281 82106 99347 82109
rect 243813 82106 243879 82109
rect 99281 82104 243879 82106
rect 99281 82048 99286 82104
rect 99342 82048 243818 82104
rect 243874 82048 243879 82104
rect 99281 82046 243879 82048
rect 99281 82043 99347 82046
rect 243813 82043 243879 82046
rect 150433 81426 150499 81429
rect 166390 81426 166396 81428
rect 150433 81424 166396 81426
rect 150433 81368 150438 81424
rect 150494 81368 166396 81424
rect 150433 81366 166396 81368
rect 150433 81363 150499 81366
rect 166390 81364 166396 81366
rect 166460 81364 166466 81428
rect 142797 80882 142863 80885
rect 243721 80882 243787 80885
rect 142797 80880 243787 80882
rect 142797 80824 142802 80880
rect 142858 80824 243726 80880
rect 243782 80824 243787 80880
rect 142797 80822 243787 80824
rect 142797 80819 142863 80822
rect 243721 80819 243787 80822
rect 12341 80746 12407 80749
rect 259085 80746 259151 80749
rect 12341 80744 259151 80746
rect 12341 80688 12346 80744
rect 12402 80688 259090 80744
rect 259146 80688 259151 80744
rect 12341 80686 259151 80688
rect 12341 80683 12407 80686
rect 259085 80683 259151 80686
rect 106917 80066 106983 80069
rect 170489 80066 170555 80069
rect 106917 80064 170555 80066
rect 106917 80008 106922 80064
rect 106978 80008 170494 80064
rect 170550 80008 170555 80064
rect 106917 80006 170555 80008
rect 106917 80003 106983 80006
rect 170489 80003 170555 80006
rect 5441 79522 5507 79525
rect 224401 79522 224467 79525
rect 5441 79520 224467 79522
rect 5441 79464 5446 79520
rect 5502 79464 224406 79520
rect 224462 79464 224467 79520
rect 5441 79462 224467 79464
rect 5441 79459 5507 79462
rect 224401 79459 224467 79462
rect 29637 79386 29703 79389
rect 265893 79386 265959 79389
rect 29637 79384 265959 79386
rect 29637 79328 29642 79384
rect 29698 79328 265898 79384
rect 265954 79328 265959 79384
rect 29637 79326 265959 79328
rect 29637 79323 29703 79326
rect 265893 79323 265959 79326
rect 101949 78570 102015 78573
rect 207657 78570 207723 78573
rect 101949 78568 207723 78570
rect 101949 78512 101954 78568
rect 102010 78512 207662 78568
rect 207718 78512 207723 78568
rect 101949 78510 207723 78512
rect 101949 78507 102015 78510
rect 207657 78507 207723 78510
rect 67449 78434 67515 78437
rect 166206 78434 166212 78436
rect 67449 78432 166212 78434
rect 67449 78376 67454 78432
rect 67510 78376 166212 78432
rect 67449 78374 166212 78376
rect 67449 78371 67515 78374
rect 166206 78372 166212 78374
rect 166276 78372 166282 78436
rect 74441 77890 74507 77893
rect 260281 77890 260347 77893
rect 74441 77888 260347 77890
rect 74441 77832 74446 77888
rect 74502 77832 260286 77888
rect 260342 77832 260347 77888
rect 74441 77830 260347 77832
rect 74441 77827 74507 77830
rect 260281 77827 260347 77830
rect 70209 76666 70275 76669
rect 255957 76666 256023 76669
rect 70209 76664 256023 76666
rect 70209 76608 70214 76664
rect 70270 76608 255962 76664
rect 256018 76608 256023 76664
rect 70209 76606 256023 76608
rect 70209 76603 70275 76606
rect 255957 76603 256023 76606
rect 26141 76530 26207 76533
rect 246573 76530 246639 76533
rect 26141 76528 246639 76530
rect 26141 76472 26146 76528
rect 26202 76472 246578 76528
rect 246634 76472 246639 76528
rect 26141 76470 246639 76472
rect 26141 76467 26207 76470
rect 246573 76467 246639 76470
rect 95141 75306 95207 75309
rect 258809 75306 258875 75309
rect 95141 75304 258875 75306
rect 95141 75248 95146 75304
rect 95202 75248 258814 75304
rect 258870 75248 258875 75304
rect 95141 75246 258875 75248
rect 95141 75243 95207 75246
rect 258809 75243 258875 75246
rect 41321 75170 41387 75173
rect 284293 75170 284359 75173
rect 41321 75168 284359 75170
rect 41321 75112 41326 75168
rect 41382 75112 284298 75168
rect 284354 75112 284359 75168
rect 41321 75110 284359 75112
rect 41321 75107 41387 75110
rect 284293 75107 284359 75110
rect 73061 73946 73127 73949
rect 256049 73946 256115 73949
rect 73061 73944 256115 73946
rect 73061 73888 73066 73944
rect 73122 73888 256054 73944
rect 256110 73888 256115 73944
rect 73061 73886 256115 73888
rect 73061 73883 73127 73886
rect 256049 73883 256115 73886
rect 41321 73810 41387 73813
rect 264421 73810 264487 73813
rect 41321 73808 264487 73810
rect 41321 73752 41326 73808
rect 41382 73752 264426 73808
rect 264482 73752 264487 73808
rect 41321 73750 264487 73752
rect 41321 73747 41387 73750
rect 264421 73747 264487 73750
rect 88977 73130 89043 73133
rect 171869 73130 171935 73133
rect 88977 73128 171935 73130
rect 88977 73072 88982 73128
rect 89038 73072 171874 73128
rect 171930 73072 171935 73128
rect 88977 73070 171935 73072
rect 88977 73067 89043 73070
rect 171869 73067 171935 73070
rect 583520 72994 584960 73084
rect 583342 72934 584960 72994
rect 583342 72858 583402 72934
rect 583520 72858 584960 72934
rect 583342 72844 584960 72858
rect 583342 72798 583586 72844
rect 583526 72722 583586 72798
rect 583845 72722 583911 72725
rect 583526 72720 583911 72722
rect 583526 72664 583850 72720
rect 583906 72664 583911 72720
rect 583526 72662 583911 72664
rect 583845 72659 583911 72662
rect 53741 72586 53807 72589
rect 278773 72586 278839 72589
rect 53741 72584 278839 72586
rect 53741 72528 53746 72584
rect 53802 72528 278778 72584
rect 278834 72528 278839 72584
rect 53741 72526 278839 72528
rect 53741 72523 53807 72526
rect 278773 72523 278839 72526
rect 17861 72450 17927 72453
rect 263133 72450 263199 72453
rect 17861 72448 263199 72450
rect 17861 72392 17866 72448
rect 17922 72392 263138 72448
rect 263194 72392 263199 72448
rect 17861 72390 263199 72392
rect 17861 72387 17927 72390
rect 263133 72387 263199 72390
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 104157 71226 104223 71229
rect 213269 71226 213335 71229
rect 104157 71224 213335 71226
rect 104157 71168 104162 71224
rect 104218 71168 213274 71224
rect 213330 71168 213335 71224
rect 104157 71166 213335 71168
rect 104157 71163 104223 71166
rect 213269 71163 213335 71166
rect 61929 71090 61995 71093
rect 255313 71090 255379 71093
rect 61929 71088 255379 71090
rect 61929 71032 61934 71088
rect 61990 71032 255318 71088
rect 255374 71032 255379 71088
rect 61929 71030 255379 71032
rect 61929 71027 61995 71030
rect 255313 71027 255379 71030
rect 64413 69730 64479 69733
rect 262213 69730 262279 69733
rect 64413 69728 262279 69730
rect 64413 69672 64418 69728
rect 64474 69672 262218 69728
rect 262274 69672 262279 69728
rect 64413 69670 262279 69672
rect 64413 69667 64479 69670
rect 262213 69667 262279 69670
rect 23381 69594 23447 69597
rect 261661 69594 261727 69597
rect 23381 69592 261727 69594
rect 23381 69536 23386 69592
rect 23442 69536 261666 69592
rect 261722 69536 261727 69592
rect 23381 69534 261727 69536
rect 23381 69531 23447 69534
rect 261661 69531 261727 69534
rect 130377 68506 130443 68509
rect 168414 68506 168420 68508
rect 130377 68504 168420 68506
rect 130377 68448 130382 68504
rect 130438 68448 168420 68504
rect 130377 68446 168420 68448
rect 130377 68443 130443 68446
rect 168414 68444 168420 68446
rect 168484 68444 168490 68508
rect 160737 68370 160803 68373
rect 239489 68370 239555 68373
rect 160737 68368 239555 68370
rect 160737 68312 160742 68368
rect 160798 68312 239494 68368
rect 239550 68312 239555 68368
rect 160737 68310 239555 68312
rect 160737 68307 160803 68310
rect 239489 68307 239555 68310
rect 4061 68234 4127 68237
rect 224902 68234 224908 68236
rect 4061 68232 224908 68234
rect 4061 68176 4066 68232
rect 4122 68176 224908 68232
rect 4061 68174 224908 68176
rect 4061 68171 4127 68174
rect 224902 68172 224908 68174
rect 224972 68172 224978 68236
rect 66110 66948 66116 67012
rect 66180 67010 66186 67012
rect 276013 67010 276079 67013
rect 66180 67008 276079 67010
rect 66180 66952 276018 67008
rect 276074 66952 276079 67008
rect 66180 66950 276079 66952
rect 66180 66948 66186 66950
rect 276013 66947 276079 66950
rect 35801 66874 35867 66877
rect 249149 66874 249215 66877
rect 35801 66872 249215 66874
rect 35801 66816 35806 66872
rect 35862 66816 249154 66872
rect 249210 66816 249215 66872
rect 35801 66814 249215 66816
rect 35801 66811 35867 66814
rect 249149 66811 249215 66814
rect 122097 65650 122163 65653
rect 265709 65650 265775 65653
rect 122097 65648 265775 65650
rect 122097 65592 122102 65648
rect 122158 65592 265714 65648
rect 265770 65592 265775 65648
rect 122097 65590 265775 65592
rect 122097 65587 122163 65590
rect 265709 65587 265775 65590
rect 56501 65514 56567 65517
rect 307753 65514 307819 65517
rect 56501 65512 307819 65514
rect 56501 65456 56506 65512
rect 56562 65456 307758 65512
rect 307814 65456 307819 65512
rect 56501 65454 307819 65456
rect 56501 65451 56567 65454
rect 307753 65451 307819 65454
rect 75821 64290 75887 64293
rect 257429 64290 257495 64293
rect 75821 64288 257495 64290
rect 75821 64232 75826 64288
rect 75882 64232 257434 64288
rect 257490 64232 257495 64288
rect 75821 64230 257495 64232
rect 75821 64227 75887 64230
rect 257429 64227 257495 64230
rect 40677 64154 40743 64157
rect 253381 64154 253447 64157
rect 40677 64152 253447 64154
rect 40677 64096 40682 64152
rect 40738 64096 253386 64152
rect 253442 64096 253447 64152
rect 40677 64094 253447 64096
rect 40677 64091 40743 64094
rect 253381 64091 253447 64094
rect 87597 62930 87663 62933
rect 265617 62930 265683 62933
rect 87597 62928 265683 62930
rect 87597 62872 87602 62928
rect 87658 62872 265622 62928
rect 265678 62872 265683 62928
rect 87597 62870 265683 62872
rect 87597 62867 87663 62870
rect 265617 62867 265683 62870
rect 33041 62794 33107 62797
rect 261569 62794 261635 62797
rect 33041 62792 261635 62794
rect 33041 62736 33046 62792
rect 33102 62736 261574 62792
rect 261630 62736 261635 62792
rect 33041 62734 261635 62736
rect 33041 62731 33107 62734
rect 261569 62731 261635 62734
rect 86861 61570 86927 61573
rect 247677 61570 247743 61573
rect 86861 61568 247743 61570
rect 86861 61512 86866 61568
rect 86922 61512 247682 61568
rect 247738 61512 247743 61568
rect 86861 61510 247743 61512
rect 86861 61507 86927 61510
rect 247677 61507 247743 61510
rect 66161 61434 66227 61437
rect 262949 61434 263015 61437
rect 66161 61432 263015 61434
rect 66161 61376 66166 61432
rect 66222 61376 262954 61432
rect 263010 61376 263015 61432
rect 66161 61374 263015 61376
rect 66161 61371 66227 61374
rect 262949 61371 263015 61374
rect 583753 60210 583819 60213
rect 583710 60208 583819 60210
rect 583710 60152 583758 60208
rect 583814 60152 583819 60208
rect 583710 60147 583819 60152
rect 15101 59938 15167 59941
rect 264094 59938 264100 59940
rect 15101 59936 264100 59938
rect 15101 59880 15106 59936
rect 15162 59880 264100 59936
rect 15101 59878 264100 59880
rect 15101 59875 15167 59878
rect 264094 59876 264100 59878
rect 264164 59876 264170 59940
rect 583710 59802 583770 60147
rect 583342 59756 583770 59802
rect 583342 59742 584960 59756
rect 583342 59666 583402 59742
rect 583520 59666 584960 59742
rect 583342 59606 584960 59666
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 89621 58578 89687 58581
rect 267774 58578 267780 58580
rect 89621 58576 267780 58578
rect 89621 58520 89626 58576
rect 89682 58520 267780 58576
rect 89621 58518 267780 58520
rect 89621 58515 89687 58518
rect 267774 58516 267780 58518
rect 267844 58516 267850 58580
rect 57881 57218 57947 57221
rect 347037 57218 347103 57221
rect 57881 57216 347103 57218
rect 57881 57160 57886 57216
rect 57942 57160 347042 57216
rect 347098 57160 347103 57216
rect 57881 57158 347103 57160
rect 57881 57155 57947 57158
rect 347037 57155 347103 57158
rect 53741 55858 53807 55861
rect 245009 55858 245075 55861
rect 53741 55856 245075 55858
rect 53741 55800 53746 55856
rect 53802 55800 245014 55856
rect 245070 55800 245075 55856
rect 53741 55798 245075 55800
rect 53741 55795 53807 55798
rect 245009 55795 245075 55798
rect 50889 54498 50955 54501
rect 266854 54498 266860 54500
rect 50889 54496 266860 54498
rect 50889 54440 50894 54496
rect 50950 54440 266860 54496
rect 50889 54438 266860 54440
rect 50889 54435 50955 54438
rect 266854 54436 266860 54438
rect 266924 54436 266930 54500
rect 68921 53138 68987 53141
rect 242014 53138 242020 53140
rect 68921 53136 242020 53138
rect 68921 53080 68926 53136
rect 68982 53080 242020 53136
rect 68921 53078 242020 53080
rect 68921 53075 68987 53078
rect 242014 53076 242020 53078
rect 242084 53076 242090 53140
rect 57881 51778 57947 51781
rect 216213 51778 216279 51781
rect 57881 51776 216279 51778
rect 57881 51720 57886 51776
rect 57942 51720 216218 51776
rect 216274 51720 216279 51776
rect 57881 51718 216279 51720
rect 57881 51715 57947 51718
rect 216213 51715 216279 51718
rect 221457 50418 221523 50421
rect 267958 50418 267964 50420
rect 221457 50416 267964 50418
rect 221457 50360 221462 50416
rect 221518 50360 267964 50416
rect 221457 50358 267964 50360
rect 221457 50355 221523 50358
rect 267958 50356 267964 50358
rect 268028 50356 268034 50420
rect 22001 50282 22067 50285
rect 227069 50282 227135 50285
rect 22001 50280 227135 50282
rect 22001 50224 22006 50280
rect 22062 50224 227074 50280
rect 227130 50224 227135 50280
rect 22001 50222 227135 50224
rect 22001 50219 22067 50222
rect 227069 50219 227135 50222
rect 34421 47562 34487 47565
rect 246389 47562 246455 47565
rect 34421 47560 246455 47562
rect 34421 47504 34426 47560
rect 34482 47504 246394 47560
rect 246450 47504 246455 47560
rect 34421 47502 246455 47504
rect 34421 47499 34487 47502
rect 246389 47499 246455 47502
rect 582833 46338 582899 46341
rect 583520 46338 584960 46428
rect 582833 46336 584960 46338
rect 582833 46280 582838 46336
rect 582894 46280 584960 46336
rect 582833 46278 584960 46280
rect 582833 46275 582899 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 37181 44842 37247 44845
rect 244917 44842 244983 44845
rect 37181 44840 244983 44842
rect 37181 44784 37186 44840
rect 37242 44784 244922 44840
rect 244978 44784 244983 44840
rect 37181 44782 244983 44784
rect 37181 44779 37247 44782
rect 244917 44779 244983 44782
rect 16481 43482 16547 43485
rect 220854 43482 220860 43484
rect 16481 43480 220860 43482
rect 16481 43424 16486 43480
rect 16542 43424 220860 43480
rect 16481 43422 220860 43424
rect 16481 43419 16547 43422
rect 220854 43420 220860 43422
rect 220924 43420 220930 43484
rect 106917 42122 106983 42125
rect 264237 42122 264303 42125
rect 106917 42120 264303 42122
rect 106917 42064 106922 42120
rect 106978 42064 264242 42120
rect 264298 42064 264303 42120
rect 106917 42062 264303 42064
rect 106917 42059 106983 42062
rect 264237 42059 264303 42062
rect 81341 40626 81407 40629
rect 240726 40626 240732 40628
rect 81341 40624 240732 40626
rect 81341 40568 81346 40624
rect 81402 40568 240732 40624
rect 81341 40566 240732 40568
rect 81341 40563 81407 40566
rect 240726 40564 240732 40566
rect 240796 40564 240802 40628
rect 197997 39266 198063 39269
rect 276105 39266 276171 39269
rect 197997 39264 276171 39266
rect 197997 39208 198002 39264
rect 198058 39208 276110 39264
rect 276166 39208 276171 39264
rect 197997 39206 276171 39208
rect 197997 39203 198063 39206
rect 276105 39203 276171 39206
rect 10961 35186 11027 35189
rect 232497 35186 232563 35189
rect 10961 35184 232563 35186
rect 10961 35128 10966 35184
rect 11022 35128 232502 35184
rect 232558 35128 232563 35184
rect 10961 35126 232563 35128
rect 10961 35123 11027 35126
rect 232497 35123 232563 35126
rect 182817 33826 182883 33829
rect 244273 33826 244339 33829
rect 182817 33824 244339 33826
rect 182817 33768 182822 33824
rect 182878 33768 244278 33824
rect 244334 33768 244339 33824
rect 182817 33766 244339 33768
rect 182817 33763 182883 33766
rect 244273 33763 244339 33766
rect 582741 33146 582807 33149
rect 583520 33146 584960 33236
rect 582741 33144 584960 33146
rect 582741 33088 582746 33144
rect 582802 33088 584960 33144
rect 582741 33086 584960 33088
rect 582741 33083 582807 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 24761 29610 24827 29613
rect 255814 29610 255820 29612
rect 24761 29608 255820 29610
rect 24761 29552 24766 29608
rect 24822 29552 255820 29608
rect 24761 29550 255820 29552
rect 24761 29547 24827 29550
rect 255814 29548 255820 29550
rect 255884 29548 255890 29612
rect 3969 28250 4035 28253
rect 260046 28250 260052 28252
rect 3969 28248 260052 28250
rect 3969 28192 3974 28248
rect 4030 28192 260052 28248
rect 3969 28190 260052 28192
rect 3969 28187 4035 28190
rect 260046 28188 260052 28190
rect 260116 28188 260122 28252
rect 46841 26890 46907 26893
rect 225597 26890 225663 26893
rect 46841 26888 225663 26890
rect 46841 26832 46846 26888
rect 46902 26832 225602 26888
rect 225658 26832 225663 26888
rect 46841 26830 225663 26832
rect 46841 26827 46907 26830
rect 225597 26827 225663 26830
rect 59261 24170 59327 24173
rect 311893 24170 311959 24173
rect 59261 24168 311959 24170
rect 59261 24112 59266 24168
rect 59322 24112 311898 24168
rect 311954 24112 311959 24168
rect 59261 24110 311959 24112
rect 59261 24107 59327 24110
rect 311893 24107 311959 24110
rect 105 22674 171 22677
rect 227662 22674 227668 22676
rect 105 22672 227668 22674
rect 105 22616 110 22672
rect 166 22616 227668 22672
rect 105 22614 227668 22616
rect 105 22611 171 22614
rect 227662 22612 227668 22614
rect 227732 22612 227738 22676
rect 185577 21314 185643 21317
rect 259453 21314 259519 21317
rect 185577 21312 259519 21314
rect 185577 21256 185582 21312
rect 185638 21256 259458 21312
rect 259514 21256 259519 21312
rect 185577 21254 259519 21256
rect 185577 21251 185643 21254
rect 259453 21251 259519 21254
rect 583845 20362 583911 20365
rect 583710 20360 583911 20362
rect 583710 20304 583850 20360
rect 583906 20304 583911 20360
rect 583710 20302 583911 20304
rect 583710 19954 583770 20302
rect 583845 20299 583911 20302
rect 583342 19908 583770 19954
rect 583342 19894 584960 19908
rect 583342 19818 583402 19894
rect 583520 19818 584960 19894
rect 583342 19758 584960 19818
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 193857 15874 193923 15877
rect 269757 15874 269823 15877
rect 193857 15872 269823 15874
rect 193857 15816 193862 15872
rect 193918 15816 269762 15872
rect 269818 15816 269823 15872
rect 193857 15814 269823 15816
rect 193857 15811 193923 15814
rect 269757 15811 269823 15814
rect 186814 14452 186820 14516
rect 186884 14514 186890 14516
rect 269665 14514 269731 14517
rect 186884 14512 269731 14514
rect 186884 14456 269670 14512
rect 269726 14456 269731 14512
rect 186884 14454 269731 14456
rect 186884 14452 186890 14454
rect 269665 14451 269731 14454
rect 188337 13018 188403 13021
rect 261753 13018 261819 13021
rect 188337 13016 261819 13018
rect 188337 12960 188342 13016
rect 188398 12960 261758 13016
rect 261814 12960 261819 13016
rect 188337 12958 261819 12960
rect 188337 12955 188403 12958
rect 261753 12955 261819 12958
rect 136449 11658 136515 11661
rect 169702 11658 169708 11660
rect 136449 11656 169708 11658
rect 136449 11600 136454 11656
rect 136510 11600 169708 11656
rect 136449 11598 169708 11600
rect 136449 11595 136515 11598
rect 169702 11596 169708 11598
rect 169772 11596 169778 11660
rect 195094 11596 195100 11660
rect 195164 11658 195170 11660
rect 268377 11658 268443 11661
rect 195164 11656 268443 11658
rect 195164 11600 268382 11656
rect 268438 11600 268443 11656
rect 195164 11598 268443 11600
rect 195164 11596 195170 11598
rect 268377 11595 268443 11598
rect 9581 10298 9647 10301
rect 160737 10298 160803 10301
rect 9581 10296 160803 10298
rect 9581 10240 9586 10296
rect 9642 10240 160742 10296
rect 160798 10240 160803 10296
rect 9581 10238 160803 10240
rect 9581 10235 9647 10238
rect 160737 10235 160803 10238
rect 184197 10298 184263 10301
rect 244089 10298 244155 10301
rect 184197 10296 244155 10298
rect 184197 10240 184202 10296
rect 184258 10240 244094 10296
rect 244150 10240 244155 10296
rect 184197 10238 244155 10240
rect 184197 10235 184263 10238
rect 244089 10235 244155 10238
rect 132953 8938 133019 8941
rect 166942 8938 166948 8940
rect 132953 8936 166948 8938
rect 132953 8880 132958 8936
rect 133014 8880 166948 8936
rect 132953 8878 166948 8880
rect 132953 8875 133019 8878
rect 166942 8876 166948 8878
rect 167012 8876 167018 8940
rect 173014 8876 173020 8940
rect 173084 8938 173090 8940
rect 281441 8938 281507 8941
rect 173084 8936 281507 8938
rect 173084 8880 281446 8936
rect 281502 8880 281507 8936
rect 173084 8878 281507 8880
rect 173084 8876 173090 8878
rect 281441 8875 281507 8878
rect 227069 7578 227135 7581
rect 298461 7578 298527 7581
rect 227069 7576 298527 7578
rect 227069 7520 227074 7576
rect 227130 7520 298466 7576
rect 298522 7520 298527 7576
rect 227069 7518 298527 7520
rect 227069 7515 227135 7518
rect 298461 7515 298527 7518
rect 13 6762 79 6765
rect 13 6760 122 6762
rect 13 6704 18 6760
rect 74 6704 122 6760
rect 13 6699 122 6704
rect 62 6626 122 6699
rect 582649 6626 582715 6629
rect 583520 6626 584960 6716
rect 62 6580 674 6626
rect -960 6566 674 6580
rect -960 6490 480 6566
rect 614 6490 674 6566
rect 582649 6624 584960 6626
rect 582649 6568 582654 6624
rect 582710 6568 584960 6624
rect 582649 6566 584960 6568
rect 582649 6563 582715 6566
rect -960 6430 674 6490
rect 583520 6476 584960 6566
rect -960 6340 480 6430
rect 39573 6218 39639 6221
rect 211797 6218 211863 6221
rect 39573 6216 211863 6218
rect 39573 6160 39578 6216
rect 39634 6160 211802 6216
rect 211858 6160 211863 6216
rect 39573 6158 211863 6160
rect 39573 6155 39639 6158
rect 211797 6155 211863 6158
rect 220077 6218 220143 6221
rect 239305 6218 239371 6221
rect 220077 6216 239371 6218
rect 220077 6160 220082 6216
rect 220138 6160 239310 6216
rect 239366 6160 239371 6216
rect 220077 6158 239371 6160
rect 220077 6155 220143 6158
rect 239305 6155 239371 6158
rect 278313 6218 278379 6221
rect 304993 6218 305059 6221
rect 278313 6216 305059 6218
rect 278313 6160 278318 6216
rect 278374 6160 304998 6216
rect 305054 6160 305059 6216
rect 278313 6158 305059 6160
rect 278313 6155 278379 6158
rect 304993 6155 305059 6158
rect 177246 4932 177252 4996
rect 177316 4994 177322 4996
rect 242893 4994 242959 4997
rect 177316 4992 242959 4994
rect 177316 4936 242898 4992
rect 242954 4936 242959 4992
rect 177316 4934 242959 4936
rect 177316 4932 177322 4934
rect 242893 4931 242959 4934
rect 178677 4858 178743 4861
rect 265341 4858 265407 4861
rect 178677 4856 265407 4858
rect 178677 4800 178682 4856
rect 178738 4800 265346 4856
rect 265402 4800 265407 4856
rect 178677 4798 265407 4800
rect 178677 4795 178743 4798
rect 265341 4795 265407 4798
rect 253054 3980 253060 4044
rect 253124 4042 253130 4044
rect 260649 4042 260715 4045
rect 253124 4040 260715 4042
rect 253124 3984 260654 4040
rect 260710 3984 260715 4040
rect 253124 3982 260715 3984
rect 253124 3980 253130 3982
rect 260649 3979 260715 3982
rect 246246 3436 246252 3500
rect 246316 3498 246322 3500
rect 247585 3498 247651 3501
rect 246316 3496 247651 3498
rect 246316 3440 247590 3496
rect 247646 3440 247651 3496
rect 246316 3438 247651 3440
rect 246316 3436 246322 3438
rect 247585 3435 247651 3438
rect 249006 3436 249012 3500
rect 249076 3498 249082 3500
rect 252369 3498 252435 3501
rect 249076 3496 252435 3498
rect 249076 3440 252374 3496
rect 252430 3440 252435 3496
rect 249076 3438 252435 3440
rect 249076 3436 249082 3438
rect 252369 3435 252435 3438
rect 285622 3436 285628 3500
rect 285692 3498 285698 3500
rect 286593 3498 286659 3501
rect 285692 3496 286659 3498
rect 285692 3440 286598 3496
rect 286654 3440 286659 3496
rect 285692 3438 286659 3440
rect 285692 3436 285698 3438
rect 286593 3435 286659 3438
rect 287094 3436 287100 3500
rect 287164 3498 287170 3500
rect 287789 3498 287855 3501
rect 287164 3496 287855 3498
rect 287164 3440 287794 3496
rect 287850 3440 287855 3496
rect 287164 3438 287855 3440
rect 287164 3436 287170 3438
rect 287789 3435 287855 3438
rect 288382 3436 288388 3500
rect 288452 3498 288458 3500
rect 288985 3498 289051 3501
rect 288452 3496 289051 3498
rect 288452 3440 288990 3496
rect 289046 3440 289051 3496
rect 288452 3438 289051 3440
rect 288452 3436 288458 3438
rect 288985 3435 289051 3438
rect 291142 3436 291148 3500
rect 291212 3498 291218 3500
rect 291377 3498 291443 3501
rect 291212 3496 291443 3498
rect 291212 3440 291382 3496
rect 291438 3440 291443 3496
rect 291212 3438 291443 3440
rect 291212 3436 291218 3438
rect 291377 3435 291443 3438
rect 298686 3436 298692 3500
rect 298756 3498 298762 3500
rect 300761 3498 300827 3501
rect 298756 3496 300827 3498
rect 298756 3440 300766 3496
rect 300822 3440 300827 3496
rect 298756 3438 300827 3440
rect 298756 3436 298762 3438
rect 300761 3435 300827 3438
rect 348049 3498 348115 3501
rect 357433 3498 357499 3501
rect 348049 3496 357499 3498
rect 348049 3440 348054 3496
rect 348110 3440 357438 3496
rect 357494 3440 357499 3496
rect 348049 3438 357499 3440
rect 348049 3435 348115 3438
rect 357433 3435 357499 3438
rect 64321 3362 64387 3365
rect 122097 3362 122163 3365
rect 64321 3360 122163 3362
rect 64321 3304 64326 3360
rect 64382 3304 122102 3360
rect 122158 3304 122163 3360
rect 64321 3302 122163 3304
rect 64321 3299 64387 3302
rect 122097 3299 122163 3302
rect 125869 3362 125935 3365
rect 191046 3362 191052 3364
rect 125869 3360 191052 3362
rect 125869 3304 125874 3360
rect 125930 3304 191052 3360
rect 125869 3302 191052 3304
rect 125869 3299 125935 3302
rect 191046 3300 191052 3302
rect 191116 3300 191122 3364
rect 196617 3362 196683 3365
rect 246389 3362 246455 3365
rect 196617 3360 246455 3362
rect 196617 3304 196622 3360
rect 196678 3304 246394 3360
rect 246450 3304 246455 3360
rect 196617 3302 246455 3304
rect 196617 3299 196683 3302
rect 246389 3299 246455 3302
rect 294873 3362 294939 3365
rect 299749 3362 299815 3365
rect 294873 3360 299815 3362
rect 294873 3304 294878 3360
rect 294934 3304 299754 3360
rect 299810 3304 299815 3360
rect 294873 3302 299815 3304
rect 294873 3299 294939 3302
rect 299749 3299 299815 3302
rect 344553 3362 344619 3365
rect 356053 3362 356119 3365
rect 344553 3360 356119 3362
rect 344553 3304 344558 3360
rect 344614 3304 356058 3360
rect 356114 3304 356119 3360
rect 344553 3302 356119 3304
rect 344553 3299 344619 3302
rect 356053 3299 356119 3302
rect 200849 2002 200915 2005
rect 254669 2002 254735 2005
rect 200849 2000 254735 2002
rect 200849 1944 200854 2000
rect 200910 1944 254674 2000
rect 254730 1944 254735 2000
rect 200849 1942 254735 1944
rect 200849 1939 200915 1942
rect 254669 1939 254735 1942
<< via3 >>
rect 69612 702476 69676 702540
rect 76052 699756 76116 699820
rect 93900 589460 93964 589524
rect 88196 588508 88260 588572
rect 67772 583748 67836 583812
rect 69428 582252 69492 582316
rect 122972 581572 123036 581636
rect 119476 580212 119540 580276
rect 111012 553420 111076 553484
rect 66668 550836 66732 550900
rect 99972 550700 100036 550764
rect 107700 542948 107764 543012
rect 76052 539548 76116 539612
rect 115060 538596 115124 538660
rect 68140 535468 68204 535532
rect 69612 535528 69676 535532
rect 69612 535472 69662 535528
rect 69662 535472 69676 535528
rect 69612 535468 69676 535472
rect 71820 535468 71884 535532
rect 106412 465700 106476 465764
rect 102180 464340 102244 464404
rect 89668 462844 89732 462908
rect 104940 462844 105004 462908
rect 115980 462844 116044 462908
rect 109172 462164 109236 462228
rect 88196 460124 88260 460188
rect 98132 458764 98196 458828
rect 96660 457404 96724 457468
rect 100708 456044 100772 456108
rect 92612 454684 92676 454748
rect 67772 453868 67836 453932
rect 68324 453868 68388 453932
rect 91324 453188 91388 453252
rect 68324 452644 68388 452708
rect 158668 451284 158732 451348
rect 111748 448564 111812 448628
rect 120028 447884 120092 447948
rect 95188 447748 95252 447812
rect 122604 447748 122668 447812
rect 155172 445980 155236 446044
rect 91140 445708 91204 445772
rect 93900 445708 93964 445772
rect 96476 445708 96540 445772
rect 97764 445708 97828 445772
rect 111564 445708 111628 445772
rect 114324 445708 114388 445772
rect 118556 445708 118620 445772
rect 109540 444816 109604 444820
rect 109540 444760 109554 444816
rect 109554 444760 109604 444816
rect 109540 444756 109604 444760
rect 133092 442308 133156 442372
rect 68324 440812 68388 440876
rect 122972 435236 123036 435300
rect 146892 435236 146956 435300
rect 120028 431428 120092 431492
rect 122604 430884 122668 430948
rect 122420 426260 122484 426324
rect 66116 424084 66180 424148
rect 122420 422316 122484 422380
rect 122788 422316 122852 422380
rect 122788 422044 122852 422108
rect 69244 419324 69308 419388
rect 122788 412856 122852 412860
rect 122788 412800 122802 412856
rect 122802 412800 122852 412856
rect 122788 412796 122852 412800
rect 122788 412388 122852 412452
rect 66668 411300 66732 411364
rect 122788 403064 122852 403068
rect 122788 403008 122802 403064
rect 122802 403008 122852 403064
rect 122788 403004 122852 403008
rect 122972 402868 123036 402932
rect 122972 394708 123036 394772
rect 122788 393408 122852 393412
rect 122788 393352 122802 393408
rect 122802 393352 122852 393408
rect 122788 393348 122852 393352
rect 122788 393272 122852 393276
rect 122788 393216 122802 393272
rect 122802 393216 122852 393272
rect 122788 393212 122852 393216
rect 92612 390900 92676 390964
rect 102180 390960 102244 390964
rect 102180 390904 102194 390960
rect 102194 390904 102244 390960
rect 102180 390900 102244 390904
rect 69612 390628 69676 390692
rect 71820 390416 71884 390420
rect 71820 390360 71870 390416
rect 71870 390360 71884 390416
rect 71820 390356 71884 390360
rect 91324 390416 91388 390420
rect 91324 390360 91374 390416
rect 91374 390360 91388 390416
rect 91324 390356 91388 390360
rect 95188 390356 95252 390420
rect 96660 390356 96724 390420
rect 98132 390356 98196 390420
rect 100708 390416 100772 390420
rect 100708 390360 100722 390416
rect 100722 390360 100772 390416
rect 100708 390356 100772 390360
rect 104940 390416 105004 390420
rect 104940 390360 104990 390416
rect 104990 390360 105004 390416
rect 104940 390356 105004 390360
rect 106412 390356 106476 390420
rect 107700 390356 107764 390420
rect 109172 390356 109236 390420
rect 115980 390416 116044 390420
rect 115980 390360 115994 390416
rect 115994 390360 116044 390416
rect 115980 390356 116044 390360
rect 120028 390356 120092 390420
rect 111012 389132 111076 389196
rect 76420 388996 76484 389060
rect 89668 388996 89732 389060
rect 111748 388996 111812 389060
rect 67772 388724 67836 388788
rect 68140 388724 68204 388788
rect 96476 388452 96540 388516
rect 99972 388316 100036 388380
rect 83412 387228 83476 387292
rect 122972 385596 123036 385660
rect 122788 383828 122852 383892
rect 122788 383616 122852 383620
rect 122788 383560 122802 383616
rect 122802 383560 122852 383616
rect 122788 383556 122852 383560
rect 115060 382256 115124 382260
rect 115060 382200 115110 382256
rect 115110 382200 115124 382256
rect 115060 382196 115124 382200
rect 89668 378796 89732 378860
rect 136588 378660 136652 378724
rect 163452 377300 163516 377364
rect 122788 374172 122852 374236
rect 122788 373960 122852 373964
rect 122788 373904 122802 373960
rect 122802 373904 122852 373960
rect 122788 373900 122852 373904
rect 244228 371316 244292 371380
rect 114324 369956 114388 370020
rect 97764 369820 97828 369884
rect 252508 369820 252572 369884
rect 169708 369004 169772 369068
rect 69796 367644 69860 367708
rect 69060 366284 69124 366348
rect 146892 365876 146956 365940
rect 222332 365740 222396 365804
rect 122972 364516 123036 364580
rect 122972 364108 123036 364172
rect 138060 362204 138124 362268
rect 111564 361796 111628 361860
rect 122604 361660 122668 361724
rect 70164 360844 70228 360908
rect 66116 359348 66180 359412
rect 91140 359272 91204 359276
rect 91140 359216 91190 359272
rect 91190 359216 91204 359272
rect 91140 359212 91204 359216
rect 109540 358940 109604 359004
rect 136036 357988 136100 358052
rect 188292 357580 188356 357644
rect 249748 357444 249812 357508
rect 111748 356628 111812 356692
rect 197860 356220 197924 356284
rect 212580 354860 212644 354924
rect 232452 354724 232516 354788
rect 139716 352548 139780 352612
rect 186820 350644 186884 350708
rect 248460 350508 248524 350572
rect 196940 349284 197004 349348
rect 69612 349148 69676 349212
rect 70164 349148 70228 349212
rect 66668 349012 66732 349076
rect 66668 347788 66732 347852
rect 118556 347652 118620 347716
rect 156460 347108 156524 347172
rect 67956 345748 68020 345812
rect 67772 345612 67836 345676
rect 230428 340988 230492 341052
rect 291148 339492 291212 339556
rect 93900 332420 93964 332484
rect 160692 331468 160756 331532
rect 61884 329972 61948 330036
rect 154252 329972 154316 330036
rect 153700 327660 153764 327724
rect 82676 327524 82740 327588
rect 145604 327116 145668 327180
rect 150388 327116 150452 327180
rect 155356 327116 155420 327180
rect 67404 326980 67468 327044
rect 160876 326436 160940 326500
rect 237420 324940 237484 325004
rect 154252 320724 154316 320788
rect 155172 318548 155236 318612
rect 155356 318140 155420 318204
rect 191604 317324 191668 317388
rect 66668 316372 66732 316436
rect 191604 316100 191668 316164
rect 69428 315556 69492 315620
rect 154252 315012 154316 315076
rect 160692 313924 160756 313988
rect 195100 313244 195164 313308
rect 284340 311884 284404 311948
rect 160876 311068 160940 311132
rect 187004 308484 187068 308548
rect 214236 308348 214300 308412
rect 67404 307940 67468 308004
rect 242940 306444 243004 306508
rect 67772 297332 67836 297396
rect 241652 297332 241716 297396
rect 221044 296788 221108 296852
rect 180012 295972 180076 296036
rect 158668 295352 158732 295356
rect 158668 295296 158682 295352
rect 158682 295296 158732 295352
rect 158668 295292 158732 295296
rect 69060 295020 69124 295084
rect 166212 292572 166276 292636
rect 199332 291348 199396 291412
rect 156460 291076 156524 291140
rect 280292 289988 280356 290052
rect 200620 288628 200684 288692
rect 233188 288628 233252 288692
rect 288572 288492 288636 288556
rect 287284 287268 287348 287332
rect 211660 287132 211724 287196
rect 226932 285908 226996 285972
rect 240364 285908 240428 285972
rect 238524 285772 238588 285836
rect 224908 285636 224972 285700
rect 236500 285636 236564 285700
rect 281580 284412 281644 284476
rect 205404 283928 205468 283932
rect 205404 283872 205418 283928
rect 205418 283872 205468 283928
rect 205404 283868 205468 283872
rect 206876 283868 206940 283932
rect 209636 283868 209700 283932
rect 214052 283928 214116 283932
rect 214052 283872 214102 283928
rect 214102 283872 214116 283928
rect 214052 283868 214116 283872
rect 215340 283868 215404 283932
rect 217180 283868 217244 283932
rect 224724 283928 224788 283932
rect 224724 283872 224738 283928
rect 224738 283872 224788 283928
rect 224724 283868 224788 283872
rect 226380 283868 226444 283932
rect 228772 283868 228836 283932
rect 229692 283868 229756 283932
rect 231716 283868 231780 283932
rect 236500 283868 236564 283932
rect 200068 282508 200132 282572
rect 197860 281556 197924 281620
rect 163452 280060 163516 280124
rect 199332 279516 199396 279580
rect 67956 279380 68020 279444
rect 243492 279108 243556 279172
rect 65932 275980 65996 276044
rect 155172 275300 155236 275364
rect 244228 275572 244292 275636
rect 173020 275164 173084 275228
rect 160692 273260 160756 273324
rect 273300 270540 273364 270604
rect 161980 269316 162044 269380
rect 67404 266868 67468 266932
rect 249932 265704 249996 265708
rect 249932 265648 249982 265704
rect 249982 265648 249996 265704
rect 249932 265644 249996 265648
rect 249748 263876 249812 263940
rect 154620 260748 154684 260812
rect 191052 260068 191116 260132
rect 191604 258980 191668 259044
rect 69428 256804 69492 256868
rect 67956 256260 68020 256324
rect 197124 255172 197188 255236
rect 66668 251908 66732 251972
rect 199884 251908 199948 251972
rect 168420 251364 168484 251428
rect 199516 249792 199580 249796
rect 199516 249736 199530 249792
rect 199530 249736 199580 249792
rect 199516 249732 199580 249736
rect 248460 249460 248524 249524
rect 187004 247148 187068 247212
rect 199884 246468 199948 246532
rect 160692 246196 160756 246260
rect 243492 246196 243556 246260
rect 69428 245108 69492 245172
rect 154436 244428 154500 244492
rect 66116 243476 66180 243540
rect 199884 243476 199948 243540
rect 195284 242932 195348 242996
rect 245884 242932 245948 242996
rect 67404 242796 67468 242860
rect 136036 242040 136100 242044
rect 136036 241984 136050 242040
rect 136050 241984 136100 242040
rect 136036 241980 136100 241984
rect 136588 241980 136652 242044
rect 138060 241980 138124 242044
rect 147444 241980 147508 242044
rect 83412 241300 83476 241364
rect 245700 240212 245764 240276
rect 214236 240076 214300 240140
rect 221044 240136 221108 240140
rect 221044 240080 221094 240136
rect 221094 240080 221108 240136
rect 221044 240076 221108 240080
rect 224908 240136 224972 240140
rect 224908 240080 224958 240136
rect 224958 240080 224972 240136
rect 224908 240076 224972 240080
rect 229692 240136 229756 240140
rect 229692 240080 229742 240136
rect 229742 240080 229756 240136
rect 229692 240076 229756 240080
rect 230428 240076 230492 240140
rect 237420 240076 237484 240140
rect 154436 239940 154500 240004
rect 199884 239396 199948 239460
rect 212580 238580 212644 238644
rect 222332 238580 222396 238644
rect 232452 238580 232516 238644
rect 241652 238580 241716 238644
rect 211660 238308 211724 238372
rect 200620 237900 200684 237964
rect 213132 237416 213196 237420
rect 213132 237360 213146 237416
rect 213146 237360 213196 237416
rect 213132 237356 213196 237360
rect 155172 237220 155236 237284
rect 196940 237220 197004 237284
rect 186820 237084 186884 237148
rect 180012 235724 180076 235788
rect 188292 235724 188356 235788
rect 195284 235180 195348 235244
rect 214052 234636 214116 234700
rect 245884 234500 245948 234564
rect 191052 234364 191116 234428
rect 252508 234500 252572 234564
rect 65932 233820 65996 233884
rect 231716 233140 231780 233204
rect 233372 233140 233436 233204
rect 139716 233004 139780 233068
rect 69612 232460 69676 232524
rect 242940 232460 243004 232524
rect 217180 231780 217244 231844
rect 76420 231644 76484 231708
rect 133092 231372 133156 231436
rect 69796 230420 69860 230484
rect 67956 229740 68020 229804
rect 61884 228380 61948 228444
rect 82676 227564 82740 227628
rect 245700 227564 245764 227628
rect 150388 224164 150452 224228
rect 285812 224164 285876 224228
rect 191052 222940 191116 223004
rect 155172 219132 155236 219196
rect 298692 218588 298756 218652
rect 209636 215868 209700 215932
rect 186820 214508 186884 214572
rect 215340 213828 215404 213892
rect 224724 213284 224788 213348
rect 213132 213148 213196 213212
rect 231900 211924 231964 211988
rect 155172 210292 155236 210356
rect 166212 210292 166276 210356
rect 66668 206212 66732 206276
rect 244228 205184 244292 205188
rect 244228 205128 244278 205184
rect 244278 205128 244292 205184
rect 244228 205124 244292 205128
rect 288388 202132 288452 202196
rect 253060 200636 253124 200700
rect 226932 196012 226996 196076
rect 234660 196012 234724 196076
rect 280292 195332 280356 195396
rect 287100 193836 287164 193900
rect 229692 191116 229756 191180
rect 226380 189892 226444 189956
rect 161980 189756 162044 189820
rect 228220 189756 228284 189820
rect 240548 189756 240612 189820
rect 284524 189620 284588 189684
rect 241468 188532 241532 188596
rect 232084 188396 232148 188460
rect 251220 187172 251284 187236
rect 244412 187036 244476 187100
rect 295380 186900 295444 186964
rect 145604 185676 145668 185740
rect 177252 185676 177316 185740
rect 206876 185676 206940 185740
rect 227668 185676 227732 185740
rect 228772 185676 228836 185740
rect 246252 185540 246316 185604
rect 290596 185540 290660 185604
rect 67772 184180 67836 184244
rect 249012 182956 249076 183020
rect 230428 181596 230492 181660
rect 237604 181460 237668 181524
rect 291332 181460 291396 181524
rect 285628 181324 285692 181388
rect 199516 178740 199580 178804
rect 278820 178604 278884 178668
rect 109540 178332 109604 178396
rect 110644 178196 110708 178260
rect 97028 177924 97092 177988
rect 98316 177516 98380 177580
rect 101996 177576 102060 177580
rect 101996 177520 102046 177576
rect 102046 177520 102060 177576
rect 101996 177516 102060 177520
rect 105676 177516 105740 177580
rect 108068 177516 108132 177580
rect 112116 177516 112180 177580
rect 120764 177516 120828 177580
rect 124444 177516 124508 177580
rect 125732 177516 125796 177580
rect 127020 177516 127084 177580
rect 132356 177576 132420 177580
rect 132356 177520 132406 177576
rect 132406 177520 132420 177576
rect 132356 177516 132420 177520
rect 133092 177516 133156 177580
rect 148180 177576 148244 177580
rect 148180 177520 148230 177576
rect 148230 177520 148244 177576
rect 148180 177516 148244 177520
rect 118372 177380 118436 177444
rect 283788 177380 283852 177444
rect 130700 177244 130764 177308
rect 104572 177108 104636 177172
rect 113220 176972 113284 177036
rect 115796 177032 115860 177036
rect 115796 176976 115846 177032
rect 115846 176976 115860 177032
rect 115796 176972 115860 176976
rect 279372 176972 279436 177036
rect 100708 176896 100772 176900
rect 100708 176840 100758 176896
rect 100758 176840 100772 176896
rect 100708 176836 100772 176840
rect 106964 176700 107028 176764
rect 121868 176760 121932 176764
rect 121868 176704 121918 176760
rect 121918 176704 121932 176760
rect 121868 176700 121932 176704
rect 123156 176700 123220 176764
rect 129412 176760 129476 176764
rect 129412 176704 129462 176760
rect 129462 176704 129476 176760
rect 129412 176700 129476 176704
rect 136036 176760 136100 176764
rect 136036 176704 136086 176760
rect 136086 176704 136100 176760
rect 136036 176700 136100 176704
rect 158852 176700 158916 176764
rect 229324 176700 229388 176764
rect 230612 176564 230676 176628
rect 99420 176428 99484 176492
rect 103284 176428 103348 176492
rect 128124 176428 128188 176492
rect 166948 175944 167012 175948
rect 166948 175888 166998 175944
rect 166998 175888 167012 175944
rect 166948 175884 167012 175888
rect 241652 176020 241716 176084
rect 273300 175944 273364 175948
rect 273300 175888 273350 175944
rect 273350 175888 273364 175944
rect 273300 175884 273364 175888
rect 114324 175476 114388 175540
rect 116900 175340 116964 175404
rect 229140 175128 229204 175132
rect 229140 175072 229154 175128
rect 229154 175072 229204 175128
rect 229140 175068 229204 175072
rect 229692 175068 229756 175132
rect 119398 174992 119462 174996
rect 119398 174936 119434 174992
rect 119434 174936 119462 174992
rect 119398 174932 119462 174936
rect 229508 174932 229572 174996
rect 134358 174796 134422 174860
rect 229140 174252 229204 174316
rect 240364 173844 240428 173908
rect 279372 173708 279436 173772
rect 238524 173300 238588 173364
rect 240364 172348 240428 172412
rect 237420 168676 237484 168740
rect 279372 168268 279436 168332
rect 236500 165140 236564 165204
rect 244412 162148 244476 162212
rect 231900 161468 231964 161532
rect 281580 157252 281644 157316
rect 244228 156708 244292 156772
rect 233556 155892 233620 155956
rect 230612 155756 230676 155820
rect 230980 155212 231044 155276
rect 233188 154804 233252 154868
rect 232084 152492 232148 152556
rect 249932 151948 249996 152012
rect 241468 150996 241532 151060
rect 230428 149636 230492 149700
rect 241836 149636 241900 149700
rect 237604 149228 237668 149292
rect 291332 149092 291396 149156
rect 240548 147188 240612 147252
rect 229324 146236 229388 146300
rect 233556 145284 233620 145348
rect 233740 145284 233804 145348
rect 283788 143516 283852 143580
rect 240364 143244 240428 143308
rect 244780 141340 244844 141404
rect 251220 140116 251284 140180
rect 260052 140116 260116 140180
rect 284340 140388 284404 140452
rect 231164 139980 231228 140044
rect 233372 139708 233436 139772
rect 234660 139164 234724 139228
rect 232452 138620 232516 138684
rect 229140 137260 229204 137324
rect 242204 135764 242268 135828
rect 280476 135900 280540 135964
rect 267780 135628 267844 135692
rect 250300 134404 250364 134468
rect 290596 133860 290660 133924
rect 230980 133452 231044 133516
rect 242020 132908 242084 132972
rect 229692 132772 229756 132836
rect 295380 132500 295444 132564
rect 231164 131548 231228 131612
rect 280292 131276 280356 131340
rect 266860 131004 266924 131068
rect 251772 128964 251836 129028
rect 255820 127196 255884 127260
rect 264100 127060 264164 127124
rect 240732 120804 240796 120868
rect 284524 116860 284588 116924
rect 262812 113732 262876 113796
rect 230980 111148 231044 111212
rect 250300 107476 250364 107540
rect 251772 106796 251836 106860
rect 288572 106252 288636 106316
rect 285812 106116 285876 106180
rect 233740 103260 233804 103324
rect 166212 102444 166276 102508
rect 287284 102172 287348 102236
rect 244780 102036 244844 102100
rect 267044 100812 267108 100876
rect 230980 98908 231044 98972
rect 262812 98636 262876 98700
rect 232452 97956 232516 98020
rect 267964 97956 268028 98020
rect 229140 97140 229204 97204
rect 229140 96596 229204 96660
rect 219204 95976 219268 95980
rect 219204 95920 219254 95976
rect 219254 95920 219268 95976
rect 219204 95916 219268 95920
rect 166396 95780 166460 95844
rect 219204 95840 219268 95844
rect 219204 95784 219218 95840
rect 219218 95784 219268 95840
rect 219204 95780 219268 95784
rect 224908 95508 224972 95572
rect 228588 95508 228652 95572
rect 205404 95100 205468 95164
rect 100630 94752 100694 94756
rect 100630 94696 100666 94752
rect 100666 94696 100694 94752
rect 100630 94692 100694 94696
rect 151308 94692 151372 94756
rect 151766 94692 151830 94756
rect 126652 94012 126716 94076
rect 111932 93876 111996 93940
rect 114876 93740 114940 93804
rect 134380 93604 134444 93668
rect 117084 93528 117148 93532
rect 117084 93472 117134 93528
rect 117134 93472 117148 93528
rect 117084 93468 117148 93472
rect 121684 93528 121748 93532
rect 121684 93472 121734 93528
rect 121734 93472 121748 93528
rect 121684 93468 121748 93472
rect 123156 93468 123220 93532
rect 133092 93332 133156 93396
rect 110092 93256 110156 93260
rect 110092 93200 110142 93256
rect 110142 93200 110156 93256
rect 110092 93196 110156 93200
rect 113772 93256 113836 93260
rect 113772 93200 113822 93256
rect 113822 93200 113836 93256
rect 113772 93196 113836 93200
rect 84332 92440 84396 92444
rect 84332 92384 84382 92440
rect 84382 92384 84396 92440
rect 84332 92380 84396 92384
rect 88932 92380 88996 92444
rect 99052 92440 99116 92444
rect 99052 92384 99102 92440
rect 99102 92384 99116 92440
rect 99052 92380 99116 92384
rect 106780 92440 106844 92444
rect 106780 92384 106830 92440
rect 106830 92384 106844 92440
rect 106780 92380 106844 92384
rect 109172 92380 109236 92444
rect 110644 92440 110708 92444
rect 110644 92384 110694 92440
rect 110694 92384 110708 92440
rect 110644 92380 110708 92384
rect 111196 92380 111260 92444
rect 124076 92440 124140 92444
rect 124076 92384 124126 92440
rect 124126 92384 124140 92440
rect 124076 92380 124140 92384
rect 136036 92440 136100 92444
rect 136036 92384 136086 92440
rect 136086 92384 136100 92440
rect 136036 92380 136100 92384
rect 151308 92380 151372 92444
rect 116716 92244 116780 92308
rect 130700 92108 130764 92172
rect 96292 91896 96356 91900
rect 96292 91840 96342 91896
rect 96342 91840 96356 91896
rect 96292 91836 96356 91840
rect 242204 91836 242268 91900
rect 92612 91700 92676 91764
rect 98132 91700 98196 91764
rect 119660 91700 119724 91764
rect 229692 91700 229756 91764
rect 104572 91564 104636 91628
rect 122788 91428 122852 91492
rect 96660 91292 96724 91356
rect 101812 91292 101876 91356
rect 113220 91292 113284 91356
rect 115796 91352 115860 91356
rect 115796 91296 115810 91352
rect 115810 91296 115860 91352
rect 115796 91292 115860 91296
rect 118004 91292 118068 91356
rect 124444 91292 124508 91356
rect 125732 91292 125796 91356
rect 151676 91292 151740 91356
rect 74764 91156 74828 91220
rect 85804 91156 85868 91220
rect 86724 91156 86788 91220
rect 88012 91156 88076 91220
rect 90220 91156 90284 91220
rect 91324 91156 91388 91220
rect 93900 91156 93964 91220
rect 97212 91156 97276 91220
rect 98500 91156 98564 91220
rect 99972 91216 100036 91220
rect 99972 91160 100022 91216
rect 100022 91160 100036 91216
rect 99972 91156 100036 91160
rect 100892 91156 100956 91220
rect 101996 91216 102060 91220
rect 101996 91160 102010 91216
rect 102010 91160 102060 91216
rect 101996 91156 102060 91160
rect 102548 91156 102612 91220
rect 102732 91156 102796 91220
rect 104204 91156 104268 91220
rect 105492 91216 105556 91220
rect 105492 91160 105542 91216
rect 105542 91160 105556 91216
rect 105492 91156 105556 91160
rect 105676 91156 105740 91220
rect 106412 91156 106476 91220
rect 108068 91156 108132 91220
rect 109540 91156 109604 91220
rect 112300 91156 112364 91220
rect 114324 91216 114388 91220
rect 114324 91160 114374 91216
rect 114374 91160 114388 91216
rect 114324 91156 114388 91160
rect 115428 91156 115492 91220
rect 118188 91156 118252 91220
rect 119292 91156 119356 91220
rect 120212 91156 120276 91220
rect 120580 91156 120644 91220
rect 122052 91156 122116 91220
rect 125364 91156 125428 91220
rect 126468 91156 126532 91220
rect 127572 91156 127636 91220
rect 129412 91156 129476 91220
rect 132356 91216 132420 91220
rect 132356 91160 132406 91216
rect 132406 91160 132420 91216
rect 132356 91156 132420 91160
rect 151492 91156 151556 91220
rect 152044 91156 152108 91220
rect 107700 90884 107764 90948
rect 95004 90748 95068 90812
rect 197124 90340 197188 90404
rect 219204 86804 219268 86868
rect 267044 86124 267108 86188
rect 166396 81364 166460 81428
rect 166212 78372 166276 78436
rect 168420 68444 168484 68508
rect 224908 68172 224972 68236
rect 66116 66948 66180 67012
rect 264100 59876 264164 59940
rect 267780 58516 267844 58580
rect 266860 54436 266924 54500
rect 242020 53076 242084 53140
rect 267964 50356 268028 50420
rect 220860 43420 220924 43484
rect 240732 40564 240796 40628
rect 255820 29548 255884 29612
rect 260052 28188 260116 28252
rect 227668 22612 227732 22676
rect 186820 14452 186884 14516
rect 169708 11596 169772 11660
rect 195100 11596 195164 11660
rect 166948 8876 167012 8940
rect 173020 8876 173084 8940
rect 177252 4932 177316 4996
rect 253060 3980 253124 4044
rect 246252 3436 246316 3500
rect 249012 3436 249076 3500
rect 285628 3436 285692 3500
rect 287100 3436 287164 3500
rect 288388 3436 288452 3500
rect 291148 3436 291212 3500
rect 298692 3436 298756 3500
rect 191052 3300 191116 3364
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 69611 702540 69677 702541
rect 69611 702476 69612 702540
rect 69676 702476 69677 702540
rect 69611 702475 69677 702476
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 591166 67574 608058
rect 69614 586530 69674 702475
rect 73794 687454 74414 704282
rect 76051 699820 76117 699821
rect 76051 699756 76052 699820
rect 76116 699756 76117 699820
rect 76051 699755 76117 699756
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 591166 74414 614898
rect 69430 586470 69674 586530
rect 67771 583812 67837 583813
rect 67771 583748 67772 583812
rect 67836 583748 67837 583812
rect 67771 583747 67837 583748
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 66667 550900 66733 550901
rect 66667 550836 66668 550900
rect 66732 550836 66733 550900
rect 66667 550835 66733 550836
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 66115 424148 66181 424149
rect 66115 424084 66116 424148
rect 66180 424084 66181 424148
rect 66115 424083 66181 424084
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 66118 359413 66178 424083
rect 66670 411365 66730 550835
rect 66954 536614 67574 537166
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 446407 67574 464058
rect 67774 453933 67834 583747
rect 69430 582317 69490 586470
rect 69427 582316 69493 582317
rect 69427 582252 69428 582316
rect 69492 582252 69493 582316
rect 69427 582251 69493 582252
rect 72679 579454 72999 579486
rect 72679 579218 72721 579454
rect 72957 579218 72999 579454
rect 72679 579134 72999 579218
rect 72679 578898 72721 579134
rect 72957 578898 72999 579134
rect 72679 578866 72999 578898
rect 75644 561454 75964 561486
rect 75644 561218 75686 561454
rect 75922 561218 75964 561454
rect 75644 561134 75964 561218
rect 75644 560898 75686 561134
rect 75922 560898 75964 561134
rect 75644 560866 75964 560898
rect 72679 543454 72999 543486
rect 72679 543218 72721 543454
rect 72957 543218 72999 543454
rect 72679 543134 72999 543218
rect 72679 542898 72721 543134
rect 72957 542898 72999 543134
rect 72679 542866 72999 542898
rect 76054 539613 76114 699755
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 591166 78134 618618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 591166 81854 622338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 591166 85574 626058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 88195 588572 88261 588573
rect 88195 588508 88196 588572
rect 88260 588508 88261 588572
rect 88195 588507 88261 588508
rect 78609 579454 78929 579486
rect 78609 579218 78651 579454
rect 78887 579218 78929 579454
rect 78609 579134 78929 579218
rect 78609 578898 78651 579134
rect 78887 578898 78929 579134
rect 78609 578866 78929 578898
rect 84540 579454 84860 579486
rect 84540 579218 84582 579454
rect 84818 579218 84860 579454
rect 84540 579134 84860 579218
rect 84540 578898 84582 579134
rect 84818 578898 84860 579134
rect 84540 578866 84860 578898
rect 81575 561454 81895 561486
rect 81575 561218 81617 561454
rect 81853 561218 81895 561454
rect 81575 561134 81895 561218
rect 81575 560898 81617 561134
rect 81853 560898 81895 561134
rect 81575 560866 81895 560898
rect 78609 543454 78929 543486
rect 78609 543218 78651 543454
rect 78887 543218 78929 543454
rect 78609 543134 78929 543218
rect 78609 542898 78651 543134
rect 78887 542898 78929 543134
rect 78609 542866 78929 542898
rect 84540 543454 84860 543486
rect 84540 543218 84582 543454
rect 84818 543218 84860 543454
rect 84540 543134 84860 543218
rect 84540 542898 84582 543134
rect 84818 542898 84860 543134
rect 84540 542866 84860 542898
rect 76051 539612 76117 539613
rect 76051 539548 76052 539612
rect 76116 539548 76117 539612
rect 76051 539547 76117 539548
rect 68139 535532 68205 535533
rect 68139 535468 68140 535532
rect 68204 535468 68205 535532
rect 68139 535467 68205 535468
rect 69611 535532 69677 535533
rect 69611 535468 69612 535532
rect 69676 535468 69677 535532
rect 69611 535467 69677 535468
rect 71819 535532 71885 535533
rect 71819 535468 71820 535532
rect 71884 535468 71885 535532
rect 71819 535467 71885 535468
rect 67771 453932 67837 453933
rect 67771 453868 67772 453932
rect 67836 453868 67837 453932
rect 67771 453867 67837 453868
rect 66667 411364 66733 411365
rect 66667 411300 66668 411364
rect 66732 411300 66733 411364
rect 66667 411299 66733 411300
rect 68142 388789 68202 535467
rect 68323 453932 68389 453933
rect 68323 453868 68324 453932
rect 68388 453868 68389 453932
rect 68323 453867 68389 453868
rect 68326 452709 68386 453867
rect 68323 452708 68389 452709
rect 68323 452644 68324 452708
rect 68388 452644 68389 452708
rect 68323 452643 68389 452644
rect 68326 440877 68386 452643
rect 68323 440876 68389 440877
rect 68323 440812 68324 440876
rect 68388 440812 68389 440876
rect 68323 440811 68389 440812
rect 69614 425070 69674 535467
rect 69062 425010 69674 425070
rect 69062 417890 69122 425010
rect 69243 419388 69309 419389
rect 69243 419324 69244 419388
rect 69308 419386 69309 419388
rect 69308 419326 69858 419386
rect 69308 419324 69309 419326
rect 69243 419323 69309 419324
rect 69062 417830 69674 417890
rect 69614 390693 69674 417830
rect 69611 390692 69677 390693
rect 69611 390628 69612 390692
rect 69676 390628 69677 390692
rect 69611 390627 69677 390628
rect 67771 388788 67837 388789
rect 67771 388724 67772 388788
rect 67836 388724 67837 388788
rect 67771 388723 67837 388724
rect 68139 388788 68205 388789
rect 68139 388724 68140 388788
rect 68204 388724 68205 388788
rect 68139 388723 68205 388724
rect 66115 359412 66181 359413
rect 66115 359348 66116 359412
rect 66180 359348 66181 359412
rect 66115 359347 66181 359348
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 61883 330036 61949 330037
rect 61883 329972 61884 330036
rect 61948 329972 61949 330036
rect 61883 329971 61949 329972
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 61886 228445 61946 329971
rect 63234 316894 63854 352338
rect 66954 356614 67574 388356
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66667 349076 66733 349077
rect 66667 349012 66668 349076
rect 66732 349012 66733 349076
rect 66667 349011 66733 349012
rect 66670 347853 66730 349011
rect 66667 347852 66733 347853
rect 66667 347788 66668 347852
rect 66732 347788 66733 347852
rect 66667 347787 66733 347788
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 66670 316437 66730 347787
rect 66954 329592 67574 356058
rect 67774 345677 67834 388723
rect 69798 367709 69858 419326
rect 71822 390421 71882 535467
rect 73794 507454 74414 537166
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 446407 74414 470898
rect 77514 511174 78134 537166
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 446407 78134 474618
rect 81234 514894 81854 537166
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 446407 81854 478338
rect 84954 518614 85574 537166
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446407 85574 482058
rect 88198 460189 88258 588507
rect 91794 561454 92414 596898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 93899 589524 93965 589525
rect 93899 589460 93900 589524
rect 93964 589460 93965 589524
rect 93899 589459 93965 589460
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 89667 462908 89733 462909
rect 89667 462844 89668 462908
rect 89732 462844 89733 462908
rect 89667 462843 89733 462844
rect 88195 460188 88261 460189
rect 88195 460124 88196 460188
rect 88260 460124 88261 460188
rect 88195 460123 88261 460124
rect 72978 435454 73298 435486
rect 72978 435218 73020 435454
rect 73256 435218 73298 435454
rect 72978 435134 73298 435218
rect 72978 434898 73020 435134
rect 73256 434898 73298 435134
rect 72978 434866 73298 434898
rect 88338 417454 88658 417486
rect 88338 417218 88380 417454
rect 88616 417218 88658 417454
rect 88338 417134 88658 417218
rect 88338 416898 88380 417134
rect 88616 416898 88658 417134
rect 88338 416866 88658 416898
rect 72978 399454 73298 399486
rect 72978 399218 73020 399454
rect 73256 399218 73298 399454
rect 72978 399134 73298 399218
rect 72978 398898 73020 399134
rect 73256 398898 73298 399134
rect 72978 398866 73298 398898
rect 71819 390420 71885 390421
rect 71819 390356 71820 390420
rect 71884 390356 71885 390420
rect 71819 390355 71885 390356
rect 89670 389061 89730 462843
rect 91794 453454 92414 488898
rect 92611 454748 92677 454749
rect 92611 454684 92612 454748
rect 92676 454684 92677 454748
rect 92611 454683 92677 454684
rect 91323 453252 91389 453253
rect 91323 453188 91324 453252
rect 91388 453188 91389 453252
rect 91323 453187 91389 453188
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91139 445772 91205 445773
rect 91139 445708 91140 445772
rect 91204 445708 91205 445772
rect 91139 445707 91205 445708
rect 76419 389060 76485 389061
rect 76419 388996 76420 389060
rect 76484 388996 76485 389060
rect 76419 388995 76485 388996
rect 89667 389060 89733 389061
rect 89667 388996 89668 389060
rect 89732 388996 89733 389060
rect 89667 388995 89733 388996
rect 69795 367708 69861 367709
rect 69795 367644 69796 367708
rect 69860 367644 69861 367708
rect 69795 367643 69861 367644
rect 69059 366348 69125 366349
rect 69059 366284 69060 366348
rect 69124 366284 69125 366348
rect 69059 366283 69125 366284
rect 67955 345812 68021 345813
rect 67955 345748 67956 345812
rect 68020 345748 68021 345812
rect 67955 345747 68021 345748
rect 67771 345676 67837 345677
rect 67771 345612 67772 345676
rect 67836 345612 67837 345676
rect 67771 345611 67837 345612
rect 67403 327044 67469 327045
rect 67403 326980 67404 327044
rect 67468 326980 67469 327044
rect 67403 326979 67469 326980
rect 66667 316436 66733 316437
rect 66667 316372 66668 316436
rect 66732 316372 66733 316436
rect 66667 316371 66733 316372
rect 63234 280894 63854 316338
rect 67406 308005 67466 326979
rect 67403 308004 67469 308005
rect 67403 307940 67404 308004
rect 67468 307940 67469 308004
rect 67403 307939 67469 307940
rect 67771 297396 67837 297397
rect 67771 297332 67772 297396
rect 67836 297332 67837 297396
rect 67771 297331 67837 297332
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 65931 276044 65997 276045
rect 65931 275980 65932 276044
rect 65996 275980 65997 276044
rect 65931 275979 65997 275980
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 61883 228444 61949 228445
rect 61883 228380 61884 228444
rect 61948 228380 61949 228444
rect 61883 228379 61949 228380
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 208894 63854 244338
rect 65934 233885 65994 275979
rect 67403 266932 67469 266933
rect 67403 266868 67404 266932
rect 67468 266868 67469 266932
rect 67403 266867 67469 266868
rect 66667 251972 66733 251973
rect 66667 251908 66668 251972
rect 66732 251908 66733 251972
rect 66667 251907 66733 251908
rect 66115 243540 66181 243541
rect 66115 243476 66116 243540
rect 66180 243476 66181 243540
rect 66115 243475 66181 243476
rect 65931 233884 65997 233885
rect 65931 233820 65932 233884
rect 65996 233820 65997 233884
rect 65931 233819 65997 233820
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 66118 67013 66178 243475
rect 66670 206277 66730 251907
rect 67406 242861 67466 266867
rect 67403 242860 67469 242861
rect 67403 242796 67404 242860
rect 67468 242796 67469 242860
rect 67403 242795 67469 242796
rect 66954 212614 67574 239592
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66667 206276 66733 206277
rect 66667 206212 66668 206276
rect 66732 206212 66733 206276
rect 66667 206211 66733 206212
rect 66954 176600 67574 212058
rect 67774 184245 67834 297331
rect 67958 279445 68018 345747
rect 69062 295085 69122 366283
rect 73794 363454 74414 388356
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 70163 360908 70229 360909
rect 70163 360844 70164 360908
rect 70228 360844 70229 360908
rect 70163 360843 70229 360844
rect 70166 349213 70226 360843
rect 69611 349212 69677 349213
rect 69611 349148 69612 349212
rect 69676 349148 69677 349212
rect 69611 349147 69677 349148
rect 70163 349212 70229 349213
rect 70163 349148 70164 349212
rect 70228 349148 70229 349212
rect 70163 349147 70229 349148
rect 69614 316050 69674 349147
rect 73794 329592 74414 362898
rect 69430 315990 69674 316050
rect 69430 315621 69490 315990
rect 69427 315620 69493 315621
rect 69427 315556 69428 315620
rect 69492 315556 69493 315620
rect 69427 315555 69493 315556
rect 69059 295084 69125 295085
rect 69059 295020 69060 295084
rect 69124 295020 69125 295084
rect 69059 295019 69125 295020
rect 72978 291454 73298 291486
rect 72978 291218 73020 291454
rect 73256 291218 73298 291454
rect 72978 291134 73298 291218
rect 72978 290898 73020 291134
rect 73256 290898 73298 291134
rect 72978 290866 73298 290898
rect 67955 279444 68021 279445
rect 67955 279380 67956 279444
rect 68020 279380 68021 279444
rect 67955 279379 68021 279380
rect 69427 256868 69493 256869
rect 69427 256804 69428 256868
rect 69492 256804 69493 256868
rect 69427 256803 69493 256804
rect 67955 256324 68021 256325
rect 67955 256260 67956 256324
rect 68020 256260 68021 256324
rect 67955 256259 68021 256260
rect 67958 229805 68018 256259
rect 69430 248430 69490 256803
rect 72978 255454 73298 255486
rect 72978 255218 73020 255454
rect 73256 255218 73298 255454
rect 72978 255134 73298 255218
rect 72978 254898 73020 255134
rect 73256 254898 73298 255134
rect 72978 254866 73298 254898
rect 69246 248370 69490 248430
rect 69246 243810 69306 248370
rect 69427 245172 69493 245173
rect 69427 245108 69428 245172
rect 69492 245170 69493 245172
rect 69492 245110 69858 245170
rect 69492 245108 69493 245110
rect 69427 245107 69493 245108
rect 69246 243750 69674 243810
rect 69614 232525 69674 243750
rect 69611 232524 69677 232525
rect 69611 232460 69612 232524
rect 69676 232460 69677 232524
rect 69611 232459 69677 232460
rect 69798 230485 69858 245110
rect 69795 230484 69861 230485
rect 69795 230420 69796 230484
rect 69860 230420 69861 230484
rect 69795 230419 69861 230420
rect 67955 229804 68021 229805
rect 67955 229740 67956 229804
rect 68020 229740 68021 229804
rect 67955 229739 68021 229740
rect 73794 219454 74414 239592
rect 76422 231709 76482 388995
rect 77514 367174 78134 388356
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 329592 78134 330618
rect 81234 370894 81854 388356
rect 83411 387292 83477 387293
rect 83411 387228 83412 387292
rect 83476 387228 83477 387292
rect 83411 387227 83477 387228
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 329592 81854 334338
rect 82675 327588 82741 327589
rect 82675 327524 82676 327588
rect 82740 327524 82741 327588
rect 82675 327523 82741 327524
rect 76419 231708 76485 231709
rect 76419 231644 76420 231708
rect 76484 231644 76485 231708
rect 76419 231643 76485 231644
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 67771 184244 67837 184245
rect 67771 184180 67772 184244
rect 67836 184180 67837 184244
rect 67771 184179 67837 184180
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 176600 74414 182898
rect 77514 223174 78134 239592
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 176600 78134 186618
rect 81234 226894 81854 239592
rect 82678 227629 82738 327523
rect 83414 241365 83474 387227
rect 84954 374614 85574 388356
rect 89670 378861 89730 388995
rect 89667 378860 89733 378861
rect 89667 378796 89668 378860
rect 89732 378796 89733 378860
rect 89667 378795 89733 378796
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 91142 359277 91202 445707
rect 91326 390421 91386 453187
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 446407 92414 452898
rect 92614 390965 92674 454683
rect 93902 445773 93962 589459
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 99971 550764 100037 550765
rect 99971 550700 99972 550764
rect 100036 550700 100037 550764
rect 99971 550699 100037 550700
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 98131 458828 98197 458829
rect 98131 458764 98132 458828
rect 98196 458764 98197 458828
rect 98131 458763 98197 458764
rect 96659 457468 96725 457469
rect 96659 457404 96660 457468
rect 96724 457404 96725 457468
rect 96659 457403 96725 457404
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95187 447812 95253 447813
rect 95187 447748 95188 447812
rect 95252 447748 95253 447812
rect 95187 447747 95253 447748
rect 93899 445772 93965 445773
rect 93899 445708 93900 445772
rect 93964 445708 93965 445772
rect 93899 445707 93965 445708
rect 92611 390964 92677 390965
rect 92611 390900 92612 390964
rect 92676 390900 92677 390964
rect 92611 390899 92677 390900
rect 91323 390420 91389 390421
rect 91323 390356 91324 390420
rect 91388 390356 91389 390420
rect 91323 390355 91389 390356
rect 91794 381454 92414 388356
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91139 359276 91205 359277
rect 91139 359212 91140 359276
rect 91204 359212 91205 359276
rect 91139 359211 91205 359212
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 329592 85574 338058
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 329592 92414 344898
rect 93902 332485 93962 445707
rect 95190 390421 95250 447747
rect 95514 446407 96134 456618
rect 96475 445772 96541 445773
rect 96475 445708 96476 445772
rect 96540 445708 96541 445772
rect 96475 445707 96541 445708
rect 95187 390420 95253 390421
rect 95187 390356 95188 390420
rect 95252 390356 95253 390420
rect 95187 390355 95253 390356
rect 96478 388517 96538 445707
rect 96662 390421 96722 457403
rect 97763 445772 97829 445773
rect 97763 445708 97764 445772
rect 97828 445708 97829 445772
rect 97763 445707 97829 445708
rect 96659 390420 96725 390421
rect 96659 390356 96660 390420
rect 96724 390356 96725 390420
rect 96659 390355 96725 390356
rect 96475 388516 96541 388517
rect 96475 388452 96476 388516
rect 96540 388452 96541 388516
rect 96475 388451 96541 388452
rect 95514 385174 96134 388356
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 97766 369885 97826 445707
rect 98134 390421 98194 458763
rect 99234 446407 99854 460338
rect 98131 390420 98197 390421
rect 98131 390356 98132 390420
rect 98196 390356 98197 390420
rect 98131 390355 98197 390356
rect 99974 388381 100034 550699
rect 102954 536614 103574 572058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 111011 553484 111077 553485
rect 111011 553420 111012 553484
rect 111076 553420 111077 553484
rect 111011 553419 111077 553420
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 107699 543012 107765 543013
rect 107699 542948 107700 543012
rect 107764 542948 107765 543012
rect 107699 542947 107765 542948
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 106411 465764 106477 465765
rect 106411 465700 106412 465764
rect 106476 465700 106477 465764
rect 106411 465699 106477 465700
rect 102179 464404 102245 464405
rect 102179 464340 102180 464404
rect 102244 464340 102245 464404
rect 102179 464339 102245 464340
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 100707 456108 100773 456109
rect 100707 456044 100708 456108
rect 100772 456044 100773 456108
rect 100707 456043 100773 456044
rect 100710 390421 100770 456043
rect 102182 390965 102242 464339
rect 102954 464294 103574 464378
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 446407 103574 464058
rect 104939 462908 105005 462909
rect 104939 462844 104940 462908
rect 105004 462844 105005 462908
rect 104939 462843 105005 462844
rect 103698 435454 104018 435486
rect 103698 435218 103740 435454
rect 103976 435218 104018 435454
rect 103698 435134 104018 435218
rect 103698 434898 103740 435134
rect 103976 434898 104018 435134
rect 103698 434866 104018 434898
rect 103698 399454 104018 399486
rect 103698 399218 103740 399454
rect 103976 399218 104018 399454
rect 103698 399134 104018 399218
rect 103698 398898 103740 399134
rect 103976 398898 104018 399134
rect 103698 398866 104018 398898
rect 102179 390964 102245 390965
rect 102179 390900 102180 390964
rect 102244 390900 102245 390964
rect 102179 390899 102245 390900
rect 104942 390421 105002 462843
rect 106414 390421 106474 465699
rect 107702 390421 107762 542947
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 109171 462228 109237 462229
rect 109171 462164 109172 462228
rect 109236 462164 109237 462228
rect 109171 462163 109237 462164
rect 109174 390421 109234 462163
rect 109794 446407 110414 470898
rect 109539 444820 109605 444821
rect 109539 444756 109540 444820
rect 109604 444756 109605 444820
rect 109539 444755 109605 444756
rect 100707 390420 100773 390421
rect 100707 390356 100708 390420
rect 100772 390356 100773 390420
rect 100707 390355 100773 390356
rect 104939 390420 105005 390421
rect 104939 390356 104940 390420
rect 105004 390356 105005 390420
rect 104939 390355 105005 390356
rect 106411 390420 106477 390421
rect 106411 390356 106412 390420
rect 106476 390356 106477 390420
rect 106411 390355 106477 390356
rect 107699 390420 107765 390421
rect 107699 390356 107700 390420
rect 107764 390356 107765 390420
rect 107699 390355 107765 390356
rect 109171 390420 109237 390421
rect 109171 390356 109172 390420
rect 109236 390356 109237 390420
rect 109171 390355 109237 390356
rect 99971 388380 100037 388381
rect 97763 369884 97829 369885
rect 97763 369820 97764 369884
rect 97828 369820 97829 369884
rect 97763 369819 97829 369820
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 93899 332484 93965 332485
rect 93899 332420 93900 332484
rect 93964 332420 93965 332484
rect 93899 332419 93965 332420
rect 95514 329592 96134 348618
rect 99234 352894 99854 388356
rect 99971 388316 99972 388380
rect 100036 388316 100037 388380
rect 99971 388315 100037 388316
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 329592 99854 352338
rect 102954 356614 103574 388356
rect 109542 359005 109602 444755
rect 111014 389197 111074 553419
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 119475 580276 119541 580277
rect 119475 580212 119476 580276
rect 119540 580212 119541 580276
rect 119475 580211 119541 580212
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 115059 538660 115125 538661
rect 115059 538596 115060 538660
rect 115124 538596 115125 538660
rect 115059 538595 115125 538596
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 111747 448628 111813 448629
rect 111747 448564 111748 448628
rect 111812 448564 111813 448628
rect 111747 448563 111813 448564
rect 111563 445772 111629 445773
rect 111563 445708 111564 445772
rect 111628 445708 111629 445772
rect 111563 445707 111629 445708
rect 111011 389196 111077 389197
rect 111011 389132 111012 389196
rect 111076 389132 111077 389196
rect 111011 389131 111077 389132
rect 109794 363454 110414 388356
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109539 359004 109605 359005
rect 109539 358940 109540 359004
rect 109604 358940 109605 359004
rect 109539 358939 109605 358940
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 329592 103574 356058
rect 109794 329592 110414 362898
rect 111566 361861 111626 445707
rect 111750 389061 111810 448563
rect 113514 446407 114134 474618
rect 114323 445772 114389 445773
rect 114323 445708 114324 445772
rect 114388 445708 114389 445772
rect 114323 445707 114389 445708
rect 111747 389060 111813 389061
rect 111747 388996 111748 389060
rect 111812 388996 111813 389060
rect 111747 388995 111813 388996
rect 111563 361860 111629 361861
rect 111563 361796 111564 361860
rect 111628 361796 111629 361860
rect 111563 361795 111629 361796
rect 111750 356693 111810 388995
rect 113514 367174 114134 388356
rect 114326 370021 114386 445707
rect 115062 382261 115122 538595
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 115979 462908 116045 462909
rect 115979 462844 115980 462908
rect 116044 462844 116045 462908
rect 115979 462843 116045 462844
rect 115982 390421 116042 462843
rect 117234 446407 117854 478338
rect 118555 445772 118621 445773
rect 118555 445708 118556 445772
rect 118620 445708 118621 445772
rect 118555 445707 118621 445708
rect 115979 390420 116045 390421
rect 115979 390356 115980 390420
rect 116044 390356 116045 390420
rect 115979 390355 116045 390356
rect 115059 382260 115125 382261
rect 115059 382196 115060 382260
rect 115124 382196 115125 382260
rect 115059 382195 115125 382196
rect 117234 370894 117854 388356
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 114323 370020 114389 370021
rect 114323 369956 114324 370020
rect 114388 369956 114389 370020
rect 114323 369955 114389 369956
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 111747 356692 111813 356693
rect 111747 356628 111748 356692
rect 111812 356628 111813 356692
rect 111747 356627 111813 356628
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 329592 114134 330618
rect 117234 334894 117854 370338
rect 118558 347717 118618 445707
rect 119478 441630 119538 580211
rect 120954 554614 121574 590058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 122971 581636 123037 581637
rect 122971 581572 122972 581636
rect 123036 581572 123037 581636
rect 122971 581571 123037 581572
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120027 447948 120093 447949
rect 120027 447884 120028 447948
rect 120092 447884 120093 447948
rect 120027 447883 120093 447884
rect 120030 441630 120090 447883
rect 120954 446407 121574 482058
rect 122603 447812 122669 447813
rect 122603 447748 122604 447812
rect 122668 447748 122669 447812
rect 122603 447747 122669 447748
rect 119478 441570 119906 441630
rect 120030 441570 120458 441630
rect 119846 431490 119906 441570
rect 120027 431492 120093 431493
rect 120027 431490 120028 431492
rect 119846 431430 120028 431490
rect 120027 431428 120028 431430
rect 120092 431428 120093 431492
rect 120027 431427 120093 431428
rect 119058 417454 119378 417486
rect 119058 417218 119100 417454
rect 119336 417218 119378 417454
rect 119058 417134 119378 417218
rect 119058 416898 119100 417134
rect 119336 416898 119378 417134
rect 119058 416866 119378 416898
rect 120398 412650 120458 441570
rect 122606 431970 122666 447747
rect 122974 435301 123034 581571
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 122971 435300 123037 435301
rect 122971 435236 122972 435300
rect 123036 435236 123037 435300
rect 122971 435235 123037 435236
rect 122422 431910 122666 431970
rect 122422 426325 122482 431910
rect 122603 430948 122669 430949
rect 122603 430884 122604 430948
rect 122668 430884 122669 430948
rect 122603 430883 122669 430884
rect 122419 426324 122485 426325
rect 122419 426260 122420 426324
rect 122484 426260 122485 426324
rect 122419 426259 122485 426260
rect 122422 422381 122482 426259
rect 122419 422380 122485 422381
rect 122419 422316 122420 422380
rect 122484 422316 122485 422380
rect 122419 422315 122485 422316
rect 120030 412590 120458 412650
rect 120030 390421 120090 412590
rect 120027 390420 120093 390421
rect 120027 390356 120028 390420
rect 120092 390356 120093 390420
rect 120027 390355 120093 390356
rect 120954 374614 121574 388356
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 118555 347716 118621 347717
rect 118555 347652 118556 347716
rect 118620 347652 118621 347716
rect 118555 347651 118621 347652
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 329592 117854 334338
rect 120954 338614 121574 374058
rect 122606 361725 122666 430883
rect 122787 422380 122853 422381
rect 122787 422316 122788 422380
rect 122852 422316 122853 422380
rect 122787 422315 122853 422316
rect 122790 422109 122850 422315
rect 122787 422108 122853 422109
rect 122787 422044 122788 422108
rect 122852 422044 122853 422108
rect 122787 422043 122853 422044
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 122787 412860 122853 412861
rect 122787 412796 122788 412860
rect 122852 412796 122853 412860
rect 122787 412795 122853 412796
rect 122790 412453 122850 412795
rect 122787 412452 122853 412453
rect 122787 412388 122788 412452
rect 122852 412388 122853 412452
rect 122787 412387 122853 412388
rect 122787 403068 122853 403069
rect 122787 403004 122788 403068
rect 122852 403004 122853 403068
rect 122787 403003 122853 403004
rect 122790 402930 122850 403003
rect 122971 402932 123037 402933
rect 122971 402930 122972 402932
rect 122790 402870 122972 402930
rect 122971 402868 122972 402870
rect 123036 402868 123037 402932
rect 122971 402867 123037 402868
rect 122971 394772 123037 394773
rect 122971 394708 122972 394772
rect 123036 394708 123037 394772
rect 122971 394707 123037 394708
rect 122787 393412 122853 393413
rect 122787 393348 122788 393412
rect 122852 393348 122853 393412
rect 122787 393347 122853 393348
rect 122790 393277 122850 393347
rect 122787 393276 122853 393277
rect 122787 393212 122788 393276
rect 122852 393212 122853 393276
rect 122787 393211 122853 393212
rect 122974 385661 123034 394707
rect 122971 385660 123037 385661
rect 122971 385596 122972 385660
rect 123036 385596 123037 385660
rect 122971 385595 123037 385596
rect 122787 383892 122853 383893
rect 122787 383828 122788 383892
rect 122852 383828 122853 383892
rect 122787 383827 122853 383828
rect 122790 383621 122850 383827
rect 122787 383620 122853 383621
rect 122787 383556 122788 383620
rect 122852 383556 122853 383620
rect 122787 383555 122853 383556
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 122787 374236 122853 374237
rect 122787 374172 122788 374236
rect 122852 374172 122853 374236
rect 122787 374171 122853 374172
rect 122790 373965 122850 374171
rect 122787 373964 122853 373965
rect 122787 373900 122788 373964
rect 122852 373900 122853 373964
rect 122787 373899 122853 373900
rect 122971 364580 123037 364581
rect 122971 364516 122972 364580
rect 123036 364516 123037 364580
rect 122971 364515 123037 364516
rect 122974 364173 123034 364515
rect 122971 364172 123037 364173
rect 122971 364108 122972 364172
rect 123036 364108 123037 364172
rect 122971 364107 123037 364108
rect 122603 361724 122669 361725
rect 122603 361660 122604 361724
rect 122668 361660 122669 361724
rect 122603 361659 122669 361660
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 329592 121574 338058
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 329592 128414 344898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 133091 442372 133157 442373
rect 133091 442308 133092 442372
rect 133156 442308 133157 442372
rect 133091 442307 133157 442308
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 329592 132134 348618
rect 88338 309454 88658 309486
rect 88338 309218 88380 309454
rect 88616 309218 88658 309454
rect 88338 309134 88658 309218
rect 88338 308898 88380 309134
rect 88616 308898 88658 309134
rect 88338 308866 88658 308898
rect 119058 309454 119378 309486
rect 119058 309218 119100 309454
rect 119336 309218 119378 309454
rect 119058 309134 119378 309218
rect 119058 308898 119100 309134
rect 119336 308898 119378 309134
rect 119058 308866 119378 308898
rect 103698 291454 104018 291486
rect 103698 291218 103740 291454
rect 103976 291218 104018 291454
rect 103698 291134 104018 291218
rect 103698 290898 103740 291134
rect 103976 290898 104018 291134
rect 103698 290866 104018 290898
rect 88338 273454 88658 273486
rect 88338 273218 88380 273454
rect 88616 273218 88658 273454
rect 88338 273134 88658 273218
rect 88338 272898 88380 273134
rect 88616 272898 88658 273134
rect 88338 272866 88658 272898
rect 119058 273454 119378 273486
rect 119058 273218 119100 273454
rect 119336 273218 119378 273454
rect 119058 273134 119378 273218
rect 119058 272898 119100 273134
rect 119336 272898 119378 273134
rect 119058 272866 119378 272898
rect 103698 255454 104018 255486
rect 103698 255218 103740 255454
rect 103976 255218 104018 255454
rect 103698 255134 104018 255218
rect 103698 254898 103740 255134
rect 103976 254898 104018 255134
rect 103698 254866 104018 254898
rect 83411 241364 83477 241365
rect 83411 241300 83412 241364
rect 83476 241300 83477 241364
rect 83411 241299 83477 241300
rect 84954 230614 85574 239592
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 82675 227628 82741 227629
rect 82675 227564 82676 227628
rect 82740 227564 82741 227628
rect 82675 227563 82741 227564
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 176600 81854 190338
rect 84954 194614 85574 230058
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 176600 85574 194058
rect 91794 237454 92414 239592
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 95514 205174 96134 239592
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 176600 96134 204618
rect 99234 208894 99854 239592
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 97027 177988 97093 177989
rect 97027 177924 97028 177988
rect 97092 177924 97093 177988
rect 97027 177923 97093 177924
rect 97030 175130 97090 177923
rect 98315 177580 98381 177581
rect 98315 177516 98316 177580
rect 98380 177516 98381 177580
rect 98315 177515 98381 177516
rect 96960 175070 97090 175130
rect 98318 175130 98378 177515
rect 99234 176600 99854 208338
rect 102954 212614 103574 239592
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 101995 177580 102061 177581
rect 101995 177516 101996 177580
rect 102060 177516 102061 177580
rect 101995 177515 102061 177516
rect 100707 176900 100773 176901
rect 100707 176836 100708 176900
rect 100772 176836 100773 176900
rect 100707 176835 100773 176836
rect 99419 176492 99485 176493
rect 99419 176428 99420 176492
rect 99484 176428 99485 176492
rect 99419 176427 99485 176428
rect 99422 175130 99482 176427
rect 98318 175070 98380 175130
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 176835
rect 101998 175130 102058 177515
rect 102954 176600 103574 212058
rect 109794 219454 110414 239592
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 109539 178396 109605 178397
rect 109539 178332 109540 178396
rect 109604 178332 109605 178396
rect 109539 178331 109605 178332
rect 105675 177580 105741 177581
rect 105675 177516 105676 177580
rect 105740 177516 105741 177580
rect 105675 177515 105741 177516
rect 108067 177580 108133 177581
rect 108067 177516 108068 177580
rect 108132 177516 108133 177580
rect 108067 177515 108133 177516
rect 104571 177172 104637 177173
rect 104571 177108 104572 177172
rect 104636 177108 104637 177172
rect 104571 177107 104637 177108
rect 103283 176492 103349 176493
rect 103283 176428 103284 176492
rect 103348 176428 103349 176492
rect 103283 176427 103349 176428
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 176427
rect 104574 175130 104634 177107
rect 105678 175130 105738 177515
rect 106963 176764 107029 176765
rect 106963 176700 106964 176764
rect 107028 176700 107029 176764
rect 106963 176699 107029 176700
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 105738 175130
rect 106966 175130 107026 176699
rect 108070 175130 108130 177515
rect 109542 175130 109602 178331
rect 109794 176600 110414 182898
rect 113514 223174 114134 239592
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 110643 178260 110709 178261
rect 110643 178196 110644 178260
rect 110708 178196 110709 178260
rect 110643 178195 110709 178196
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109472 175070 109602 175130
rect 110646 175130 110706 178195
rect 112115 177580 112181 177581
rect 112115 177516 112116 177580
rect 112180 177516 112181 177580
rect 112115 177515 112181 177516
rect 112118 175130 112178 177515
rect 113219 177036 113285 177037
rect 113219 176972 113220 177036
rect 113284 176972 113285 177036
rect 113219 176971 113285 176972
rect 113222 175130 113282 176971
rect 113514 176600 114134 186618
rect 117234 226894 117854 239592
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 115795 177036 115861 177037
rect 115795 176972 115796 177036
rect 115860 176972 115861 177036
rect 115795 176971 115861 176972
rect 114323 175540 114389 175541
rect 114323 175476 114324 175540
rect 114388 175476 114389 175540
rect 114323 175475 114389 175476
rect 110646 175070 110756 175130
rect 109472 174494 109532 175070
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 113144 175070 113282 175130
rect 114326 175130 114386 175475
rect 115798 175130 115858 176971
rect 117234 176600 117854 190338
rect 120954 230614 121574 239592
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 120763 177580 120829 177581
rect 120763 177516 120764 177580
rect 120828 177516 120829 177580
rect 120763 177515 120829 177516
rect 118371 177444 118437 177445
rect 118371 177380 118372 177444
rect 118436 177380 118437 177444
rect 118371 177379 118437 177380
rect 116899 175404 116965 175405
rect 116899 175340 116900 175404
rect 116964 175340 116965 175404
rect 116899 175339 116965 175340
rect 114326 175070 114428 175130
rect 112056 174494 112116 175070
rect 113144 174494 113204 175070
rect 114368 174494 114428 175070
rect 115728 175070 115858 175130
rect 116902 175130 116962 175339
rect 118374 175130 118434 177379
rect 120766 175130 120826 177515
rect 120954 176600 121574 194058
rect 127794 237454 128414 239592
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 124443 177580 124509 177581
rect 124443 177516 124444 177580
rect 124508 177516 124509 177580
rect 124443 177515 124509 177516
rect 125731 177580 125797 177581
rect 125731 177516 125732 177580
rect 125796 177516 125797 177580
rect 125731 177515 125797 177516
rect 127019 177580 127085 177581
rect 127019 177516 127020 177580
rect 127084 177516 127085 177580
rect 127019 177515 127085 177516
rect 121867 176764 121933 176765
rect 121867 176700 121868 176764
rect 121932 176700 121933 176764
rect 121867 176699 121933 176700
rect 123155 176764 123221 176765
rect 123155 176700 123156 176764
rect 123220 176700 123221 176764
rect 123155 176699 123221 176700
rect 121870 175130 121930 176699
rect 123158 175130 123218 176699
rect 124446 175130 124506 177515
rect 125734 175130 125794 177515
rect 127022 175130 127082 177515
rect 127794 176600 128414 200898
rect 131514 205174 132134 239592
rect 133094 231437 133154 442307
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 136587 378724 136653 378725
rect 136587 378660 136588 378724
rect 136652 378660 136653 378724
rect 136587 378659 136653 378660
rect 136035 358052 136101 358053
rect 136035 357988 136036 358052
rect 136100 357988 136101 358052
rect 136035 357987 136101 357988
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 329592 135854 352338
rect 134418 291454 134738 291486
rect 134418 291218 134460 291454
rect 134696 291218 134738 291454
rect 134418 291134 134738 291218
rect 134418 290898 134460 291134
rect 134696 290898 134738 291134
rect 134418 290866 134738 290898
rect 134418 255454 134738 255486
rect 134418 255218 134460 255454
rect 134696 255218 134738 255454
rect 134418 255134 134738 255218
rect 134418 254898 134460 255134
rect 134696 254898 134738 255134
rect 134418 254866 134738 254898
rect 136038 242045 136098 357987
rect 136590 242045 136650 378659
rect 138059 362268 138125 362269
rect 138059 362204 138060 362268
rect 138124 362204 138125 362268
rect 138059 362203 138125 362204
rect 138062 242045 138122 362203
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 329592 139574 356058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 146891 435300 146957 435301
rect 146891 435236 146892 435300
rect 146956 435236 146957 435300
rect 146891 435235 146957 435236
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 146894 365941 146954 435235
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 146891 365940 146957 365941
rect 146891 365876 146892 365940
rect 146956 365876 146957 365940
rect 146891 365875 146957 365876
rect 146894 364350 146954 365875
rect 146894 364290 147506 364350
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 139715 352612 139781 352613
rect 139715 352548 139716 352612
rect 139780 352548 139781 352612
rect 139715 352547 139781 352548
rect 136035 242044 136101 242045
rect 136035 241980 136036 242044
rect 136100 241980 136101 242044
rect 136035 241979 136101 241980
rect 136587 242044 136653 242045
rect 136587 241980 136588 242044
rect 136652 241980 136653 242044
rect 136587 241979 136653 241980
rect 138059 242044 138125 242045
rect 138059 241980 138060 242044
rect 138124 241980 138125 242044
rect 138059 241979 138125 241980
rect 133091 231436 133157 231437
rect 133091 231372 133092 231436
rect 133156 231372 133157 231436
rect 133091 231371 133157 231372
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 130699 177308 130765 177309
rect 130699 177244 130700 177308
rect 130764 177244 130765 177308
rect 130699 177243 130765 177244
rect 129411 176764 129477 176765
rect 129411 176700 129412 176764
rect 129476 176700 129477 176764
rect 129411 176699 129477 176700
rect 128123 176492 128189 176493
rect 128123 176428 128124 176492
rect 128188 176428 128189 176492
rect 128123 176427 128189 176428
rect 128126 175130 128186 176427
rect 116902 175070 117012 175130
rect 115728 174494 115788 175070
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 123072 175070 123218 175130
rect 124432 175070 124506 175130
rect 125656 175070 125794 175130
rect 127016 175070 127082 175130
rect 128104 175070 128186 175130
rect 129414 175130 129474 176699
rect 130702 175130 130762 177243
rect 131514 176600 132134 204618
rect 135234 208894 135854 239592
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 132355 177580 132421 177581
rect 132355 177516 132356 177580
rect 132420 177516 132421 177580
rect 132355 177515 132421 177516
rect 133091 177580 133157 177581
rect 133091 177516 133092 177580
rect 133156 177516 133157 177580
rect 133091 177515 133157 177516
rect 132358 175130 132418 177515
rect 129414 175070 129524 175130
rect 118312 174494 118372 175070
rect 119397 174996 119463 174997
rect 119397 174932 119398 174996
rect 119462 174932 119463 174996
rect 119397 174931 119463 174932
rect 119400 174494 119460 174931
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123072 174494 123132 175070
rect 124432 174494 124492 175070
rect 125656 174494 125716 175070
rect 127016 174494 127076 175070
rect 128104 174494 128164 175070
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 132048 175070 132418 175130
rect 133094 175130 133154 177515
rect 135234 176600 135854 208338
rect 138954 212614 139574 239592
rect 139718 233069 139778 352547
rect 145794 329592 146414 362898
rect 145603 327180 145669 327181
rect 145603 327116 145604 327180
rect 145668 327116 145669 327180
rect 145603 327115 145669 327116
rect 139715 233068 139781 233069
rect 139715 233004 139716 233068
rect 139780 233004 139781 233068
rect 139715 233003 139781 233004
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 136035 176764 136101 176765
rect 136035 176700 136036 176764
rect 136100 176700 136101 176764
rect 136035 176699 136101 176700
rect 136038 175130 136098 176699
rect 138954 176600 139574 212058
rect 145606 185741 145666 327115
rect 147446 242045 147506 364290
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 329592 150134 330618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 158667 451348 158733 451349
rect 158667 451284 158668 451348
rect 158732 451284 158733 451348
rect 158667 451283 158733 451284
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 155171 446044 155237 446045
rect 155171 445980 155172 446044
rect 155236 445980 155237 446044
rect 155171 445979 155237 445980
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 329592 153854 334338
rect 154251 330036 154317 330037
rect 154251 329972 154252 330036
rect 154316 329972 154317 330036
rect 154251 329971 154317 329972
rect 153699 327724 153765 327725
rect 153699 327660 153700 327724
rect 153764 327660 153765 327724
rect 153699 327659 153765 327660
rect 150387 327180 150453 327181
rect 150387 327116 150388 327180
rect 150452 327116 150453 327180
rect 150387 327115 150453 327116
rect 149778 309454 150098 309486
rect 149778 309218 149820 309454
rect 150056 309218 150098 309454
rect 149778 309134 150098 309218
rect 149778 308898 149820 309134
rect 150056 308898 150098 309134
rect 149778 308866 150098 308898
rect 149778 273454 150098 273486
rect 149778 273218 149820 273454
rect 150056 273218 150098 273454
rect 149778 273134 150098 273218
rect 149778 272898 149820 273134
rect 150056 272898 150098 273134
rect 149778 272866 150098 272898
rect 147443 242044 147509 242045
rect 147443 241980 147444 242044
rect 147508 241980 147509 242044
rect 147443 241979 147509 241980
rect 145794 219454 146414 239592
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145603 185740 145669 185741
rect 145603 185676 145604 185740
rect 145668 185676 145669 185740
rect 145603 185675 145669 185676
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 149514 223174 150134 239592
rect 150390 224229 150450 327115
rect 153702 316050 153762 327659
rect 154254 320789 154314 329971
rect 154251 320788 154317 320789
rect 154251 320724 154252 320788
rect 154316 320724 154317 320788
rect 154251 320723 154317 320724
rect 155174 318613 155234 445979
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156459 347172 156525 347173
rect 156459 347108 156460 347172
rect 156524 347108 156525 347172
rect 156459 347107 156525 347108
rect 155355 327180 155421 327181
rect 155355 327116 155356 327180
rect 155420 327116 155421 327180
rect 155355 327115 155421 327116
rect 155171 318612 155237 318613
rect 155171 318548 155172 318612
rect 155236 318548 155237 318612
rect 155171 318547 155237 318548
rect 155358 318205 155418 327115
rect 155355 318204 155421 318205
rect 155355 318140 155356 318204
rect 155420 318140 155421 318204
rect 155355 318139 155421 318140
rect 153702 315990 154314 316050
rect 154254 315077 154314 315990
rect 154251 315076 154317 315077
rect 154251 315012 154252 315076
rect 154316 315012 154317 315076
rect 154251 315011 154317 315012
rect 156462 291141 156522 347107
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156459 291140 156525 291141
rect 156459 291076 156460 291140
rect 156524 291076 156525 291140
rect 156459 291075 156525 291076
rect 155171 275364 155237 275365
rect 155171 275300 155172 275364
rect 155236 275300 155237 275364
rect 155171 275299 155237 275300
rect 154619 260812 154685 260813
rect 154619 260748 154620 260812
rect 154684 260748 154685 260812
rect 154619 260747 154685 260748
rect 154435 244492 154501 244493
rect 154435 244428 154436 244492
rect 154500 244428 154501 244492
rect 154435 244427 154501 244428
rect 154438 240005 154498 244427
rect 154435 240004 154501 240005
rect 154435 239940 154436 240004
rect 154500 239940 154501 240004
rect 154435 239939 154501 239940
rect 153234 226894 153854 239592
rect 154622 229110 154682 260747
rect 155174 237285 155234 275299
rect 156954 266614 157574 302058
rect 158670 295357 158730 451283
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163451 377364 163517 377365
rect 163451 377300 163452 377364
rect 163516 377300 163517 377364
rect 163451 377299 163517 377300
rect 160691 331532 160757 331533
rect 160691 331468 160692 331532
rect 160756 331468 160757 331532
rect 160691 331467 160757 331468
rect 160694 313989 160754 331467
rect 160875 326500 160941 326501
rect 160875 326436 160876 326500
rect 160940 326436 160941 326500
rect 160875 326435 160941 326436
rect 160691 313988 160757 313989
rect 160691 313924 160692 313988
rect 160756 313924 160757 313988
rect 160691 313923 160757 313924
rect 160878 311133 160938 326435
rect 160875 311132 160941 311133
rect 160875 311068 160876 311132
rect 160940 311068 160941 311132
rect 160875 311067 160941 311068
rect 158667 295356 158733 295357
rect 158667 295292 158668 295356
rect 158732 295292 158733 295356
rect 158667 295291 158733 295292
rect 163454 280125 163514 377299
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163451 280124 163517 280125
rect 163451 280060 163452 280124
rect 163516 280060 163517 280124
rect 163451 280059 163517 280060
rect 163794 273454 164414 308898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 169707 369068 169773 369069
rect 169707 369004 169708 369068
rect 169772 369004 169773 369068
rect 169707 369003 169773 369004
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 166211 292636 166277 292637
rect 166211 292572 166212 292636
rect 166276 292572 166277 292636
rect 166211 292571 166277 292572
rect 160691 273324 160757 273325
rect 160691 273260 160692 273324
rect 160756 273260 160757 273324
rect 160691 273259 160757 273260
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 155171 237284 155237 237285
rect 155171 237220 155172 237284
rect 155236 237220 155237 237284
rect 155171 237219 155237 237220
rect 156954 230614 157574 266058
rect 160694 246261 160754 273259
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 161979 269380 162045 269381
rect 161979 269316 161980 269380
rect 162044 269316 162045 269380
rect 161979 269315 162045 269316
rect 160691 246260 160757 246261
rect 160691 246196 160692 246260
rect 160756 246196 160757 246260
rect 160691 246195 160757 246196
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 154622 229050 155234 229110
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 150387 224228 150453 224229
rect 150387 224164 150388 224228
rect 150452 224164 150453 224228
rect 150387 224163 150453 224164
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 148179 177580 148245 177581
rect 148179 177516 148180 177580
rect 148244 177516 148245 177580
rect 148179 177515 148245 177516
rect 133094 175070 133196 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 135720 175070 136098 175130
rect 148182 175130 148242 177515
rect 149514 176600 150134 186618
rect 153234 190894 153854 226338
rect 155174 219197 155234 229050
rect 155171 219196 155237 219197
rect 155171 219132 155172 219196
rect 155236 219132 155237 219196
rect 155171 219131 155237 219132
rect 155174 210357 155234 219131
rect 155171 210356 155237 210357
rect 155171 210292 155172 210356
rect 155236 210292 155237 210356
rect 155171 210291 155237 210292
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 176600 153854 190338
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 176600 157574 194058
rect 161982 189821 162042 269315
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 166214 210357 166274 292571
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 168419 251428 168485 251429
rect 168419 251364 168420 251428
rect 168484 251364 168485 251428
rect 168419 251363 168485 251364
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 166211 210356 166277 210357
rect 166211 210292 166212 210356
rect 166276 210292 166277 210356
rect 166211 210291 166277 210292
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 161979 189820 162045 189821
rect 161979 189756 161980 189820
rect 162044 189756 162045 189820
rect 161979 189755 162045 189756
rect 158851 176764 158917 176765
rect 158851 176700 158852 176764
rect 158916 176700 158917 176764
rect 158851 176699 158917 176700
rect 158854 175130 158914 176699
rect 163794 176600 164414 200898
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 166947 175948 167013 175949
rect 166947 175884 166948 175948
rect 167012 175884 167013 175948
rect 166947 175883 167013 175884
rect 148182 175070 148292 175130
rect 134357 174860 134423 174861
rect 134357 174796 134358 174860
rect 134422 174796 134423 174860
rect 134357 174795 134423 174796
rect 134360 174494 134420 174795
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 69072 165454 69420 165486
rect 69072 165218 69128 165454
rect 69364 165218 69420 165454
rect 69072 165134 69420 165218
rect 69072 164898 69128 165134
rect 69364 164898 69420 165134
rect 69072 164866 69420 164898
rect 164136 165454 164484 165486
rect 164136 165218 164192 165454
rect 164428 165218 164484 165454
rect 164136 165134 164484 165218
rect 164136 164898 164192 165134
rect 164428 164898 164484 165134
rect 164136 164866 164484 164898
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 69072 129454 69420 129486
rect 69072 129218 69128 129454
rect 69364 129218 69420 129454
rect 69072 129134 69420 129218
rect 69072 128898 69128 129134
rect 69364 128898 69420 129134
rect 69072 128866 69420 128898
rect 164136 129454 164484 129486
rect 164136 129218 164192 129454
rect 164428 129218 164484 129454
rect 164136 129134 164484 129218
rect 164136 128898 164192 129134
rect 164428 128898 164484 129134
rect 164136 128866 164484 128898
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 166211 102508 166277 102509
rect 166211 102444 166212 102508
rect 166276 102444 166277 102508
rect 166211 102443 166277 102444
rect 74656 94890 74716 95200
rect 84312 94890 84372 95200
rect 85536 94890 85596 95200
rect 86624 94890 86684 95200
rect 87984 94890 88044 95200
rect 88936 94890 88996 95200
rect 74656 94830 74826 94890
rect 84312 94830 84394 94890
rect 85536 94830 85866 94890
rect 86624 94830 86786 94890
rect 87984 94830 88074 94890
rect 66954 68614 67574 93100
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66115 67012 66181 67013
rect 66115 66948 66116 67012
rect 66180 66948 66181 67012
rect 66115 66947 66181 66948
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 75454 74414 93100
rect 74766 91221 74826 94830
rect 74763 91220 74829 91221
rect 74763 91156 74764 91220
rect 74828 91156 74829 91220
rect 74763 91155 74829 91156
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 93100
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 93100
rect 84334 92445 84394 94830
rect 84331 92444 84397 92445
rect 84331 92380 84332 92444
rect 84396 92380 84397 92444
rect 84331 92379 84397 92380
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 93100
rect 85806 91221 85866 94830
rect 86726 91221 86786 94830
rect 88014 91221 88074 94830
rect 88934 94830 88996 94890
rect 90160 94890 90220 95200
rect 91384 94890 91444 95200
rect 90160 94830 90282 94890
rect 88934 92445 88994 94830
rect 88931 92444 88997 92445
rect 88931 92380 88932 92444
rect 88996 92380 88997 92444
rect 88931 92379 88997 92380
rect 90222 91221 90282 94830
rect 91326 94830 91444 94890
rect 92472 94890 92532 95200
rect 93832 94890 93892 95200
rect 94920 94890 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 92472 94830 92674 94890
rect 93832 94830 93962 94890
rect 94920 94830 95066 94890
rect 96008 94830 96354 94890
rect 91326 91221 91386 94830
rect 85803 91220 85869 91221
rect 85803 91156 85804 91220
rect 85868 91156 85869 91220
rect 85803 91155 85869 91156
rect 86723 91220 86789 91221
rect 86723 91156 86724 91220
rect 86788 91156 86789 91220
rect 86723 91155 86789 91156
rect 88011 91220 88077 91221
rect 88011 91156 88012 91220
rect 88076 91156 88077 91220
rect 88011 91155 88077 91156
rect 90219 91220 90285 91221
rect 90219 91156 90220 91220
rect 90284 91156 90285 91220
rect 90219 91155 90285 91156
rect 91323 91220 91389 91221
rect 91323 91156 91324 91220
rect 91388 91156 91389 91220
rect 91323 91155 91389 91156
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 93100
rect 92614 91765 92674 94830
rect 92611 91764 92677 91765
rect 92611 91700 92612 91764
rect 92676 91700 92677 91764
rect 92611 91699 92677 91700
rect 93902 91221 93962 94830
rect 93899 91220 93965 91221
rect 93899 91156 93900 91220
rect 93964 91156 93965 91220
rect 93899 91155 93965 91156
rect 95006 90813 95066 94830
rect 95003 90812 95069 90813
rect 95003 90748 95004 90812
rect 95068 90748 95069 90812
rect 95003 90747 95069 90748
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 93100
rect 96294 91901 96354 94830
rect 96662 94830 96748 94890
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 96291 91900 96357 91901
rect 96291 91836 96292 91900
rect 96356 91836 96357 91900
rect 96291 91835 96357 91836
rect 96662 91357 96722 94830
rect 96659 91356 96725 91357
rect 96659 91292 96660 91356
rect 96724 91292 96725 91356
rect 96659 91291 96725 91292
rect 97214 91221 97274 94830
rect 98134 91765 98194 94830
rect 98131 91764 98197 91765
rect 98131 91700 98132 91764
rect 98196 91700 98197 91764
rect 98131 91699 98197 91700
rect 98502 91221 98562 94830
rect 99054 94830 99196 94890
rect 99544 94890 99604 95200
rect 99544 94830 100034 94890
rect 99054 92445 99114 94830
rect 99051 92444 99117 92445
rect 99051 92380 99052 92444
rect 99116 92380 99117 92444
rect 99051 92379 99117 92380
rect 97211 91220 97277 91221
rect 97211 91156 97212 91220
rect 97276 91156 97277 91220
rect 97211 91155 97277 91156
rect 98499 91220 98565 91221
rect 98499 91156 98500 91220
rect 98564 91156 98565 91220
rect 98499 91155 98565 91156
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 93100
rect 99974 91221 100034 94830
rect 100632 94757 100692 95200
rect 100768 94890 100828 95200
rect 101856 94890 101916 95200
rect 100768 94830 100954 94890
rect 100629 94756 100695 94757
rect 100629 94692 100630 94756
rect 100694 94692 100695 94756
rect 100629 94691 100695 94692
rect 100894 91221 100954 94830
rect 101814 94830 101916 94890
rect 101992 94890 102052 95200
rect 102944 94890 103004 95200
rect 103216 94890 103276 95200
rect 104304 94890 104364 95200
rect 101992 94830 102058 94890
rect 101814 91357 101874 94830
rect 101811 91356 101877 91357
rect 101811 91292 101812 91356
rect 101876 91292 101877 91356
rect 101811 91291 101877 91292
rect 101998 91221 102058 94830
rect 102550 94830 103004 94890
rect 103102 94830 103276 94890
rect 104206 94830 104364 94890
rect 104440 94890 104500 95200
rect 105392 94890 105452 95200
rect 105664 94890 105724 95200
rect 106480 94890 106540 95200
rect 104440 94830 104634 94890
rect 105392 94830 105554 94890
rect 105664 94830 105738 94890
rect 102550 91221 102610 94830
rect 103102 93870 103162 94830
rect 102734 93810 103162 93870
rect 102734 91221 102794 93810
rect 99971 91220 100037 91221
rect 99971 91156 99972 91220
rect 100036 91156 100037 91220
rect 99971 91155 100037 91156
rect 100891 91220 100957 91221
rect 100891 91156 100892 91220
rect 100956 91156 100957 91220
rect 100891 91155 100957 91156
rect 101995 91220 102061 91221
rect 101995 91156 101996 91220
rect 102060 91156 102061 91220
rect 101995 91155 102061 91156
rect 102547 91220 102613 91221
rect 102547 91156 102548 91220
rect 102612 91156 102613 91220
rect 102547 91155 102613 91156
rect 102731 91220 102797 91221
rect 102731 91156 102732 91220
rect 102796 91156 102797 91220
rect 102731 91155 102797 91156
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 93100
rect 104206 91221 104266 94830
rect 104574 91629 104634 94830
rect 104571 91628 104637 91629
rect 104571 91564 104572 91628
rect 104636 91564 104637 91628
rect 104571 91563 104637 91564
rect 105494 91221 105554 94830
rect 105678 91221 105738 94830
rect 106414 94830 106540 94890
rect 106616 94890 106676 95200
rect 107704 94890 107764 95200
rect 108112 94890 108172 95200
rect 106616 94830 106842 94890
rect 106414 91221 106474 94830
rect 106782 92445 106842 94830
rect 107702 94830 107764 94890
rect 108070 94830 108172 94890
rect 109064 94890 109124 95200
rect 109472 94890 109532 95200
rect 110152 94890 110212 95200
rect 110696 94890 110756 95200
rect 111240 94890 111300 95200
rect 109064 94830 109234 94890
rect 109472 94830 109602 94890
rect 106779 92444 106845 92445
rect 106779 92380 106780 92444
rect 106844 92380 106845 92444
rect 106779 92379 106845 92380
rect 104203 91220 104269 91221
rect 104203 91156 104204 91220
rect 104268 91156 104269 91220
rect 104203 91155 104269 91156
rect 105491 91220 105557 91221
rect 105491 91156 105492 91220
rect 105556 91156 105557 91220
rect 105491 91155 105557 91156
rect 105675 91220 105741 91221
rect 105675 91156 105676 91220
rect 105740 91156 105741 91220
rect 105675 91155 105741 91156
rect 106411 91220 106477 91221
rect 106411 91156 106412 91220
rect 106476 91156 106477 91220
rect 106411 91155 106477 91156
rect 107702 90949 107762 94830
rect 108070 91221 108130 94830
rect 109174 92445 109234 94830
rect 109171 92444 109237 92445
rect 109171 92380 109172 92444
rect 109236 92380 109237 92444
rect 109171 92379 109237 92380
rect 109542 91221 109602 94830
rect 110094 94830 110212 94890
rect 110646 94830 110756 94890
rect 111198 94830 111300 94890
rect 111920 94890 111980 95200
rect 112328 94890 112388 95200
rect 111920 94830 111994 94890
rect 110094 93261 110154 94830
rect 110091 93260 110157 93261
rect 110091 93196 110092 93260
rect 110156 93196 110157 93260
rect 110091 93195 110157 93196
rect 108067 91220 108133 91221
rect 108067 91156 108068 91220
rect 108132 91156 108133 91220
rect 108067 91155 108133 91156
rect 109539 91220 109605 91221
rect 109539 91156 109540 91220
rect 109604 91156 109605 91220
rect 109539 91155 109605 91156
rect 107699 90948 107765 90949
rect 107699 90884 107700 90948
rect 107764 90884 107765 90948
rect 107699 90883 107765 90884
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 75454 110414 93100
rect 110646 92445 110706 94830
rect 111198 92445 111258 94830
rect 111934 93941 111994 94830
rect 112302 94830 112388 94890
rect 113144 94890 113204 95200
rect 113688 94890 113748 95200
rect 114368 94890 114428 95200
rect 113144 94830 113282 94890
rect 113688 94830 113834 94890
rect 111931 93940 111997 93941
rect 111931 93876 111932 93940
rect 111996 93876 111997 93940
rect 111931 93875 111997 93876
rect 110643 92444 110709 92445
rect 110643 92380 110644 92444
rect 110708 92380 110709 92444
rect 110643 92379 110709 92380
rect 111195 92444 111261 92445
rect 111195 92380 111196 92444
rect 111260 92380 111261 92444
rect 111195 92379 111261 92380
rect 112302 91221 112362 94830
rect 113222 91357 113282 94830
rect 113774 93261 113834 94830
rect 114326 94830 114428 94890
rect 114776 94890 114836 95200
rect 115456 94890 115516 95200
rect 115864 94890 115924 95200
rect 114776 94830 114938 94890
rect 113771 93260 113837 93261
rect 113771 93196 113772 93260
rect 113836 93196 113837 93260
rect 113771 93195 113837 93196
rect 113219 91356 113285 91357
rect 113219 91292 113220 91356
rect 113284 91292 113285 91356
rect 113219 91291 113285 91292
rect 112299 91220 112365 91221
rect 112299 91156 112300 91220
rect 112364 91156 112365 91220
rect 112299 91155 112365 91156
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 79174 114134 93100
rect 114326 91221 114386 94830
rect 114878 93805 114938 94830
rect 115430 94830 115516 94890
rect 115798 94830 115924 94890
rect 116680 94890 116740 95200
rect 117088 94890 117148 95200
rect 116680 94830 116778 94890
rect 114875 93804 114941 93805
rect 114875 93740 114876 93804
rect 114940 93740 114941 93804
rect 114875 93739 114941 93740
rect 115430 91221 115490 94830
rect 115798 91357 115858 94830
rect 116718 92309 116778 94830
rect 117086 94830 117148 94890
rect 117904 94890 117964 95200
rect 118176 94890 118236 95200
rect 119400 94890 119460 95200
rect 117904 94830 118066 94890
rect 118176 94830 118250 94890
rect 117086 93533 117146 94830
rect 117083 93532 117149 93533
rect 117083 93468 117084 93532
rect 117148 93468 117149 93532
rect 117083 93467 117149 93468
rect 116715 92308 116781 92309
rect 116715 92244 116716 92308
rect 116780 92244 116781 92308
rect 116715 92243 116781 92244
rect 115795 91356 115861 91357
rect 115795 91292 115796 91356
rect 115860 91292 115861 91356
rect 115795 91291 115861 91292
rect 114323 91220 114389 91221
rect 114323 91156 114324 91220
rect 114388 91156 114389 91220
rect 114323 91155 114389 91156
rect 115427 91220 115493 91221
rect 115427 91156 115428 91220
rect 115492 91156 115493 91220
rect 115427 91155 115493 91156
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 82894 117854 93100
rect 118006 91357 118066 94830
rect 118003 91356 118069 91357
rect 118003 91292 118004 91356
rect 118068 91292 118069 91356
rect 118003 91291 118069 91292
rect 118190 91221 118250 94830
rect 119294 94830 119460 94890
rect 119536 94890 119596 95200
rect 120216 94890 120276 95200
rect 120624 94890 120684 95200
rect 121712 94890 121772 95200
rect 119536 94830 119722 94890
rect 119294 91221 119354 94830
rect 119662 91765 119722 94830
rect 120214 94830 120276 94890
rect 120582 94830 120684 94890
rect 121686 94830 121772 94890
rect 121984 94890 122044 95200
rect 122800 94890 122860 95200
rect 123208 94890 123268 95200
rect 121984 94830 122114 94890
rect 122800 94830 123034 94890
rect 119659 91764 119725 91765
rect 119659 91700 119660 91764
rect 119724 91700 119725 91764
rect 119659 91699 119725 91700
rect 120214 91221 120274 94830
rect 120582 91221 120642 94830
rect 121686 93533 121746 94830
rect 121683 93532 121749 93533
rect 121683 93468 121684 93532
rect 121748 93468 121749 93532
rect 121683 93467 121749 93468
rect 118187 91220 118253 91221
rect 118187 91156 118188 91220
rect 118252 91156 118253 91220
rect 118187 91155 118253 91156
rect 119291 91220 119357 91221
rect 119291 91156 119292 91220
rect 119356 91156 119357 91220
rect 119291 91155 119357 91156
rect 120211 91220 120277 91221
rect 120211 91156 120212 91220
rect 120276 91156 120277 91220
rect 120211 91155 120277 91156
rect 120579 91220 120645 91221
rect 120579 91156 120580 91220
rect 120644 91156 120645 91220
rect 120579 91155 120645 91156
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 86614 121574 93100
rect 122054 91221 122114 94830
rect 122974 93870 123034 94830
rect 122606 93810 123034 93870
rect 123158 94830 123268 94890
rect 124024 94890 124084 95200
rect 124432 94890 124492 95200
rect 125384 94890 125444 95200
rect 124024 94830 124138 94890
rect 124432 94830 124506 94890
rect 122606 91490 122666 93810
rect 123158 93533 123218 94830
rect 123155 93532 123221 93533
rect 123155 93468 123156 93532
rect 123220 93468 123221 93532
rect 123155 93467 123221 93468
rect 124078 92445 124138 94830
rect 124075 92444 124141 92445
rect 124075 92380 124076 92444
rect 124140 92380 124141 92444
rect 124075 92379 124141 92380
rect 122787 91492 122853 91493
rect 122787 91490 122788 91492
rect 122606 91430 122788 91490
rect 122787 91428 122788 91430
rect 122852 91428 122853 91492
rect 122787 91427 122853 91428
rect 124446 91357 124506 94830
rect 125366 94830 125444 94890
rect 125656 94890 125716 95200
rect 126472 94890 126532 95200
rect 125656 94830 125794 94890
rect 124443 91356 124509 91357
rect 124443 91292 124444 91356
rect 124508 91292 124509 91356
rect 124443 91291 124509 91292
rect 125366 91221 125426 94830
rect 125734 91357 125794 94830
rect 126470 94830 126532 94890
rect 126608 94890 126668 95200
rect 128104 94890 128164 95200
rect 126608 94830 126714 94890
rect 125731 91356 125797 91357
rect 125731 91292 125732 91356
rect 125796 91292 125797 91356
rect 125731 91291 125797 91292
rect 126470 91221 126530 94830
rect 126654 94077 126714 94830
rect 127574 94830 128164 94890
rect 129328 94890 129388 95200
rect 130688 94890 130748 95200
rect 131912 94890 131972 95200
rect 133136 94890 133196 95200
rect 129328 94830 129474 94890
rect 130688 94830 130762 94890
rect 131912 94830 132418 94890
rect 126651 94076 126717 94077
rect 126651 94012 126652 94076
rect 126716 94012 126717 94076
rect 126651 94011 126717 94012
rect 127574 91221 127634 94830
rect 122051 91220 122117 91221
rect 122051 91156 122052 91220
rect 122116 91156 122117 91220
rect 122051 91155 122117 91156
rect 125363 91220 125429 91221
rect 125363 91156 125364 91220
rect 125428 91156 125429 91220
rect 125363 91155 125429 91156
rect 126467 91220 126533 91221
rect 126467 91156 126468 91220
rect 126532 91156 126533 91220
rect 126467 91155 126533 91156
rect 127571 91220 127637 91221
rect 127571 91156 127572 91220
rect 127636 91156 127637 91220
rect 127571 91155 127637 91156
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 93100
rect 129414 91221 129474 94830
rect 130702 92173 130762 94830
rect 130699 92172 130765 92173
rect 130699 92108 130700 92172
rect 130764 92108 130765 92172
rect 130699 92107 130765 92108
rect 129411 91220 129477 91221
rect 129411 91156 129412 91220
rect 129476 91156 129477 91220
rect 129411 91155 129477 91156
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 61174 132134 93100
rect 132358 91221 132418 94830
rect 133094 94830 133196 94890
rect 134360 94890 134420 95200
rect 135584 94890 135644 95200
rect 151496 94890 151556 95200
rect 134360 94830 134442 94890
rect 135584 94830 136098 94890
rect 133094 93397 133154 94830
rect 134382 93669 134442 94830
rect 134379 93668 134445 93669
rect 134379 93604 134380 93668
rect 134444 93604 134445 93668
rect 134379 93603 134445 93604
rect 133091 93396 133157 93397
rect 133091 93332 133092 93396
rect 133156 93332 133157 93396
rect 133091 93331 133157 93332
rect 132355 91220 132421 91221
rect 132355 91156 132356 91220
rect 132420 91156 132421 91220
rect 132355 91155 132421 91156
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 64894 135854 93100
rect 136038 92445 136098 94830
rect 151494 94830 151556 94890
rect 151307 94756 151373 94757
rect 151307 94692 151308 94756
rect 151372 94692 151373 94756
rect 151307 94691 151373 94692
rect 136035 92444 136101 92445
rect 136035 92380 136036 92444
rect 136100 92380 136101 92444
rect 136035 92379 136101 92380
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 68614 139574 93100
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 79174 150134 93100
rect 151310 92445 151370 94691
rect 151307 92444 151373 92445
rect 151307 92380 151308 92444
rect 151372 92380 151373 92444
rect 151307 92379 151373 92380
rect 151494 91221 151554 94830
rect 151632 94210 151692 95200
rect 151768 94757 151828 95200
rect 151904 94890 151964 95200
rect 151904 94830 152106 94890
rect 151765 94756 151831 94757
rect 151765 94692 151766 94756
rect 151830 94692 151831 94756
rect 151765 94691 151831 94692
rect 151632 94150 151738 94210
rect 151678 91357 151738 94150
rect 151675 91356 151741 91357
rect 151675 91292 151676 91356
rect 151740 91292 151741 91356
rect 151675 91291 151741 91292
rect 152046 91221 152106 94830
rect 151491 91220 151557 91221
rect 151491 91156 151492 91220
rect 151556 91156 151557 91220
rect 151491 91155 151557 91156
rect 152043 91220 152109 91221
rect 152043 91156 152044 91220
rect 152108 91156 152109 91220
rect 152043 91155 152109 91156
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 82894 153854 93100
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 86614 157574 93100
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 93100
rect 166214 78437 166274 102443
rect 166395 95844 166461 95845
rect 166395 95780 166396 95844
rect 166460 95780 166461 95844
rect 166395 95779 166461 95780
rect 166398 81429 166458 95779
rect 166395 81428 166461 81429
rect 166395 81364 166396 81428
rect 166460 81364 166461 81428
rect 166395 81363 166461 81364
rect 166211 78436 166277 78437
rect 166211 78372 166212 78436
rect 166276 78372 166277 78436
rect 166211 78371 166277 78372
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 166950 8941 167010 175883
rect 167514 169174 168134 204618
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 168422 68509 168482 251363
rect 168419 68508 168485 68509
rect 168419 68444 168420 68508
rect 168484 68444 168485 68508
rect 168419 68443 168485 68444
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 166947 8940 167013 8941
rect 166947 8876 166948 8940
rect 167012 8876 167013 8940
rect 166947 8875 167013 8876
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 -3226 168134 24618
rect 169710 11661 169770 369003
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 180011 296036 180077 296037
rect 180011 295972 180012 296036
rect 180076 295972 180077 296036
rect 180011 295971 180077 295972
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 173019 275228 173085 275229
rect 173019 275164 173020 275228
rect 173084 275164 173085 275228
rect 173019 275163 173085 275164
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 169707 11660 169773 11661
rect 169707 11596 169708 11660
rect 169772 11596 169773 11660
rect 169707 11595 169773 11596
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 -5146 171854 28338
rect 173022 8941 173082 275163
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 180014 235789 180074 295971
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 180011 235788 180077 235789
rect 180011 235724 180012 235788
rect 180076 235724 180077 235788
rect 180011 235723 180077 235724
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 177251 185740 177317 185741
rect 177251 185676 177252 185740
rect 177316 185676 177317 185740
rect 177251 185675 177317 185676
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 173019 8940 173085 8941
rect 173019 8876 173020 8940
rect 173084 8876 173085 8940
rect 173019 8875 173085 8876
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 177254 4997 177314 185675
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 177251 4996 177317 4997
rect 177251 4932 177252 4996
rect 177316 4932 177317 4996
rect 177251 4931 177317 4932
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 188291 357644 188357 357645
rect 188291 357580 188292 357644
rect 188356 357580 188357 357644
rect 188291 357579 188357 357580
rect 186819 350708 186885 350709
rect 186819 350644 186820 350708
rect 186884 350644 186885 350708
rect 186819 350643 186885 350644
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 186822 237149 186882 350643
rect 187003 308548 187069 308549
rect 187003 308484 187004 308548
rect 187068 308484 187069 308548
rect 187003 308483 187069 308484
rect 187006 247213 187066 308483
rect 187003 247212 187069 247213
rect 187003 247148 187004 247212
rect 187068 247148 187069 247212
rect 187003 247147 187069 247148
rect 186819 237148 186885 237149
rect 186819 237084 186820 237148
rect 186884 237084 186885 237148
rect 186819 237083 186885 237084
rect 188294 235789 188354 357579
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 197859 356284 197925 356285
rect 197859 356220 197860 356284
rect 197924 356220 197925 356284
rect 197859 356219 197925 356220
rect 196939 349348 197005 349349
rect 196939 349284 196940 349348
rect 197004 349284 197005 349348
rect 196939 349283 197005 349284
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 191603 317388 191669 317389
rect 191603 317324 191604 317388
rect 191668 317324 191669 317388
rect 191603 317323 191669 317324
rect 191606 316165 191666 317323
rect 191603 316164 191669 316165
rect 191603 316100 191604 316164
rect 191668 316100 191669 316164
rect 191603 316099 191669 316100
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 188291 235788 188357 235789
rect 188291 235724 188292 235788
rect 188356 235724 188357 235788
rect 188291 235723 188357 235724
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 189234 226894 189854 262338
rect 191051 260132 191117 260133
rect 191051 260068 191052 260132
rect 191116 260068 191117 260132
rect 191051 260067 191117 260068
rect 191054 234429 191114 260067
rect 191606 259045 191666 316099
rect 192954 302614 193574 338058
rect 195099 313308 195165 313309
rect 195099 313244 195100 313308
rect 195164 313244 195165 313308
rect 195099 313243 195165 313244
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 191603 259044 191669 259045
rect 191603 258980 191604 259044
rect 191668 258980 191669 259044
rect 191603 258979 191669 258980
rect 191051 234428 191117 234429
rect 191051 234364 191052 234428
rect 191116 234364 191117 234428
rect 191051 234363 191117 234364
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 186819 214572 186885 214573
rect 186819 214508 186820 214572
rect 186884 214508 186885 214572
rect 186819 214507 186885 214508
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 186822 14517 186882 214507
rect 189234 190894 189854 226338
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 191051 223004 191117 223005
rect 191051 222940 191052 223004
rect 191116 222940 191117 223004
rect 191051 222939 191117 222940
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 186819 14516 186885 14517
rect 186819 14452 186820 14516
rect 186884 14452 186885 14516
rect 186819 14451 186885 14452
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 191054 3365 191114 222939
rect 192954 194614 193574 230058
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 191051 3364 191117 3365
rect 191051 3300 191052 3364
rect 191116 3300 191117 3364
rect 191051 3299 191117 3300
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 195102 11661 195162 313243
rect 195283 242996 195349 242997
rect 195283 242932 195284 242996
rect 195348 242932 195349 242996
rect 195283 242931 195349 242932
rect 195286 235245 195346 242931
rect 196942 237285 197002 349283
rect 197862 281621 197922 356219
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199331 291412 199397 291413
rect 199331 291348 199332 291412
rect 199396 291348 199397 291412
rect 199331 291347 199397 291348
rect 197859 281620 197925 281621
rect 197859 281556 197860 281620
rect 197924 281556 197925 281620
rect 197859 281555 197925 281556
rect 199334 279581 199394 291347
rect 199794 286182 200414 308898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 200619 288692 200685 288693
rect 200619 288628 200620 288692
rect 200684 288628 200685 288692
rect 200619 288627 200685 288628
rect 200067 282572 200133 282573
rect 200067 282508 200068 282572
rect 200132 282570 200133 282572
rect 200622 282570 200682 288627
rect 203514 286182 204134 312618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 286182 207854 316338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 212579 354924 212645 354925
rect 212579 354860 212580 354924
rect 212644 354860 212645 354924
rect 212579 354859 212645 354860
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 286182 211574 320058
rect 211659 287196 211725 287197
rect 211659 287132 211660 287196
rect 211724 287132 211725 287196
rect 211659 287131 211725 287132
rect 205403 283932 205469 283933
rect 205403 283868 205404 283932
rect 205468 283868 205469 283932
rect 205403 283867 205469 283868
rect 206875 283932 206941 283933
rect 206875 283868 206876 283932
rect 206940 283868 206941 283932
rect 206875 283867 206941 283868
rect 209635 283932 209701 283933
rect 209635 283868 209636 283932
rect 209700 283868 209701 283932
rect 209635 283867 209701 283868
rect 200132 282510 200682 282570
rect 200132 282508 200133 282510
rect 200067 282507 200133 282508
rect 199331 279580 199397 279581
rect 199331 279516 199332 279580
rect 199396 279516 199397 279580
rect 199331 279515 199397 279516
rect 204408 255454 204728 255486
rect 197123 255236 197189 255237
rect 197123 255172 197124 255236
rect 197188 255172 197189 255236
rect 197123 255171 197189 255172
rect 204408 255218 204450 255454
rect 204686 255218 204728 255454
rect 196939 237284 197005 237285
rect 196939 237220 196940 237284
rect 197004 237220 197005 237284
rect 196939 237219 197005 237220
rect 195283 235244 195349 235245
rect 195283 235180 195284 235244
rect 195348 235180 195349 235244
rect 195283 235179 195349 235180
rect 197126 90405 197186 255171
rect 204408 255134 204728 255218
rect 204408 254898 204450 255134
rect 204686 254898 204728 255134
rect 204408 254866 204728 254898
rect 199883 251972 199949 251973
rect 199883 251908 199884 251972
rect 199948 251908 199949 251972
rect 199883 251907 199949 251908
rect 199886 251190 199946 251907
rect 199886 251130 200682 251190
rect 199515 249796 199581 249797
rect 199515 249732 199516 249796
rect 199580 249732 199581 249796
rect 199515 249731 199581 249732
rect 199518 178805 199578 249731
rect 199883 246532 199949 246533
rect 199883 246468 199884 246532
rect 199948 246468 199949 246532
rect 199883 246467 199949 246468
rect 199886 243541 199946 246467
rect 199883 243540 199949 243541
rect 199883 243476 199884 243540
rect 199948 243476 199949 243540
rect 199883 243475 199949 243476
rect 199886 239461 199946 243475
rect 199883 239460 199949 239461
rect 199883 239396 199884 239460
rect 199948 239396 199949 239460
rect 199883 239395 199949 239396
rect 199794 237454 200414 238182
rect 200622 237965 200682 251130
rect 200619 237964 200685 237965
rect 200619 237900 200620 237964
rect 200684 237900 200685 237964
rect 200619 237899 200685 237900
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199515 178804 199581 178805
rect 199515 178740 199516 178804
rect 199580 178740 199581 178804
rect 199515 178739 199581 178740
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 197123 90404 197189 90405
rect 197123 90340 197124 90404
rect 197188 90340 197189 90404
rect 197123 90339 197189 90340
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 195099 11660 195165 11661
rect 195099 11596 195100 11660
rect 195164 11596 195165 11660
rect 195099 11595 195165 11596
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 205174 204134 238182
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 203514 61174 204134 96618
rect 205406 95165 205466 283867
rect 206878 185741 206938 283867
rect 207234 208894 207854 238182
rect 209638 215933 209698 283867
rect 211662 238373 211722 287131
rect 212582 238645 212642 354859
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 214235 308412 214301 308413
rect 214235 308348 214236 308412
rect 214300 308348 214301 308412
rect 214235 308347 214301 308348
rect 214051 283932 214117 283933
rect 214051 283868 214052 283932
rect 214116 283868 214117 283932
rect 214051 283867 214117 283868
rect 212579 238644 212645 238645
rect 212579 238580 212580 238644
rect 212644 238580 212645 238644
rect 212579 238579 212645 238580
rect 211659 238372 211725 238373
rect 211659 238308 211660 238372
rect 211724 238308 211725 238372
rect 211659 238307 211725 238308
rect 209635 215932 209701 215933
rect 209635 215868 209636 215932
rect 209700 215868 209701 215932
rect 209635 215867 209701 215868
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 206875 185740 206941 185741
rect 206875 185676 206876 185740
rect 206940 185676 206941 185740
rect 206875 185675 206941 185676
rect 207234 172894 207854 208338
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 205403 95164 205469 95165
rect 205403 95100 205404 95164
rect 205468 95100 205469 95164
rect 205403 95099 205469 95100
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 212614 211574 238182
rect 213131 237420 213197 237421
rect 213131 237356 213132 237420
rect 213196 237356 213197 237420
rect 213131 237355 213197 237356
rect 213134 213213 213194 237355
rect 214054 234701 214114 283867
rect 214238 240141 214298 308347
rect 217794 291454 218414 326898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 222331 365804 222397 365805
rect 222331 365740 222332 365804
rect 222396 365740 222397 365804
rect 222331 365739 222397 365740
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221043 296852 221109 296853
rect 221043 296788 221044 296852
rect 221108 296788 221109 296852
rect 221043 296787 221109 296788
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 286182 218414 290898
rect 215339 283932 215405 283933
rect 215339 283868 215340 283932
rect 215404 283868 215405 283932
rect 215339 283867 215405 283868
rect 217179 283932 217245 283933
rect 217179 283868 217180 283932
rect 217244 283868 217245 283932
rect 217179 283867 217245 283868
rect 214235 240140 214301 240141
rect 214235 240076 214236 240140
rect 214300 240076 214301 240140
rect 214235 240075 214301 240076
rect 214051 234700 214117 234701
rect 214051 234636 214052 234700
rect 214116 234636 214117 234700
rect 214051 234635 214117 234636
rect 215342 213893 215402 283867
rect 217182 231845 217242 283867
rect 219768 273454 220088 273486
rect 219768 273218 219810 273454
rect 220046 273218 220088 273454
rect 219768 273134 220088 273218
rect 219768 272898 219810 273134
rect 220046 272898 220088 273134
rect 219768 272866 220088 272898
rect 221046 240141 221106 296787
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 286182 222134 294618
rect 221043 240140 221109 240141
rect 221043 240076 221044 240140
rect 221108 240076 221109 240140
rect 221043 240075 221109 240076
rect 222334 238645 222394 365739
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 286182 225854 298338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 232451 354788 232517 354789
rect 232451 354724 232452 354788
rect 232516 354724 232517 354788
rect 232451 354723 232517 354724
rect 230427 341052 230493 341053
rect 230427 340988 230428 341052
rect 230492 340988 230493 341052
rect 230427 340987 230493 340988
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 286182 229574 302058
rect 226931 285972 226997 285973
rect 226931 285908 226932 285972
rect 226996 285908 226997 285972
rect 226931 285907 226997 285908
rect 224907 285700 224973 285701
rect 224907 285636 224908 285700
rect 224972 285636 224973 285700
rect 224907 285635 224973 285636
rect 224723 283932 224789 283933
rect 224723 283868 224724 283932
rect 224788 283868 224789 283932
rect 224723 283867 224789 283868
rect 222331 238644 222397 238645
rect 222331 238580 222332 238644
rect 222396 238580 222397 238644
rect 222331 238579 222397 238580
rect 217179 231844 217245 231845
rect 217179 231780 217180 231844
rect 217244 231780 217245 231844
rect 217179 231779 217245 231780
rect 217794 219454 218414 238182
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 215339 213892 215405 213893
rect 215339 213828 215340 213892
rect 215404 213828 215405 213892
rect 215339 213827 215405 213828
rect 213131 213212 213197 213213
rect 213131 213148 213132 213212
rect 213196 213148 213197 213212
rect 213131 213147 213197 213148
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210954 176614 211574 212058
rect 217794 183454 218414 218898
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 178000 218414 182898
rect 221514 223174 222134 238182
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221514 187174 222134 222618
rect 224726 213349 224786 283867
rect 224910 240141 224970 285635
rect 226379 283932 226445 283933
rect 226379 283868 226380 283932
rect 226444 283868 226445 283932
rect 226379 283867 226445 283868
rect 224907 240140 224973 240141
rect 224907 240076 224908 240140
rect 224972 240076 224973 240140
rect 224907 240075 224973 240076
rect 225234 226894 225854 238182
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 224723 213348 224789 213349
rect 224723 213284 224724 213348
rect 224788 213284 224789 213348
rect 224723 213283 224789 213284
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 178000 222134 186618
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 178000 225854 190338
rect 226382 189957 226442 283867
rect 226934 196077 226994 285907
rect 228771 283932 228837 283933
rect 228771 283868 228772 283932
rect 228836 283868 228837 283932
rect 228771 283867 228837 283868
rect 229691 283932 229757 283933
rect 229691 283868 229692 283932
rect 229756 283868 229757 283932
rect 229691 283867 229757 283868
rect 226931 196076 226997 196077
rect 226931 196012 226932 196076
rect 226996 196012 226997 196076
rect 226931 196011 226997 196012
rect 226379 189956 226445 189957
rect 226379 189892 226380 189956
rect 226444 189892 226445 189956
rect 226379 189891 226445 189892
rect 228219 189820 228285 189821
rect 228219 189756 228220 189820
rect 228284 189756 228285 189820
rect 228219 189755 228285 189756
rect 227667 185740 227733 185741
rect 227667 185676 227668 185740
rect 227732 185676 227733 185740
rect 227667 185675 227733 185676
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 227670 174450 227730 185675
rect 228222 175130 228282 189755
rect 228774 185741 228834 283867
rect 229694 240141 229754 283867
rect 230430 240141 230490 340987
rect 231715 283932 231781 283933
rect 231715 283868 231716 283932
rect 231780 283868 231781 283932
rect 231715 283867 231781 283868
rect 229691 240140 229757 240141
rect 229691 240076 229692 240140
rect 229756 240076 229757 240140
rect 229691 240075 229757 240076
rect 230427 240140 230493 240141
rect 230427 240076 230428 240140
rect 230492 240076 230493 240140
rect 230427 240075 230493 240076
rect 228954 230614 229574 238182
rect 231718 233205 231778 283867
rect 232454 238645 232514 354723
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 237419 325004 237485 325005
rect 237419 324940 237420 325004
rect 237484 324940 237485 325004
rect 237419 324939 237485 324940
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 233187 288692 233253 288693
rect 233187 288628 233188 288692
rect 233252 288628 233253 288692
rect 233187 288627 233253 288628
rect 232451 238644 232517 238645
rect 232451 238580 232452 238644
rect 232516 238580 232517 238644
rect 232451 238579 232517 238580
rect 231715 233204 231781 233205
rect 231715 233140 231716 233204
rect 231780 233140 231781 233204
rect 231715 233139 231781 233140
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 231899 211988 231965 211989
rect 231899 211924 231900 211988
rect 231964 211924 231965 211988
rect 231899 211923 231965 211924
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228771 185740 228837 185741
rect 228771 185676 228772 185740
rect 228836 185676 228837 185740
rect 228771 185675 228837 185676
rect 228954 178000 229574 194058
rect 229691 191180 229757 191181
rect 229691 191116 229692 191180
rect 229756 191116 229757 191180
rect 229691 191115 229757 191116
rect 229323 176764 229389 176765
rect 229323 176700 229324 176764
rect 229388 176700 229389 176764
rect 229323 176699 229389 176700
rect 229139 175132 229205 175133
rect 229139 175130 229140 175132
rect 228222 175070 229140 175130
rect 229139 175068 229140 175070
rect 229204 175068 229205 175132
rect 229139 175067 229205 175068
rect 227670 174390 229202 174450
rect 229142 174317 229202 174390
rect 229139 174316 229205 174317
rect 229139 174252 229140 174316
rect 229204 174252 229205 174316
rect 229139 174251 229205 174252
rect 229326 173770 229386 176699
rect 229694 175133 229754 191115
rect 230427 181660 230493 181661
rect 230427 181596 230428 181660
rect 230492 181596 230493 181660
rect 230427 181595 230493 181596
rect 229691 175132 229757 175133
rect 229691 175068 229692 175132
rect 229756 175068 229757 175132
rect 229691 175067 229757 175068
rect 229507 174996 229573 174997
rect 229507 174932 229508 174996
rect 229572 174932 229573 174996
rect 229507 174931 229573 174932
rect 229142 173710 229386 173770
rect 221207 165454 221527 165486
rect 221207 165218 221249 165454
rect 221485 165218 221527 165454
rect 221207 165134 221527 165218
rect 221207 164898 221249 165134
rect 221485 164898 221527 165134
rect 221207 164866 221527 164898
rect 224471 165454 224791 165486
rect 224471 165218 224513 165454
rect 224749 165218 224791 165454
rect 224471 165134 224791 165218
rect 224471 164898 224513 165134
rect 224749 164898 224791 165134
rect 224471 164866 224791 164898
rect 219575 147454 219895 147486
rect 219575 147218 219617 147454
rect 219853 147218 219895 147454
rect 219575 147134 219895 147218
rect 219575 146898 219617 147134
rect 219853 146898 219895 147134
rect 219575 146866 219895 146898
rect 222839 147454 223159 147486
rect 222839 147218 222881 147454
rect 223117 147218 223159 147454
rect 222839 147134 223159 147218
rect 222839 146898 222881 147134
rect 223117 146898 223159 147134
rect 222839 146866 223159 146898
rect 226103 147454 226423 147486
rect 226103 147218 226145 147454
rect 226381 147218 226423 147454
rect 226103 147134 226423 147218
rect 226103 146898 226145 147134
rect 226381 146898 226423 147134
rect 226103 146866 226423 146898
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 229142 137325 229202 173710
rect 229510 161490 229570 174931
rect 229326 161430 229570 161490
rect 229326 146301 229386 161430
rect 230430 149701 230490 181595
rect 230611 176628 230677 176629
rect 230611 176564 230612 176628
rect 230676 176564 230677 176628
rect 230611 176563 230677 176564
rect 230614 155821 230674 176563
rect 231902 161533 231962 211923
rect 232083 188460 232149 188461
rect 232083 188396 232084 188460
rect 232148 188396 232149 188460
rect 232083 188395 232149 188396
rect 231899 161532 231965 161533
rect 231899 161468 231900 161532
rect 231964 161468 231965 161532
rect 231899 161467 231965 161468
rect 230611 155820 230677 155821
rect 230611 155756 230612 155820
rect 230676 155756 230677 155820
rect 230611 155755 230677 155756
rect 230979 155276 231045 155277
rect 230979 155212 230980 155276
rect 231044 155212 231045 155276
rect 230979 155211 231045 155212
rect 230427 149700 230493 149701
rect 230427 149636 230428 149700
rect 230492 149636 230493 149700
rect 230427 149635 230493 149636
rect 229323 146300 229389 146301
rect 229323 146236 229324 146300
rect 229388 146236 229389 146300
rect 229323 146235 229389 146236
rect 229139 137324 229205 137325
rect 229139 137260 229140 137324
rect 229204 137260 229205 137324
rect 229139 137259 229205 137260
rect 230982 133517 231042 155211
rect 232086 152557 232146 188395
rect 233190 154869 233250 288627
rect 235794 286182 236414 308898
rect 236499 285700 236565 285701
rect 236499 285636 236500 285700
rect 236564 285636 236565 285700
rect 236499 285635 236565 285636
rect 236502 283933 236562 285635
rect 236499 283932 236565 283933
rect 236499 283868 236500 283932
rect 236564 283868 236565 283932
rect 236499 283867 236565 283868
rect 235128 255454 235448 255486
rect 235128 255218 235170 255454
rect 235406 255218 235448 255454
rect 235128 255134 235448 255218
rect 235128 254898 235170 255134
rect 235406 254898 235448 255134
rect 235128 254866 235448 254898
rect 235794 237454 236414 238182
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 233371 233204 233437 233205
rect 233371 233140 233372 233204
rect 233436 233140 233437 233204
rect 233371 233139 233437 233140
rect 233187 154868 233253 154869
rect 233187 154804 233188 154868
rect 233252 154804 233253 154868
rect 233187 154803 233253 154804
rect 232083 152556 232149 152557
rect 232083 152492 232084 152556
rect 232148 152492 232149 152556
rect 232083 152491 232149 152492
rect 231163 140044 231229 140045
rect 231163 139980 231164 140044
rect 231228 139980 231229 140044
rect 231163 139979 231229 139980
rect 230979 133516 231045 133517
rect 230979 133452 230980 133516
rect 231044 133452 231045 133516
rect 230979 133451 231045 133452
rect 229691 132836 229757 132837
rect 229691 132772 229692 132836
rect 229756 132772 229757 132836
rect 229691 132771 229757 132772
rect 221207 129454 221527 129486
rect 221207 129218 221249 129454
rect 221485 129218 221527 129454
rect 221207 129134 221527 129218
rect 221207 128898 221249 129134
rect 221485 128898 221527 129134
rect 221207 128866 221527 128898
rect 224471 129454 224791 129486
rect 224471 129218 224513 129454
rect 224749 129218 224791 129454
rect 224471 129134 224791 129218
rect 224471 128898 224513 129134
rect 224749 128898 224791 129134
rect 224471 128866 224791 128898
rect 219575 111454 219895 111486
rect 219575 111218 219617 111454
rect 219853 111218 219895 111454
rect 219575 111134 219895 111218
rect 219575 110898 219617 111134
rect 219853 110898 219895 111134
rect 219575 110866 219895 110898
rect 222839 111454 223159 111486
rect 222839 111218 222881 111454
rect 223117 111218 223159 111454
rect 222839 111134 223159 111218
rect 222839 110898 222881 111134
rect 223117 110898 223159 111134
rect 222839 110866 223159 110898
rect 226103 111454 226423 111486
rect 226103 111218 226145 111454
rect 226381 111218 226423 111454
rect 226103 111134 226423 111218
rect 226103 110898 226145 111134
rect 226381 110898 226423 111134
rect 226103 110866 226423 110898
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 229139 97204 229205 97205
rect 229139 97140 229140 97204
rect 229204 97140 229205 97204
rect 229139 97139 229205 97140
rect 229142 96930 229202 97139
rect 219206 96870 220922 96930
rect 219206 95981 219266 96870
rect 219203 95980 219269 95981
rect 219203 95916 219204 95980
rect 219268 95916 219269 95980
rect 219203 95915 219269 95916
rect 219203 95844 219269 95845
rect 219203 95780 219204 95844
rect 219268 95780 219269 95844
rect 219203 95779 219269 95780
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 94000
rect 219206 86869 219266 95779
rect 219203 86868 219269 86869
rect 219203 86804 219204 86868
rect 219268 86804 219269 86868
rect 219203 86803 219269 86804
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 220862 43485 220922 96870
rect 228590 96870 229202 96930
rect 228590 95573 228650 96870
rect 229139 96660 229205 96661
rect 229139 96630 229140 96660
rect 228958 96596 229140 96630
rect 229204 96596 229205 96660
rect 228958 96595 229205 96596
rect 228958 96570 229202 96595
rect 224907 95572 224973 95573
rect 224907 95508 224908 95572
rect 224972 95508 224973 95572
rect 224907 95507 224973 95508
rect 228587 95572 228653 95573
rect 228587 95508 228588 95572
rect 228652 95508 228653 95572
rect 228587 95507 228653 95508
rect 221514 79174 222134 94000
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 220859 43484 220925 43485
rect 220859 43420 220860 43484
rect 220924 43420 220925 43484
rect 220859 43419 220925 43420
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 78618
rect 224910 68237 224970 95507
rect 228958 94890 229018 96570
rect 227670 94830 229018 94890
rect 225234 82894 225854 94000
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 224907 68236 224973 68237
rect 224907 68172 224908 68236
rect 224972 68172 224973 68236
rect 224907 68171 224973 68172
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 227670 22677 227730 94830
rect 228954 86614 229574 94000
rect 229694 91765 229754 132771
rect 231166 131613 231226 139979
rect 233374 139773 233434 233139
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 234659 196076 234725 196077
rect 234659 196012 234660 196076
rect 234724 196012 234725 196076
rect 234659 196011 234725 196012
rect 233555 155956 233621 155957
rect 233555 155892 233556 155956
rect 233620 155892 233621 155956
rect 233555 155891 233621 155892
rect 233558 145349 233618 155891
rect 233555 145348 233621 145349
rect 233555 145284 233556 145348
rect 233620 145284 233621 145348
rect 233555 145283 233621 145284
rect 233739 145348 233805 145349
rect 233739 145284 233740 145348
rect 233804 145284 233805 145348
rect 233739 145283 233805 145284
rect 233371 139772 233437 139773
rect 233371 139708 233372 139772
rect 233436 139708 233437 139772
rect 233371 139707 233437 139708
rect 232451 138684 232517 138685
rect 232451 138620 232452 138684
rect 232516 138620 232517 138684
rect 232451 138619 232517 138620
rect 231163 131612 231229 131613
rect 231163 131548 231164 131612
rect 231228 131548 231229 131612
rect 231163 131547 231229 131548
rect 230979 111212 231045 111213
rect 230979 111148 230980 111212
rect 231044 111148 231045 111212
rect 230979 111147 231045 111148
rect 230982 98973 231042 111147
rect 230979 98972 231045 98973
rect 230979 98908 230980 98972
rect 231044 98908 231045 98972
rect 230979 98907 231045 98908
rect 232454 98021 232514 138619
rect 233742 103325 233802 145283
rect 234662 139229 234722 196011
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 236502 165205 236562 283867
rect 237422 240141 237482 324939
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 286182 240134 312618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 244227 371380 244293 371381
rect 244227 371316 244228 371380
rect 244292 371316 244293 371380
rect 244227 371315 244293 371316
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 242939 306508 243005 306509
rect 242939 306444 242940 306508
rect 243004 306444 243005 306508
rect 242939 306443 243005 306444
rect 241651 297396 241717 297397
rect 241651 297332 241652 297396
rect 241716 297332 241717 297396
rect 241651 297331 241717 297332
rect 240363 285972 240429 285973
rect 240363 285908 240364 285972
rect 240428 285908 240429 285972
rect 240363 285907 240429 285908
rect 238523 285836 238589 285837
rect 238523 285772 238524 285836
rect 238588 285772 238589 285836
rect 238523 285771 238589 285772
rect 237419 240140 237485 240141
rect 237419 240076 237420 240140
rect 237484 240076 237485 240140
rect 237419 240075 237485 240076
rect 237422 168741 237482 240075
rect 237603 181524 237669 181525
rect 237603 181460 237604 181524
rect 237668 181460 237669 181524
rect 237603 181459 237669 181460
rect 237419 168740 237485 168741
rect 237419 168676 237420 168740
rect 237484 168676 237485 168740
rect 237419 168675 237485 168676
rect 236499 165204 236565 165205
rect 236499 165140 236500 165204
rect 236564 165140 236565 165204
rect 236499 165139 236565 165140
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 234659 139228 234725 139229
rect 234659 139164 234660 139228
rect 234724 139164 234725 139228
rect 234659 139163 234725 139164
rect 235794 129454 236414 164898
rect 237606 149293 237666 181459
rect 238526 173365 238586 285771
rect 239514 205174 240134 238182
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 238523 173364 238589 173365
rect 238523 173300 238524 173364
rect 238588 173300 238589 173364
rect 238523 173299 238589 173300
rect 239514 169174 240134 204618
rect 240366 173909 240426 285907
rect 241654 238645 241714 297331
rect 242942 279170 243002 306443
rect 243234 286182 243854 316338
rect 243491 279172 243557 279173
rect 243491 279170 243492 279172
rect 242942 279110 243492 279170
rect 243491 279108 243492 279110
rect 243556 279108 243557 279172
rect 243491 279107 243557 279108
rect 244230 275637 244290 371315
rect 246954 356614 247574 392058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 252507 369884 252573 369885
rect 252507 369820 252508 369884
rect 252572 369820 252573 369884
rect 252507 369819 252573 369820
rect 249747 357508 249813 357509
rect 249747 357444 249748 357508
rect 249812 357444 249813 357508
rect 249747 357443 249813 357444
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 248459 350572 248525 350573
rect 248459 350508 248460 350572
rect 248524 350508 248525 350572
rect 248459 350507 248525 350508
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 284614 247574 320058
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 244227 275636 244293 275637
rect 244227 275572 244228 275636
rect 244292 275572 244293 275636
rect 244227 275571 244293 275572
rect 246954 248614 247574 284058
rect 248462 249525 248522 350507
rect 249750 263941 249810 357443
rect 249931 265708 249997 265709
rect 249931 265644 249932 265708
rect 249996 265644 249997 265708
rect 249931 265643 249997 265644
rect 249747 263940 249813 263941
rect 249747 263876 249748 263940
rect 249812 263876 249813 263940
rect 249747 263875 249813 263876
rect 248459 249524 248525 249525
rect 248459 249460 248460 249524
rect 248524 249460 248525 249524
rect 248459 249459 248525 249460
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 243491 246260 243557 246261
rect 243491 246196 243492 246260
rect 243556 246196 243557 246260
rect 243491 246195 243557 246196
rect 243494 238770 243554 246195
rect 245883 242996 245949 242997
rect 245883 242932 245884 242996
rect 245948 242932 245949 242996
rect 245883 242931 245949 242932
rect 245699 240276 245765 240277
rect 245699 240212 245700 240276
rect 245764 240212 245765 240276
rect 245699 240211 245765 240212
rect 242942 238710 243554 238770
rect 241651 238644 241717 238645
rect 241651 238580 241652 238644
rect 241716 238580 241717 238644
rect 241651 238579 241717 238580
rect 242942 232525 243002 238710
rect 242939 232524 243005 232525
rect 242939 232460 242940 232524
rect 243004 232460 243005 232524
rect 242939 232459 243005 232460
rect 243234 208894 243854 238182
rect 245702 227629 245762 240211
rect 245886 234565 245946 242931
rect 245883 234564 245949 234565
rect 245883 234500 245884 234564
rect 245948 234500 245949 234564
rect 245883 234499 245949 234500
rect 245699 227628 245765 227629
rect 245699 227564 245700 227628
rect 245764 227564 245765 227628
rect 245699 227563 245765 227564
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 240547 189820 240613 189821
rect 240547 189756 240548 189820
rect 240612 189756 240613 189820
rect 240547 189755 240613 189756
rect 240363 173908 240429 173909
rect 240363 173844 240364 173908
rect 240428 173844 240429 173908
rect 240363 173843 240429 173844
rect 240363 172412 240429 172413
rect 240363 172348 240364 172412
rect 240428 172348 240429 172412
rect 240363 172347 240429 172348
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 237603 149292 237669 149293
rect 237603 149228 237604 149292
rect 237668 149228 237669 149292
rect 237603 149227 237669 149228
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 233739 103324 233805 103325
rect 233739 103260 233740 103324
rect 233804 103260 233805 103324
rect 233739 103259 233805 103260
rect 232451 98020 232517 98021
rect 232451 97956 232452 98020
rect 232516 97956 232517 98020
rect 232451 97955 232517 97956
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 229691 91764 229757 91765
rect 229691 91700 229692 91764
rect 229756 91700 229757 91764
rect 229691 91699 229757 91700
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 227667 22676 227733 22677
rect 227667 22612 227668 22676
rect 227732 22612 227733 22676
rect 227667 22611 227733 22612
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 133174 240134 168618
rect 240366 143309 240426 172347
rect 240550 147253 240610 189755
rect 241467 188596 241533 188597
rect 241467 188532 241468 188596
rect 241532 188532 241533 188596
rect 241467 188531 241533 188532
rect 241470 151061 241530 188531
rect 241651 176084 241717 176085
rect 241651 176020 241652 176084
rect 241716 176020 241717 176084
rect 241651 176019 241717 176020
rect 241654 171150 241714 176019
rect 243234 172894 243854 208338
rect 246954 212614 247574 248058
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 244227 205188 244293 205189
rect 244227 205124 244228 205188
rect 244292 205124 244293 205188
rect 244227 205123 244293 205124
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 241654 171090 241898 171150
rect 241467 151060 241533 151061
rect 241467 150996 241468 151060
rect 241532 150996 241533 151060
rect 241467 150995 241533 150996
rect 241838 149701 241898 171090
rect 241835 149700 241901 149701
rect 241835 149636 241836 149700
rect 241900 149636 241901 149700
rect 241835 149635 241901 149636
rect 240547 147252 240613 147253
rect 240547 147188 240548 147252
rect 240612 147188 240613 147252
rect 240547 147187 240613 147188
rect 240363 143308 240429 143309
rect 240363 143244 240364 143308
rect 240428 143244 240429 143308
rect 240363 143243 240429 143244
rect 243234 136894 243854 172338
rect 244230 156773 244290 205123
rect 244411 187100 244477 187101
rect 244411 187036 244412 187100
rect 244476 187036 244477 187100
rect 244411 187035 244477 187036
rect 244414 162213 244474 187035
rect 246251 185604 246317 185605
rect 246251 185540 246252 185604
rect 246316 185540 246317 185604
rect 246251 185539 246317 185540
rect 244411 162212 244477 162213
rect 244411 162148 244412 162212
rect 244476 162148 244477 162212
rect 244411 162147 244477 162148
rect 244227 156772 244293 156773
rect 244227 156708 244228 156772
rect 244292 156708 244293 156772
rect 244227 156707 244293 156708
rect 244779 141404 244845 141405
rect 244779 141340 244780 141404
rect 244844 141340 244845 141404
rect 244779 141339 244845 141340
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 242203 135828 242269 135829
rect 242203 135764 242204 135828
rect 242268 135764 242269 135828
rect 242203 135763 242269 135764
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 242019 132972 242085 132973
rect 242019 132908 242020 132972
rect 242084 132908 242085 132972
rect 242019 132907 242085 132908
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 240731 120868 240797 120869
rect 240731 120804 240732 120868
rect 240796 120804 240797 120868
rect 240731 120803 240797 120804
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 240734 40629 240794 120803
rect 242022 53141 242082 132907
rect 242206 91901 242266 135763
rect 243234 100894 243854 136338
rect 244782 102101 244842 141339
rect 244779 102100 244845 102101
rect 244779 102036 244780 102100
rect 244844 102036 244845 102100
rect 244779 102035 244845 102036
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 242203 91900 242269 91901
rect 242203 91836 242204 91900
rect 242268 91836 242269 91900
rect 242203 91835 242269 91836
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 242019 53140 242085 53141
rect 242019 53076 242020 53140
rect 242084 53076 242085 53140
rect 242019 53075 242085 53076
rect 240731 40628 240797 40629
rect 240731 40564 240732 40628
rect 240796 40564 240797 40628
rect 240731 40563 240797 40564
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 246254 3501 246314 185539
rect 246954 176614 247574 212058
rect 249011 183020 249077 183021
rect 249011 182956 249012 183020
rect 249076 182956 249077 183020
rect 249011 182955 249077 182956
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 246251 3500 246317 3501
rect 246251 3436 246252 3500
rect 246316 3436 246317 3500
rect 246251 3435 246317 3436
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 249014 3501 249074 182955
rect 249934 152013 249994 265643
rect 252510 234565 252570 369819
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 252507 234564 252573 234565
rect 252507 234500 252508 234564
rect 252572 234500 252573 234564
rect 252507 234499 252573 234500
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253059 200700 253125 200701
rect 253059 200636 253060 200700
rect 253124 200636 253125 200700
rect 253059 200635 253125 200636
rect 251219 187236 251285 187237
rect 251219 187172 251220 187236
rect 251284 187172 251285 187236
rect 251219 187171 251285 187172
rect 249931 152012 249997 152013
rect 249931 151948 249932 152012
rect 249996 151948 249997 152012
rect 249931 151947 249997 151948
rect 251222 140181 251282 187171
rect 251219 140180 251285 140181
rect 251219 140116 251220 140180
rect 251284 140116 251285 140180
rect 251219 140115 251285 140116
rect 250299 134468 250365 134469
rect 250299 134404 250300 134468
rect 250364 134404 250365 134468
rect 250299 134403 250365 134404
rect 250302 107541 250362 134403
rect 251771 129028 251837 129029
rect 251771 128964 251772 129028
rect 251836 128964 251837 129028
rect 251771 128963 251837 128964
rect 250299 107540 250365 107541
rect 250299 107476 250300 107540
rect 250364 107476 250365 107540
rect 250299 107475 250365 107476
rect 251774 106861 251834 128963
rect 251771 106860 251837 106861
rect 251771 106796 251772 106860
rect 251836 106796 251837 106860
rect 251771 106795 251837 106796
rect 253062 4045 253122 200635
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 255819 127260 255885 127261
rect 255819 127196 255820 127260
rect 255884 127196 255885 127260
rect 255819 127195 255885 127196
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253059 4044 253125 4045
rect 253059 3980 253060 4044
rect 253124 3980 253125 4044
rect 253059 3979 253125 3980
rect 249011 3500 249077 3501
rect 249011 3436 249012 3500
rect 249076 3436 249077 3500
rect 249011 3435 249077 3436
rect 253794 3454 254414 38898
rect 255822 29613 255882 127195
rect 257514 115174 258134 150618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 260051 140180 260117 140181
rect 260051 140116 260052 140180
rect 260116 140116 260117 140180
rect 260051 140115 260117 140116
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 255819 29612 255885 29613
rect 255819 29548 255820 29612
rect 255884 29548 255885 29612
rect 255819 29547 255885 29548
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 7174 258134 42618
rect 260054 28253 260114 140115
rect 261234 118894 261854 154338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 273299 270604 273365 270605
rect 273299 270540 273300 270604
rect 273364 270540 273365 270604
rect 273299 270539 273365 270540
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 178000 272414 200898
rect 273302 175949 273362 270539
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 178000 276134 204618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 280291 290052 280357 290053
rect 280291 289988 280292 290052
rect 280356 289988 280357 290052
rect 280291 289987 280357 289988
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 278819 178668 278885 178669
rect 278819 178604 278820 178668
rect 278884 178604 278885 178668
rect 278819 178603 278885 178604
rect 273299 175948 273365 175949
rect 273299 175884 273300 175948
rect 273364 175884 273365 175948
rect 273299 175883 273365 175884
rect 278822 171150 278882 178603
rect 279234 178000 279854 208338
rect 280294 200130 280354 289987
rect 282954 284614 283574 320058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 291147 339556 291213 339557
rect 291147 339492 291148 339556
rect 291212 339492 291213 339556
rect 291147 339491 291213 339492
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 284339 311948 284405 311949
rect 284339 311884 284340 311948
rect 284404 311884 284405 311948
rect 284339 311883 284405 311884
rect 281579 284476 281645 284477
rect 281579 284412 281580 284476
rect 281644 284412 281645 284476
rect 281579 284411 281645 284412
rect 280110 200070 280354 200130
rect 279371 177036 279437 177037
rect 279371 176972 279372 177036
rect 279436 176972 279437 177036
rect 279371 176971 279437 176972
rect 279374 173773 279434 176971
rect 279371 173772 279437 173773
rect 279371 173708 279372 173772
rect 279436 173708 279437 173772
rect 279371 173707 279437 173708
rect 278822 171090 279434 171150
rect 279374 168333 279434 171090
rect 279371 168332 279437 168333
rect 279371 168268 279372 168332
rect 279436 168268 279437 168332
rect 279371 168267 279437 168268
rect 272207 165454 272527 165486
rect 272207 165218 272249 165454
rect 272485 165218 272527 165454
rect 272207 165134 272527 165218
rect 272207 164898 272249 165134
rect 272485 164898 272527 165134
rect 272207 164866 272527 164898
rect 275471 165454 275791 165486
rect 275471 165218 275513 165454
rect 275749 165218 275791 165454
rect 275471 165134 275791 165218
rect 275471 164898 275513 165134
rect 275749 164898 275791 165134
rect 275471 164866 275791 164898
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264099 127124 264165 127125
rect 264099 127060 264100 127124
rect 264164 127060 264165 127124
rect 264099 127059 264165 127060
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 262811 113796 262877 113797
rect 262811 113732 262812 113796
rect 262876 113732 262877 113796
rect 262811 113731 262877 113732
rect 262814 98701 262874 113731
rect 262811 98700 262877 98701
rect 262811 98636 262812 98700
rect 262876 98636 262877 98700
rect 262811 98635 262877 98636
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 264102 59941 264162 127059
rect 264954 122614 265574 158058
rect 270575 147454 270895 147486
rect 270575 147218 270617 147454
rect 270853 147218 270895 147454
rect 270575 147134 270895 147218
rect 270575 146898 270617 147134
rect 270853 146898 270895 147134
rect 270575 146866 270895 146898
rect 273839 147454 274159 147486
rect 273839 147218 273881 147454
rect 274117 147218 274159 147454
rect 273839 147134 274159 147218
rect 273839 146898 273881 147134
rect 274117 146898 274159 147134
rect 273839 146866 274159 146898
rect 277103 147454 277423 147486
rect 277103 147218 277145 147454
rect 277381 147218 277423 147454
rect 277103 147134 277423 147218
rect 277103 146898 277145 147134
rect 277381 146898 277423 147134
rect 277103 146866 277423 146898
rect 280110 142170 280170 200070
rect 280291 195396 280357 195397
rect 280291 195332 280292 195396
rect 280356 195332 280357 195396
rect 280291 195331 280357 195332
rect 280294 151830 280354 195331
rect 281582 157317 281642 284411
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 283787 177444 283853 177445
rect 283787 177380 283788 177444
rect 283852 177380 283853 177444
rect 283787 177379 283853 177380
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 281579 157316 281645 157317
rect 281579 157252 281580 157316
rect 281644 157252 281645 157316
rect 281579 157251 281645 157252
rect 280294 151770 280538 151830
rect 280110 142110 280354 142170
rect 267779 135692 267845 135693
rect 267779 135628 267780 135692
rect 267844 135628 267845 135692
rect 267779 135627 267845 135628
rect 266859 131068 266925 131069
rect 266859 131004 266860 131068
rect 266924 131004 266925 131068
rect 266859 131003 266925 131004
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264099 59940 264165 59941
rect 264099 59876 264100 59940
rect 264164 59876 264165 59940
rect 264099 59875 264165 59876
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 260051 28252 260117 28253
rect 260051 28188 260052 28252
rect 260116 28188 260117 28252
rect 260051 28187 260117 28188
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 50614 265574 86058
rect 266862 54501 266922 131003
rect 267043 100876 267109 100877
rect 267043 100812 267044 100876
rect 267108 100812 267109 100876
rect 267043 100811 267109 100812
rect 267046 86189 267106 100811
rect 267043 86188 267109 86189
rect 267043 86124 267044 86188
rect 267108 86124 267109 86188
rect 267043 86123 267109 86124
rect 267782 58581 267842 135627
rect 280294 131341 280354 142110
rect 280478 135965 280538 151770
rect 282954 140614 283574 176058
rect 283790 143581 283850 177379
rect 283787 143580 283853 143581
rect 283787 143516 283788 143580
rect 283852 143516 283853 143580
rect 283787 143515 283853 143516
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 284342 140453 284402 311883
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 288571 288556 288637 288557
rect 288571 288492 288572 288556
rect 288636 288492 288637 288556
rect 288571 288491 288637 288492
rect 287283 287332 287349 287333
rect 287283 287268 287284 287332
rect 287348 287268 287349 287332
rect 287283 287267 287349 287268
rect 285811 224228 285877 224229
rect 285811 224164 285812 224228
rect 285876 224164 285877 224228
rect 285811 224163 285877 224164
rect 284523 189684 284589 189685
rect 284523 189620 284524 189684
rect 284588 189620 284589 189684
rect 284523 189619 284589 189620
rect 284339 140452 284405 140453
rect 284339 140388 284340 140452
rect 284404 140388 284405 140452
rect 284339 140387 284405 140388
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 280475 135964 280541 135965
rect 280475 135900 280476 135964
rect 280540 135900 280541 135964
rect 280475 135899 280541 135900
rect 280291 131340 280357 131341
rect 280291 131276 280292 131340
rect 280356 131276 280357 131340
rect 280291 131275 280357 131276
rect 272207 129454 272527 129486
rect 272207 129218 272249 129454
rect 272485 129218 272527 129454
rect 272207 129134 272527 129218
rect 272207 128898 272249 129134
rect 272485 128898 272527 129134
rect 272207 128866 272527 128898
rect 275471 129454 275791 129486
rect 275471 129218 275513 129454
rect 275749 129218 275791 129454
rect 275471 129134 275791 129218
rect 275471 128898 275513 129134
rect 275749 128898 275791 129134
rect 275471 128866 275791 128898
rect 270575 111454 270895 111486
rect 270575 111218 270617 111454
rect 270853 111218 270895 111454
rect 270575 111134 270895 111218
rect 270575 110898 270617 111134
rect 270853 110898 270895 111134
rect 270575 110866 270895 110898
rect 273839 111454 274159 111486
rect 273839 111218 273881 111454
rect 274117 111218 274159 111454
rect 273839 111134 274159 111218
rect 273839 110898 273881 111134
rect 274117 110898 274159 111134
rect 273839 110866 274159 110898
rect 277103 111454 277423 111486
rect 277103 111218 277145 111454
rect 277381 111218 277423 111454
rect 277103 111134 277423 111218
rect 277103 110898 277145 111134
rect 277381 110898 277423 111134
rect 277103 110866 277423 110898
rect 282954 104614 283574 140058
rect 284526 116925 284586 189619
rect 285627 181388 285693 181389
rect 285627 181324 285628 181388
rect 285692 181324 285693 181388
rect 285627 181323 285693 181324
rect 284523 116924 284589 116925
rect 284523 116860 284524 116924
rect 284588 116860 284589 116924
rect 284523 116859 284589 116860
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 267963 98020 268029 98021
rect 267963 97956 267964 98020
rect 268028 97956 268029 98020
rect 267963 97955 268029 97956
rect 267779 58580 267845 58581
rect 267779 58516 267780 58580
rect 267844 58516 267845 58580
rect 267779 58515 267845 58516
rect 266859 54500 266925 54501
rect 266859 54436 266860 54500
rect 266924 54436 266925 54500
rect 266859 54435 266925 54436
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 267966 50421 268026 97955
rect 271794 93454 272414 94000
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 264954 50294 265574 50378
rect 267963 50420 268029 50421
rect 267963 50356 267964 50420
rect 268028 50356 268029 50420
rect 267963 50355 268029 50356
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 61174 276134 94000
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 64894 279854 94000
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 285630 3501 285690 181323
rect 285814 106181 285874 224163
rect 287099 193900 287165 193901
rect 287099 193836 287100 193900
rect 287164 193836 287165 193900
rect 287099 193835 287165 193836
rect 285811 106180 285877 106181
rect 285811 106116 285812 106180
rect 285876 106116 285877 106180
rect 285811 106115 285877 106116
rect 287102 3501 287162 193835
rect 287286 102237 287346 287267
rect 288387 202196 288453 202197
rect 288387 202132 288388 202196
rect 288452 202132 288453 202196
rect 288387 202131 288453 202132
rect 287283 102236 287349 102237
rect 287283 102172 287284 102236
rect 287348 102172 287349 102236
rect 287283 102171 287349 102172
rect 288390 3501 288450 202131
rect 288574 106317 288634 288491
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 290595 185604 290661 185605
rect 290595 185540 290596 185604
rect 290660 185540 290661 185604
rect 290595 185539 290661 185540
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 290598 133925 290658 185539
rect 290595 133924 290661 133925
rect 290595 133860 290596 133924
rect 290660 133860 290661 133924
rect 290595 133859 290661 133860
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 288571 106316 288637 106317
rect 288571 106252 288572 106316
rect 288636 106252 288637 106316
rect 288571 106251 288637 106252
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 285627 3500 285693 3501
rect 285627 3436 285628 3500
rect 285692 3436 285693 3500
rect 285627 3435 285693 3436
rect 287099 3500 287165 3501
rect 287099 3436 287100 3500
rect 287164 3436 287165 3500
rect 287099 3435 287165 3436
rect 288387 3500 288453 3501
rect 288387 3436 288388 3500
rect 288452 3436 288453 3500
rect 288387 3435 288453 3436
rect 289794 3454 290414 38898
rect 291150 3501 291210 339491
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 298691 218652 298757 218653
rect 298691 218588 298692 218652
rect 298756 218588 298757 218652
rect 298691 218587 298757 218588
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 293514 186854 294134 186938
rect 295379 186964 295445 186965
rect 295379 186900 295380 186964
rect 295444 186900 295445 186964
rect 295379 186899 295445 186900
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 291331 181524 291397 181525
rect 291331 181460 291332 181524
rect 291396 181460 291397 181524
rect 291331 181459 291397 181460
rect 291334 149157 291394 181459
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 291331 149156 291397 149157
rect 291331 149092 291332 149156
rect 291396 149092 291397 149156
rect 291331 149091 291397 149092
rect 293514 115174 294134 150618
rect 295382 132565 295442 186899
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 295379 132564 295445 132565
rect 295379 132500 295380 132564
rect 295444 132500 295445 132564
rect 295379 132499 295445 132500
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 291147 3500 291213 3501
rect 291147 3436 291148 3500
rect 291212 3436 291213 3500
rect 291147 3435 291213 3436
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 298694 3501 298754 218587
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 298691 3500 298757 3501
rect 298691 3436 298692 3500
rect 298756 3436 298757 3500
rect 298691 3435 298757 3436
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 72721 579218 72957 579454
rect 72721 578898 72957 579134
rect 75686 561218 75922 561454
rect 75686 560898 75922 561134
rect 72721 543218 72957 543454
rect 72721 542898 72957 543134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 78651 579218 78887 579454
rect 78651 578898 78887 579134
rect 84582 579218 84818 579454
rect 84582 578898 84818 579134
rect 81617 561218 81853 561454
rect 81617 560898 81853 561134
rect 78651 543218 78887 543454
rect 78651 542898 78887 543134
rect 84582 543218 84818 543454
rect 84582 542898 84818 543134
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 73020 435218 73256 435454
rect 73020 434898 73256 435134
rect 88380 417218 88616 417454
rect 88380 416898 88616 417134
rect 73020 399218 73256 399454
rect 73020 398898 73256 399134
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73020 291218 73256 291454
rect 73020 290898 73256 291134
rect 73020 255218 73256 255454
rect 73020 254898 73256 255134
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 103740 435218 103976 435454
rect 103740 434898 103976 435134
rect 103740 399218 103976 399454
rect 103740 398898 103976 399134
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 119100 417218 119336 417454
rect 119100 416898 119336 417134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 88380 309218 88616 309454
rect 88380 308898 88616 309134
rect 119100 309218 119336 309454
rect 119100 308898 119336 309134
rect 103740 291218 103976 291454
rect 103740 290898 103976 291134
rect 88380 273218 88616 273454
rect 88380 272898 88616 273134
rect 119100 273218 119336 273454
rect 119100 272898 119336 273134
rect 103740 255218 103976 255454
rect 103740 254898 103976 255134
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 134460 291218 134696 291454
rect 134460 290898 134696 291134
rect 134460 255218 134696 255454
rect 134460 254898 134696 255134
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 149820 309218 150056 309454
rect 149820 308898 150056 309134
rect 149820 273218 150056 273454
rect 149820 272898 150056 273134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 69128 165218 69364 165454
rect 69128 164898 69364 165134
rect 164192 165218 164428 165454
rect 164192 164898 164428 165134
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 69128 129218 69364 129454
rect 69128 128898 69364 129134
rect 164192 129218 164428 129454
rect 164192 128898 164428 129134
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 204450 255218 204686 255454
rect 204450 254898 204686 255134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 219810 273218 220046 273454
rect 219810 272898 220046 273134
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 221249 165218 221485 165454
rect 221249 164898 221485 165134
rect 224513 165218 224749 165454
rect 224513 164898 224749 165134
rect 219617 147218 219853 147454
rect 219617 146898 219853 147134
rect 222881 147218 223117 147454
rect 222881 146898 223117 147134
rect 226145 147218 226381 147454
rect 226145 146898 226381 147134
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 235170 255218 235406 255454
rect 235170 254898 235406 255134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 221249 129218 221485 129454
rect 221249 128898 221485 129134
rect 224513 129218 224749 129454
rect 224513 128898 224749 129134
rect 219617 111218 219853 111454
rect 219617 110898 219853 111134
rect 222881 111218 223117 111454
rect 222881 110898 223117 111134
rect 226145 111218 226381 111454
rect 226145 110898 226381 111134
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 272249 165218 272485 165454
rect 272249 164898 272485 165134
rect 275513 165218 275749 165454
rect 275513 164898 275749 165134
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 270617 147218 270853 147454
rect 270617 146898 270853 147134
rect 273881 147218 274117 147454
rect 273881 146898 274117 147134
rect 277145 147218 277381 147454
rect 277145 146898 277381 147134
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 272249 129218 272485 129454
rect 272249 128898 272485 129134
rect 275513 129218 275749 129454
rect 275513 128898 275749 129134
rect 270617 111218 270853 111454
rect 270617 110898 270853 111134
rect 273881 111218 274117 111454
rect 273881 110898 274117 111134
rect 277145 111218 277381 111454
rect 277145 110898 277381 111134
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 72721 579454
rect 72957 579218 78651 579454
rect 78887 579218 84582 579454
rect 84818 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 72721 579134
rect 72957 578898 78651 579134
rect 78887 578898 84582 579134
rect 84818 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 75686 561454
rect 75922 561218 81617 561454
rect 81853 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 75686 561134
rect 75922 560898 81617 561134
rect 81853 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 72721 543454
rect 72957 543218 78651 543454
rect 78887 543218 84582 543454
rect 84818 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 72721 543134
rect 72957 542898 78651 543134
rect 78887 542898 84582 543134
rect 84818 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73020 435454
rect 73256 435218 103740 435454
rect 103976 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73020 435134
rect 73256 434898 103740 435134
rect 103976 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 88380 417454
rect 88616 417218 119100 417454
rect 119336 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 88380 417134
rect 88616 416898 119100 417134
rect 119336 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73020 399454
rect 73256 399218 103740 399454
rect 103976 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73020 399134
rect 73256 398898 103740 399134
rect 103976 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 88380 309454
rect 88616 309218 119100 309454
rect 119336 309218 149820 309454
rect 150056 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 88380 309134
rect 88616 308898 119100 309134
rect 119336 308898 149820 309134
rect 150056 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73020 291454
rect 73256 291218 103740 291454
rect 103976 291218 134460 291454
rect 134696 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73020 291134
rect 73256 290898 103740 291134
rect 103976 290898 134460 291134
rect 134696 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 88380 273454
rect 88616 273218 119100 273454
rect 119336 273218 149820 273454
rect 150056 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 219810 273454
rect 220046 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 88380 273134
rect 88616 272898 119100 273134
rect 119336 272898 149820 273134
rect 150056 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 219810 273134
rect 220046 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73020 255454
rect 73256 255218 103740 255454
rect 103976 255218 134460 255454
rect 134696 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 204450 255454
rect 204686 255218 235170 255454
rect 235406 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73020 255134
rect 73256 254898 103740 255134
rect 103976 254898 134460 255134
rect 134696 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 204450 255134
rect 204686 254898 235170 255134
rect 235406 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 69128 165454
rect 69364 165218 164192 165454
rect 164428 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 221249 165454
rect 221485 165218 224513 165454
rect 224749 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 272249 165454
rect 272485 165218 275513 165454
rect 275749 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 69128 165134
rect 69364 164898 164192 165134
rect 164428 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 221249 165134
rect 221485 164898 224513 165134
rect 224749 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 272249 165134
rect 272485 164898 275513 165134
rect 275749 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 219617 147454
rect 219853 147218 222881 147454
rect 223117 147218 226145 147454
rect 226381 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 270617 147454
rect 270853 147218 273881 147454
rect 274117 147218 277145 147454
rect 277381 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 219617 147134
rect 219853 146898 222881 147134
rect 223117 146898 226145 147134
rect 226381 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 270617 147134
rect 270853 146898 273881 147134
rect 274117 146898 277145 147134
rect 277381 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 69128 129454
rect 69364 129218 164192 129454
rect 164428 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 221249 129454
rect 221485 129218 224513 129454
rect 224749 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 272249 129454
rect 272485 129218 275513 129454
rect 275749 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 69128 129134
rect 69364 128898 164192 129134
rect 164428 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 221249 129134
rect 221485 128898 224513 129134
rect 224749 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 272249 129134
rect 272485 128898 275513 129134
rect 275749 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 219617 111454
rect 219853 111218 222881 111454
rect 223117 111218 226145 111454
rect 226381 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 270617 111454
rect 270853 111218 273881 111454
rect 274117 111218 277145 111454
rect 277381 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 219617 111134
rect 219853 110898 222881 111134
rect 223117 110898 226145 111134
rect 226381 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 270617 111134
rect 270853 110898 273881 111134
rect 274117 110898 277145 111134
rect 277381 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use wrapped_spell  wrapped_spell_1
timestamp 1640263499
transform 1 0 68770 0 1 241592
box 0 0 86000 86000
use wrapped_ppm_decoder  wrapped_ppm_decoder_3
timestamp 1640263499
transform 1 0 68770 0 1 539166
box 0 0 20000 50000
use wrapped_ppm_coder  wrapped_ppm_coder_2
timestamp 1640263499
transform 1 0 68770 0 1 390356
box 0 0 51907 54051
use wrapped_function_generator  wrapped_function_generator_0
timestamp 1640263499
transform 1 0 200200 0 1 240182
box 0 0 44000 44000
use wb_openram_wrapper  wb_openram_wrapper
timestamp 1640263499
transform 1 0 217000 0 1 96000
box 0 144 12000 79688
use wb_bridge_2way  wb_bridge_2way
timestamp 1640263499
transform 1 0 268000 0 1 96000
box 0 0 12000 79688
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 1640263499
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 94000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 178000 218414 238182 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 176600 74414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 176600 110414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 176600 146414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 329592 74414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 329592 110414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 446407 74414 537166 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 591166 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 446407 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 329592 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 286182 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 94000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 178000 222134 238182 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 176600 78134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 176600 114134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 176600 150134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 329592 78134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 329592 114134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 446407 78134 537166 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 591166 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 446407 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 329592 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 286182 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 94000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 178000 225854 238182 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 176600 81854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 176600 117854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 176600 153854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 329592 81854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 329592 117854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 446407 81854 537166 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 591166 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 446407 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 329592 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 286182 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 94000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 178000 229574 238182 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 176600 85574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 176600 121574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 329592 85574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 329592 121574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 446407 85574 537166 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 591166 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 446407 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 176600 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 286182 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 238182 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 238182 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 176600 99854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 176600 135854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 329592 99854 388356 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 446407 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 329592 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 286182 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 286182 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 178000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 238182 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 176600 67574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 176600 103574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 176600 139574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 329592 67574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 329592 103574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 446407 67574 537166 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 591166 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 446407 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 329592 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 286182 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 238182 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 238182 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 176600 92414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 176600 128414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 329592 92414 388356 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 446407 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 329592 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 176600 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 286182 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 286182 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 178000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 238182 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 238182 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 176600 96134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 176600 132134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 329592 96134 388356 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 446407 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 329592 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 286182 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 286182 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 178000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
