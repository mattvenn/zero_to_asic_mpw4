* NGSPICE file created from user_project_wrapper.ext - technology: sky130A

* Black-box entry subcircuit for wrapped_keyvalue abstract view
.subckt wrapped_keyvalue active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la1_data_in[0] la1_data_in[10] la1_data_in[11] la1_data_in[12] la1_data_in[13] la1_data_in[14]
+ la1_data_in[15] la1_data_in[16] la1_data_in[17] la1_data_in[18] la1_data_in[19]
+ la1_data_in[1] la1_data_in[20] la1_data_in[21] la1_data_in[22] la1_data_in[23] la1_data_in[24]
+ la1_data_in[25] la1_data_in[26] la1_data_in[27] la1_data_in[28] la1_data_in[29]
+ la1_data_in[2] la1_data_in[30] la1_data_in[31] la1_data_in[3] la1_data_in[4] la1_data_in[5]
+ la1_data_in[6] la1_data_in[7] la1_data_in[8] la1_data_in[9] la1_data_out[0] la1_data_out[10]
+ la1_data_out[11] la1_data_out[12] la1_data_out[13] la1_data_out[14] la1_data_out[15]
+ la1_data_out[16] la1_data_out[17] la1_data_out[18] la1_data_out[19] la1_data_out[1]
+ la1_data_out[20] la1_data_out[21] la1_data_out[22] la1_data_out[23] la1_data_out[24]
+ la1_data_out[25] la1_data_out[26] la1_data_out[27] la1_data_out[28] la1_data_out[29]
+ la1_data_out[2] la1_data_out[30] la1_data_out[31] la1_data_out[3] la1_data_out[4]
+ la1_data_out[5] la1_data_out[6] la1_data_out[7] la1_data_out[8] la1_data_out[9]
+ la1_oenb[0] la1_oenb[10] la1_oenb[11] la1_oenb[12] la1_oenb[13] la1_oenb[14] la1_oenb[15]
+ la1_oenb[16] la1_oenb[17] la1_oenb[18] la1_oenb[19] la1_oenb[1] la1_oenb[20] la1_oenb[21]
+ la1_oenb[22] la1_oenb[23] la1_oenb[24] la1_oenb[25] la1_oenb[26] la1_oenb[27] la1_oenb[28]
+ la1_oenb[29] la1_oenb[2] la1_oenb[30] la1_oenb[31] la1_oenb[3] la1_oenb[4] la1_oenb[5]
+ la1_oenb[6] la1_oenb[7] la1_oenb[8] la1_oenb[9] vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o
+ wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
.ends

* Black-box entry subcircuit for wrapped_ppm_coder abstract view
.subckt wrapped_ppm_coder active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] vccd1 vssd1 wb_clk_i
.ends

* Black-box entry subcircuit for wrapped_silife abstract view
.subckt wrapped_silife active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la1_data_in[0] la1_data_in[10] la1_data_in[11] la1_data_in[12] la1_data_in[13] la1_data_in[14]
+ la1_data_in[15] la1_data_in[16] la1_data_in[17] la1_data_in[18] la1_data_in[19]
+ la1_data_in[1] la1_data_in[20] la1_data_in[21] la1_data_in[22] la1_data_in[23] la1_data_in[24]
+ la1_data_in[25] la1_data_in[26] la1_data_in[27] la1_data_in[28] la1_data_in[29]
+ la1_data_in[2] la1_data_in[30] la1_data_in[31] la1_data_in[3] la1_data_in[4] la1_data_in[5]
+ la1_data_in[6] la1_data_in[7] la1_data_in[8] la1_data_in[9] la1_data_out[0] la1_data_out[10]
+ la1_data_out[11] la1_data_out[12] la1_data_out[13] la1_data_out[14] la1_data_out[15]
+ la1_data_out[16] la1_data_out[17] la1_data_out[18] la1_data_out[19] la1_data_out[1]
+ la1_data_out[20] la1_data_out[21] la1_data_out[22] la1_data_out[23] la1_data_out[24]
+ la1_data_out[25] la1_data_out[26] la1_data_out[27] la1_data_out[28] la1_data_out[29]
+ la1_data_out[2] la1_data_out[30] la1_data_out[31] la1_data_out[3] la1_data_out[4]
+ la1_data_out[5] la1_data_out[6] la1_data_out[7] la1_data_out[8] la1_data_out[9]
+ la1_oenb[0] la1_oenb[10] la1_oenb[11] la1_oenb[12] la1_oenb[13] la1_oenb[14] la1_oenb[15]
+ la1_oenb[16] la1_oenb[17] la1_oenb[18] la1_oenb[19] la1_oenb[1] la1_oenb[20] la1_oenb[21]
+ la1_oenb[22] la1_oenb[23] la1_oenb[24] la1_oenb[25] la1_oenb[26] la1_oenb[27] la1_oenb[28]
+ la1_oenb[29] la1_oenb[2] la1_oenb[30] la1_oenb[31] la1_oenb[3] la1_oenb[4] la1_oenb[5]
+ la1_oenb[6] la1_oenb[7] la1_oenb[8] la1_oenb[9] vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o
+ wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14]
+ wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1]
+ wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25]
+ wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30]
+ wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8]
+ wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13]
+ wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19]
+ wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24]
+ wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2]
+ wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6]
+ wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11]
+ wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17]
+ wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22]
+ wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28]
+ wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4]
+ wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1]
+ wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
.ends

* Black-box entry subcircuit for wrapped_spraid abstract view
.subckt wrapped_spraid active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
.ends

* Black-box entry subcircuit for wb_bridge_2way abstract view
.subckt wb_bridge_2way vccd1 vssd1 wb_clk_i wb_rst_i wbm_a_ack_i wbm_a_adr_o[0] wbm_a_adr_o[10]
+ wbm_a_adr_o[11] wbm_a_adr_o[12] wbm_a_adr_o[13] wbm_a_adr_o[14] wbm_a_adr_o[15]
+ wbm_a_adr_o[16] wbm_a_adr_o[17] wbm_a_adr_o[18] wbm_a_adr_o[19] wbm_a_adr_o[1] wbm_a_adr_o[20]
+ wbm_a_adr_o[21] wbm_a_adr_o[22] wbm_a_adr_o[23] wbm_a_adr_o[24] wbm_a_adr_o[25]
+ wbm_a_adr_o[26] wbm_a_adr_o[27] wbm_a_adr_o[28] wbm_a_adr_o[29] wbm_a_adr_o[2] wbm_a_adr_o[30]
+ wbm_a_adr_o[31] wbm_a_adr_o[3] wbm_a_adr_o[4] wbm_a_adr_o[5] wbm_a_adr_o[6] wbm_a_adr_o[7]
+ wbm_a_adr_o[8] wbm_a_adr_o[9] wbm_a_cyc_o wbm_a_dat_i[0] wbm_a_dat_i[10] wbm_a_dat_i[11]
+ wbm_a_dat_i[12] wbm_a_dat_i[13] wbm_a_dat_i[14] wbm_a_dat_i[15] wbm_a_dat_i[16]
+ wbm_a_dat_i[17] wbm_a_dat_i[18] wbm_a_dat_i[19] wbm_a_dat_i[1] wbm_a_dat_i[20] wbm_a_dat_i[21]
+ wbm_a_dat_i[22] wbm_a_dat_i[23] wbm_a_dat_i[24] wbm_a_dat_i[25] wbm_a_dat_i[26]
+ wbm_a_dat_i[27] wbm_a_dat_i[28] wbm_a_dat_i[29] wbm_a_dat_i[2] wbm_a_dat_i[30] wbm_a_dat_i[31]
+ wbm_a_dat_i[3] wbm_a_dat_i[4] wbm_a_dat_i[5] wbm_a_dat_i[6] wbm_a_dat_i[7] wbm_a_dat_i[8]
+ wbm_a_dat_i[9] wbm_a_dat_o[0] wbm_a_dat_o[10] wbm_a_dat_o[11] wbm_a_dat_o[12] wbm_a_dat_o[13]
+ wbm_a_dat_o[14] wbm_a_dat_o[15] wbm_a_dat_o[16] wbm_a_dat_o[17] wbm_a_dat_o[18]
+ wbm_a_dat_o[19] wbm_a_dat_o[1] wbm_a_dat_o[20] wbm_a_dat_o[21] wbm_a_dat_o[22] wbm_a_dat_o[23]
+ wbm_a_dat_o[24] wbm_a_dat_o[25] wbm_a_dat_o[26] wbm_a_dat_o[27] wbm_a_dat_o[28]
+ wbm_a_dat_o[29] wbm_a_dat_o[2] wbm_a_dat_o[30] wbm_a_dat_o[31] wbm_a_dat_o[3] wbm_a_dat_o[4]
+ wbm_a_dat_o[5] wbm_a_dat_o[6] wbm_a_dat_o[7] wbm_a_dat_o[8] wbm_a_dat_o[9] wbm_a_sel_o[0]
+ wbm_a_sel_o[1] wbm_a_sel_o[2] wbm_a_sel_o[3] wbm_a_stb_o wbm_a_we_o wbm_b_ack_i
+ wbm_b_adr_o[0] wbm_b_adr_o[1] wbm_b_adr_o[2] wbm_b_adr_o[3] wbm_b_adr_o[4] wbm_b_adr_o[5]
+ wbm_b_adr_o[6] wbm_b_adr_o[7] wbm_b_adr_o[8] wbm_b_adr_o[9] wbm_b_cyc_o wbm_b_dat_i[0]
+ wbm_b_dat_i[10] wbm_b_dat_i[11] wbm_b_dat_i[12] wbm_b_dat_i[13] wbm_b_dat_i[14]
+ wbm_b_dat_i[15] wbm_b_dat_i[16] wbm_b_dat_i[17] wbm_b_dat_i[18] wbm_b_dat_i[19]
+ wbm_b_dat_i[1] wbm_b_dat_i[20] wbm_b_dat_i[21] wbm_b_dat_i[22] wbm_b_dat_i[23] wbm_b_dat_i[24]
+ wbm_b_dat_i[25] wbm_b_dat_i[26] wbm_b_dat_i[27] wbm_b_dat_i[28] wbm_b_dat_i[29]
+ wbm_b_dat_i[2] wbm_b_dat_i[30] wbm_b_dat_i[31] wbm_b_dat_i[3] wbm_b_dat_i[4] wbm_b_dat_i[5]
+ wbm_b_dat_i[6] wbm_b_dat_i[7] wbm_b_dat_i[8] wbm_b_dat_i[9] wbm_b_dat_o[0] wbm_b_dat_o[10]
+ wbm_b_dat_o[11] wbm_b_dat_o[12] wbm_b_dat_o[13] wbm_b_dat_o[14] wbm_b_dat_o[15]
+ wbm_b_dat_o[16] wbm_b_dat_o[17] wbm_b_dat_o[18] wbm_b_dat_o[19] wbm_b_dat_o[1] wbm_b_dat_o[20]
+ wbm_b_dat_o[21] wbm_b_dat_o[22] wbm_b_dat_o[23] wbm_b_dat_o[24] wbm_b_dat_o[25]
+ wbm_b_dat_o[26] wbm_b_dat_o[27] wbm_b_dat_o[28] wbm_b_dat_o[29] wbm_b_dat_o[2] wbm_b_dat_o[30]
+ wbm_b_dat_o[31] wbm_b_dat_o[3] wbm_b_dat_o[4] wbm_b_dat_o[5] wbm_b_dat_o[6] wbm_b_dat_o[7]
+ wbm_b_dat_o[8] wbm_b_dat_o[9] wbm_b_sel_o[0] wbm_b_sel_o[1] wbm_b_sel_o[2] wbm_b_sel_o[3]
+ wbm_b_stb_o wbm_b_we_o wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
.ends

* Black-box entry subcircuit for sky130_sram_1kbyte_1rw1r_32x256_8 abstract view
.subckt sky130_sram_1kbyte_1rw1r_32x256_8 din0[0] din0[1] din0[2] din0[3] din0[4]
+ din0[5] din0[6] din0[7] din0[8] din0[9] din0[10] din0[11] din0[12] din0[13] din0[14]
+ din0[15] din0[16] din0[17] din0[18] din0[19] din0[20] din0[21] din0[22] din0[23]
+ din0[24] din0[25] din0[26] din0[27] din0[28] din0[29] din0[30] din0[31] addr0[0]
+ addr0[1] addr0[2] addr0[3] addr0[4] addr0[5] addr0[6] addr0[7] addr1[0] addr1[1]
+ addr1[2] addr1[3] addr1[4] addr1[5] addr1[6] addr1[7] csb0 csb1 web0 clk0 clk1 wmask0[0]
+ wmask0[1] wmask0[2] wmask0[3] dout0[0] dout0[1] dout0[2] dout0[3] dout0[4] dout0[5]
+ dout0[6] dout0[7] dout0[8] dout0[9] dout0[10] dout0[11] dout0[12] dout0[13] dout0[14]
+ dout0[15] dout0[16] dout0[17] dout0[18] dout0[19] dout0[20] dout0[21] dout0[22]
+ dout0[23] dout0[24] dout0[25] dout0[26] dout0[27] dout0[28] dout0[29] dout0[30]
+ dout0[31] dout1[0] dout1[1] dout1[2] dout1[3] dout1[4] dout1[5] dout1[6] dout1[7]
+ dout1[8] dout1[9] dout1[10] dout1[11] dout1[12] dout1[13] dout1[14] dout1[15] dout1[16]
+ dout1[17] dout1[18] dout1[19] dout1[20] dout1[21] dout1[22] dout1[23] dout1[24]
+ dout1[25] dout1[26] dout1[27] dout1[28] dout1[29] dout1[30] dout1[31] vccd1 vssd1
.ends

* Black-box entry subcircuit for wrapped_skullfet abstract view
.subckt wrapped_skullfet active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la1_data_in[0] la1_data_in[10] la1_data_in[11] la1_data_in[12] la1_data_in[13] la1_data_in[14]
+ la1_data_in[15] la1_data_in[16] la1_data_in[17] la1_data_in[18] la1_data_in[19]
+ la1_data_in[1] la1_data_in[20] la1_data_in[21] la1_data_in[22] la1_data_in[23] la1_data_in[24]
+ la1_data_in[25] la1_data_in[26] la1_data_in[27] la1_data_in[28] la1_data_in[29]
+ la1_data_in[2] la1_data_in[30] la1_data_in[31] la1_data_in[3] la1_data_in[4] la1_data_in[5]
+ la1_data_in[6] la1_data_in[7] la1_data_in[8] la1_data_in[9] la1_data_out[0] la1_data_out[10]
+ la1_data_out[11] la1_data_out[12] la1_data_out[13] la1_data_out[14] la1_data_out[15]
+ la1_data_out[16] la1_data_out[17] la1_data_out[18] la1_data_out[19] la1_data_out[1]
+ la1_data_out[20] la1_data_out[21] la1_data_out[22] la1_data_out[23] la1_data_out[24]
+ la1_data_out[25] la1_data_out[26] la1_data_out[27] la1_data_out[28] la1_data_out[29]
+ la1_data_out[2] la1_data_out[30] la1_data_out[31] la1_data_out[3] la1_data_out[4]
+ la1_data_out[5] la1_data_out[6] la1_data_out[7] la1_data_out[8] la1_data_out[9]
+ la1_oenb[0] la1_oenb[10] la1_oenb[11] la1_oenb[12] la1_oenb[13] la1_oenb[14] la1_oenb[15]
+ la1_oenb[16] la1_oenb[17] la1_oenb[18] la1_oenb[19] la1_oenb[1] la1_oenb[20] la1_oenb[21]
+ la1_oenb[22] la1_oenb[23] la1_oenb[24] la1_oenb[25] la1_oenb[26] la1_oenb[27] la1_oenb[28]
+ la1_oenb[29] la1_oenb[2] la1_oenb[30] la1_oenb[31] la1_oenb[3] la1_oenb[4] la1_oenb[5]
+ la1_oenb[6] la1_oenb[7] la1_oenb[8] la1_oenb[9] vccd1 vssd1 wb_clk_i
.ends

* Black-box entry subcircuit for wb_openram_wrapper abstract view
.subckt wb_openram_wrapper ram_addr0[0] ram_addr0[1] ram_addr0[2] ram_addr0[3] ram_addr0[4]
+ ram_addr0[5] ram_addr0[6] ram_addr0[7] ram_addr1[0] ram_addr1[1] ram_addr1[2] ram_addr1[3]
+ ram_addr1[4] ram_addr1[5] ram_addr1[6] ram_addr1[7] ram_clk0 ram_clk1 ram_csb0 ram_csb1
+ ram_din0[0] ram_din0[10] ram_din0[11] ram_din0[12] ram_din0[13] ram_din0[14] ram_din0[15]
+ ram_din0[16] ram_din0[17] ram_din0[18] ram_din0[19] ram_din0[1] ram_din0[20] ram_din0[21]
+ ram_din0[22] ram_din0[23] ram_din0[24] ram_din0[25] ram_din0[26] ram_din0[27] ram_din0[28]
+ ram_din0[29] ram_din0[2] ram_din0[30] ram_din0[31] ram_din0[3] ram_din0[4] ram_din0[5]
+ ram_din0[6] ram_din0[7] ram_din0[8] ram_din0[9] ram_dout0[0] ram_dout0[10] ram_dout0[11]
+ ram_dout0[12] ram_dout0[13] ram_dout0[14] ram_dout0[15] ram_dout0[16] ram_dout0[17]
+ ram_dout0[18] ram_dout0[19] ram_dout0[1] ram_dout0[20] ram_dout0[21] ram_dout0[22]
+ ram_dout0[23] ram_dout0[24] ram_dout0[25] ram_dout0[26] ram_dout0[27] ram_dout0[28]
+ ram_dout0[29] ram_dout0[2] ram_dout0[30] ram_dout0[31] ram_dout0[3] ram_dout0[4]
+ ram_dout0[5] ram_dout0[6] ram_dout0[7] ram_dout0[8] ram_dout0[9] ram_dout1[0] ram_dout1[10]
+ ram_dout1[11] ram_dout1[12] ram_dout1[13] ram_dout1[14] ram_dout1[15] ram_dout1[16]
+ ram_dout1[17] ram_dout1[18] ram_dout1[19] ram_dout1[1] ram_dout1[20] ram_dout1[21]
+ ram_dout1[22] ram_dout1[23] ram_dout1[24] ram_dout1[25] ram_dout1[26] ram_dout1[27]
+ ram_dout1[28] ram_dout1[29] ram_dout1[2] ram_dout1[30] ram_dout1[31] ram_dout1[3]
+ ram_dout1[4] ram_dout1[5] ram_dout1[6] ram_dout1[7] ram_dout1[8] ram_dout1[9] ram_web0
+ ram_wmask0[0] ram_wmask0[1] ram_wmask0[2] ram_wmask0[3] vccd1 vssd1 wb_a_clk_i wb_a_rst_i
+ wb_b_clk_i wb_b_rst_i wbs_a_ack_o wbs_a_adr_i[0] wbs_a_adr_i[1] wbs_a_adr_i[2] wbs_a_adr_i[3]
+ wbs_a_adr_i[4] wbs_a_adr_i[5] wbs_a_adr_i[6] wbs_a_adr_i[7] wbs_a_adr_i[8] wbs_a_adr_i[9]
+ wbs_a_cyc_i wbs_a_dat_i[0] wbs_a_dat_i[10] wbs_a_dat_i[11] wbs_a_dat_i[12] wbs_a_dat_i[13]
+ wbs_a_dat_i[14] wbs_a_dat_i[15] wbs_a_dat_i[16] wbs_a_dat_i[17] wbs_a_dat_i[18]
+ wbs_a_dat_i[19] wbs_a_dat_i[1] wbs_a_dat_i[20] wbs_a_dat_i[21] wbs_a_dat_i[22] wbs_a_dat_i[23]
+ wbs_a_dat_i[24] wbs_a_dat_i[25] wbs_a_dat_i[26] wbs_a_dat_i[27] wbs_a_dat_i[28]
+ wbs_a_dat_i[29] wbs_a_dat_i[2] wbs_a_dat_i[30] wbs_a_dat_i[31] wbs_a_dat_i[3] wbs_a_dat_i[4]
+ wbs_a_dat_i[5] wbs_a_dat_i[6] wbs_a_dat_i[7] wbs_a_dat_i[8] wbs_a_dat_i[9] wbs_a_dat_o[0]
+ wbs_a_dat_o[10] wbs_a_dat_o[11] wbs_a_dat_o[12] wbs_a_dat_o[13] wbs_a_dat_o[14]
+ wbs_a_dat_o[15] wbs_a_dat_o[16] wbs_a_dat_o[17] wbs_a_dat_o[18] wbs_a_dat_o[19]
+ wbs_a_dat_o[1] wbs_a_dat_o[20] wbs_a_dat_o[21] wbs_a_dat_o[22] wbs_a_dat_o[23] wbs_a_dat_o[24]
+ wbs_a_dat_o[25] wbs_a_dat_o[26] wbs_a_dat_o[27] wbs_a_dat_o[28] wbs_a_dat_o[29]
+ wbs_a_dat_o[2] wbs_a_dat_o[30] wbs_a_dat_o[31] wbs_a_dat_o[3] wbs_a_dat_o[4] wbs_a_dat_o[5]
+ wbs_a_dat_o[6] wbs_a_dat_o[7] wbs_a_dat_o[8] wbs_a_dat_o[9] wbs_a_sel_i[0] wbs_a_sel_i[1]
+ wbs_a_sel_i[2] wbs_a_sel_i[3] wbs_a_stb_i wbs_a_we_i wbs_b_ack_o wbs_b_adr_i[0]
+ wbs_b_adr_i[1] wbs_b_adr_i[2] wbs_b_adr_i[3] wbs_b_adr_i[4] wbs_b_adr_i[5] wbs_b_adr_i[6]
+ wbs_b_adr_i[7] wbs_b_adr_i[8] wbs_b_adr_i[9] wbs_b_cyc_i wbs_b_dat_i[0] wbs_b_dat_i[10]
+ wbs_b_dat_i[11] wbs_b_dat_i[12] wbs_b_dat_i[13] wbs_b_dat_i[14] wbs_b_dat_i[15]
+ wbs_b_dat_i[16] wbs_b_dat_i[17] wbs_b_dat_i[18] wbs_b_dat_i[19] wbs_b_dat_i[1] wbs_b_dat_i[20]
+ wbs_b_dat_i[21] wbs_b_dat_i[22] wbs_b_dat_i[23] wbs_b_dat_i[24] wbs_b_dat_i[25]
+ wbs_b_dat_i[26] wbs_b_dat_i[27] wbs_b_dat_i[28] wbs_b_dat_i[29] wbs_b_dat_i[2] wbs_b_dat_i[30]
+ wbs_b_dat_i[31] wbs_b_dat_i[3] wbs_b_dat_i[4] wbs_b_dat_i[5] wbs_b_dat_i[6] wbs_b_dat_i[7]
+ wbs_b_dat_i[8] wbs_b_dat_i[9] wbs_b_dat_o[0] wbs_b_dat_o[10] wbs_b_dat_o[11] wbs_b_dat_o[12]
+ wbs_b_dat_o[13] wbs_b_dat_o[14] wbs_b_dat_o[15] wbs_b_dat_o[16] wbs_b_dat_o[17]
+ wbs_b_dat_o[18] wbs_b_dat_o[19] wbs_b_dat_o[1] wbs_b_dat_o[20] wbs_b_dat_o[21] wbs_b_dat_o[22]
+ wbs_b_dat_o[23] wbs_b_dat_o[24] wbs_b_dat_o[25] wbs_b_dat_o[26] wbs_b_dat_o[27]
+ wbs_b_dat_o[28] wbs_b_dat_o[29] wbs_b_dat_o[2] wbs_b_dat_o[30] wbs_b_dat_o[31] wbs_b_dat_o[3]
+ wbs_b_dat_o[4] wbs_b_dat_o[5] wbs_b_dat_o[6] wbs_b_dat_o[7] wbs_b_dat_o[8] wbs_b_dat_o[9]
+ wbs_b_sel_i[0] wbs_b_sel_i[1] wbs_b_sel_i[2] wbs_b_sel_i[3] wbs_b_stb_i wbs_b_we_i
+ writable_port_req
.ends

* Black-box entry subcircuit for wrapped_ppm_decoder abstract view
.subckt wrapped_ppm_decoder active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] vccd1 vssd1 wb_clk_i
.ends

* Black-box entry subcircuit for wrapped_function_generator abstract view
.subckt wrapped_function_generator active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] rambus_wb_ack_i rambus_wb_adr_o[0] rambus_wb_adr_o[1] rambus_wb_adr_o[2]
+ rambus_wb_adr_o[3] rambus_wb_adr_o[4] rambus_wb_adr_o[5] rambus_wb_adr_o[6] rambus_wb_adr_o[7]
+ rambus_wb_adr_o[8] rambus_wb_adr_o[9] rambus_wb_clk_o rambus_wb_cyc_o rambus_wb_dat_i[0]
+ rambus_wb_dat_i[10] rambus_wb_dat_i[11] rambus_wb_dat_i[12] rambus_wb_dat_i[13]
+ rambus_wb_dat_i[14] rambus_wb_dat_i[15] rambus_wb_dat_i[16] rambus_wb_dat_i[17]
+ rambus_wb_dat_i[18] rambus_wb_dat_i[19] rambus_wb_dat_i[1] rambus_wb_dat_i[20] rambus_wb_dat_i[21]
+ rambus_wb_dat_i[22] rambus_wb_dat_i[23] rambus_wb_dat_i[24] rambus_wb_dat_i[25]
+ rambus_wb_dat_i[26] rambus_wb_dat_i[27] rambus_wb_dat_i[28] rambus_wb_dat_i[29]
+ rambus_wb_dat_i[2] rambus_wb_dat_i[30] rambus_wb_dat_i[31] rambus_wb_dat_i[3] rambus_wb_dat_i[4]
+ rambus_wb_dat_i[5] rambus_wb_dat_i[6] rambus_wb_dat_i[7] rambus_wb_dat_i[8] rambus_wb_dat_i[9]
+ rambus_wb_dat_o[0] rambus_wb_dat_o[10] rambus_wb_dat_o[11] rambus_wb_dat_o[12] rambus_wb_dat_o[13]
+ rambus_wb_dat_o[14] rambus_wb_dat_o[15] rambus_wb_dat_o[16] rambus_wb_dat_o[17]
+ rambus_wb_dat_o[18] rambus_wb_dat_o[19] rambus_wb_dat_o[1] rambus_wb_dat_o[20] rambus_wb_dat_o[21]
+ rambus_wb_dat_o[22] rambus_wb_dat_o[23] rambus_wb_dat_o[24] rambus_wb_dat_o[25]
+ rambus_wb_dat_o[26] rambus_wb_dat_o[27] rambus_wb_dat_o[28] rambus_wb_dat_o[29]
+ rambus_wb_dat_o[2] rambus_wb_dat_o[30] rambus_wb_dat_o[31] rambus_wb_dat_o[3] rambus_wb_dat_o[4]
+ rambus_wb_dat_o[5] rambus_wb_dat_o[6] rambus_wb_dat_o[7] rambus_wb_dat_o[8] rambus_wb_dat_o[9]
+ rambus_wb_rst_o rambus_wb_sel_o[0] rambus_wb_sel_o[1] rambus_wb_sel_o[2] rambus_wb_sel_o[3]
+ rambus_wb_stb_o rambus_wb_we_o vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
.ends

* Black-box entry subcircuit for wrapped_spell abstract view
.subckt wrapped_spell active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la1_data_in[0] la1_data_in[10] la1_data_in[11] la1_data_in[12] la1_data_in[13] la1_data_in[14]
+ la1_data_in[15] la1_data_in[16] la1_data_in[17] la1_data_in[18] la1_data_in[19]
+ la1_data_in[1] la1_data_in[20] la1_data_in[21] la1_data_in[22] la1_data_in[23] la1_data_in[24]
+ la1_data_in[25] la1_data_in[26] la1_data_in[27] la1_data_in[28] la1_data_in[29]
+ la1_data_in[2] la1_data_in[30] la1_data_in[31] la1_data_in[3] la1_data_in[4] la1_data_in[5]
+ la1_data_in[6] la1_data_in[7] la1_data_in[8] la1_data_in[9] la1_data_out[0] la1_data_out[10]
+ la1_data_out[11] la1_data_out[12] la1_data_out[13] la1_data_out[14] la1_data_out[15]
+ la1_data_out[16] la1_data_out[17] la1_data_out[18] la1_data_out[19] la1_data_out[1]
+ la1_data_out[20] la1_data_out[21] la1_data_out[22] la1_data_out[23] la1_data_out[24]
+ la1_data_out[25] la1_data_out[26] la1_data_out[27] la1_data_out[28] la1_data_out[29]
+ la1_data_out[2] la1_data_out[30] la1_data_out[31] la1_data_out[3] la1_data_out[4]
+ la1_data_out[5] la1_data_out[6] la1_data_out[7] la1_data_out[8] la1_data_out[9]
+ la1_oenb[0] la1_oenb[10] la1_oenb[11] la1_oenb[12] la1_oenb[13] la1_oenb[14] la1_oenb[15]
+ la1_oenb[16] la1_oenb[17] la1_oenb[18] la1_oenb[19] la1_oenb[1] la1_oenb[20] la1_oenb[21]
+ la1_oenb[22] la1_oenb[23] la1_oenb[24] la1_oenb[25] la1_oenb[26] la1_oenb[27] la1_oenb[28]
+ la1_oenb[29] la1_oenb[2] la1_oenb[30] la1_oenb[31] la1_oenb[3] la1_oenb[4] la1_oenb[5]
+ la1_oenb[6] la1_oenb[7] la1_oenb[8] la1_oenb[9] rambus_wb_ack_i rambus_wb_adr_o[0]
+ rambus_wb_adr_o[1] rambus_wb_adr_o[2] rambus_wb_adr_o[3] rambus_wb_adr_o[4] rambus_wb_adr_o[5]
+ rambus_wb_adr_o[6] rambus_wb_adr_o[7] rambus_wb_adr_o[8] rambus_wb_adr_o[9] rambus_wb_clk_o
+ rambus_wb_cyc_o rambus_wb_dat_i[0] rambus_wb_dat_i[10] rambus_wb_dat_i[11] rambus_wb_dat_i[12]
+ rambus_wb_dat_i[13] rambus_wb_dat_i[14] rambus_wb_dat_i[15] rambus_wb_dat_i[16]
+ rambus_wb_dat_i[17] rambus_wb_dat_i[18] rambus_wb_dat_i[19] rambus_wb_dat_i[1] rambus_wb_dat_i[20]
+ rambus_wb_dat_i[21] rambus_wb_dat_i[22] rambus_wb_dat_i[23] rambus_wb_dat_i[24]
+ rambus_wb_dat_i[25] rambus_wb_dat_i[26] rambus_wb_dat_i[27] rambus_wb_dat_i[28]
+ rambus_wb_dat_i[29] rambus_wb_dat_i[2] rambus_wb_dat_i[30] rambus_wb_dat_i[31] rambus_wb_dat_i[3]
+ rambus_wb_dat_i[4] rambus_wb_dat_i[5] rambus_wb_dat_i[6] rambus_wb_dat_i[7] rambus_wb_dat_i[8]
+ rambus_wb_dat_i[9] rambus_wb_dat_o[0] rambus_wb_dat_o[10] rambus_wb_dat_o[11] rambus_wb_dat_o[12]
+ rambus_wb_dat_o[13] rambus_wb_dat_o[14] rambus_wb_dat_o[15] rambus_wb_dat_o[16]
+ rambus_wb_dat_o[17] rambus_wb_dat_o[18] rambus_wb_dat_o[19] rambus_wb_dat_o[1] rambus_wb_dat_o[20]
+ rambus_wb_dat_o[21] rambus_wb_dat_o[22] rambus_wb_dat_o[23] rambus_wb_dat_o[24]
+ rambus_wb_dat_o[25] rambus_wb_dat_o[26] rambus_wb_dat_o[27] rambus_wb_dat_o[28]
+ rambus_wb_dat_o[29] rambus_wb_dat_o[2] rambus_wb_dat_o[30] rambus_wb_dat_o[31] rambus_wb_dat_o[3]
+ rambus_wb_dat_o[4] rambus_wb_dat_o[5] rambus_wb_dat_o[6] rambus_wb_dat_o[7] rambus_wb_dat_o[8]
+ rambus_wb_dat_o[9] rambus_wb_rst_o rambus_wb_sel_o[0] rambus_wb_sel_o[1] rambus_wb_sel_o[2]
+ rambus_wb_sel_o[3] rambus_wb_stb_o rambus_wb_we_o user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
.ends

* Black-box entry subcircuit for wrapped_bin_mult abstract view
.subckt wrapped_bin_mult active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
.ends

* Black-box entry subcircuit for wrapped_asic_watch abstract view
.subckt wrapped_asic_watch active io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] la1_data_in[0] la1_data_in[10] la1_data_in[11] la1_data_in[12]
+ la1_data_in[13] la1_data_in[14] la1_data_in[15] la1_data_in[16] la1_data_in[17]
+ la1_data_in[18] la1_data_in[19] la1_data_in[1] la1_data_in[20] la1_data_in[21] la1_data_in[22]
+ la1_data_in[23] la1_data_in[24] la1_data_in[25] la1_data_in[26] la1_data_in[27]
+ la1_data_in[28] la1_data_in[29] la1_data_in[2] la1_data_in[30] la1_data_in[31] la1_data_in[3]
+ la1_data_in[4] la1_data_in[5] la1_data_in[6] la1_data_in[7] la1_data_in[8] la1_data_in[9]
+ la1_data_out[0] la1_data_out[10] la1_data_out[11] la1_data_out[12] la1_data_out[13]
+ la1_data_out[14] la1_data_out[15] la1_data_out[16] la1_data_out[17] la1_data_out[18]
+ la1_data_out[19] la1_data_out[1] la1_data_out[20] la1_data_out[21] la1_data_out[22]
+ la1_data_out[23] la1_data_out[24] la1_data_out[25] la1_data_out[26] la1_data_out[27]
+ la1_data_out[28] la1_data_out[29] la1_data_out[2] la1_data_out[30] la1_data_out[31]
+ la1_data_out[3] la1_data_out[4] la1_data_out[5] la1_data_out[6] la1_data_out[7]
+ la1_data_out[8] la1_data_out[9] la1_oenb[0] la1_oenb[10] la1_oenb[11] la1_oenb[12]
+ la1_oenb[13] la1_oenb[14] la1_oenb[15] la1_oenb[16] la1_oenb[17] la1_oenb[18] la1_oenb[19]
+ la1_oenb[1] la1_oenb[20] la1_oenb[21] la1_oenb[22] la1_oenb[23] la1_oenb[24] la1_oenb[25]
+ la1_oenb[26] la1_oenb[27] la1_oenb[28] la1_oenb[29] la1_oenb[2] la1_oenb[30] la1_oenb[31]
+ la1_oenb[3] la1_oenb[4] la1_oenb[5] la1_oenb[6] la1_oenb[7] la1_oenb[8] la1_oenb[9]
+ vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
.ends

.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[2]
+ analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7] analog_io[8] analog_io[9]
+ io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14] io_in[15] io_in[16] io_in[17]
+ io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22] io_in[23] io_in[24] io_in[25]
+ io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33]
+ io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7]
+ io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14]
+ io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21]
+ io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29]
+ io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36]
+ io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9]
+ io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15] io_out[16]
+ io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22] io_out[23]
+ io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29] io_out[2] io_out[30]
+ io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36] io_out[37] io_out[3]
+ io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100]
+ la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105]
+ la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110]
+ la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115]
+ la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120]
+ la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125]
+ la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15]
+ la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20]
+ la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26]
+ la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31]
+ la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42]
+ la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48]
+ la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53]
+ la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59]
+ la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64]
+ la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6]
+ la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75]
+ la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80]
+ la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86]
+ la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91]
+ la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97]
+ la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101]
+ la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106]
+ la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110]
+ la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115]
+ la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11]
+ la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124]
+ la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13]
+ la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18]
+ la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23]
+ la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28]
+ la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33]
+ la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43]
+ la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48]
+ la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63]
+ la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68]
+ la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73]
+ la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78]
+ la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83]
+ la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88]
+ la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93]
+ la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98]
+ la_data_out[99] la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102]
+ la_oenb[103] la_oenb[104] la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109]
+ la_oenb[10] la_oenb[110] la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115]
+ la_oenb[116] la_oenb[117] la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121]
+ la_oenb[122] la_oenb[123] la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12]
+ la_oenb[13] la_oenb[14] la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19]
+ la_oenb[1] la_oenb[20] la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25]
+ la_oenb[26] la_oenb[27] la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31]
+ la_oenb[32] la_oenb[33] la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38]
+ la_oenb[39] la_oenb[3] la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44]
+ la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50]
+ la_oenb[51] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57]
+ la_oenb[58] la_oenb[59] la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63]
+ la_oenb[64] la_oenb[65] la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6]
+ la_oenb[70] la_oenb[71] la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76]
+ la_oenb[77] la_oenb[78] la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82]
+ la_oenb[83] la_oenb[84] la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89]
+ la_oenb[8] la_oenb[90] la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95]
+ la_oenb[96] la_oenb[97] la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0]
+ user_irq[1] user_irq[2] vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i
+ wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13]
+ wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19]
+ wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24]
+ wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2]
+ wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6]
+ wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11]
+ wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17]
+ wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22]
+ wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28]
+ wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4]
+ wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10]
+ wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16]
+ wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21]
+ wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27]
+ wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3]
+ wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0]
+ wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
Xwrapped_keyvalue_12 la_data_in[12] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] la_data_in[32] la_data_in[42] la_data_in[43] la_data_in[44]
+ la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[50]
+ la_data_in[51] la_data_in[33] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55]
+ la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[60] la_data_in[61]
+ la_data_in[34] la_data_in[62] la_data_in[63] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[40] la_data_in[41] la_data_out[32] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[50] la_data_out[51] la_data_out[33]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[60] la_data_out[61]
+ la_data_out[34] la_data_out[62] la_data_out[63] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[40] la_data_out[41]
+ la_oenb[32] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47]
+ la_oenb[48] la_oenb[49] la_oenb[50] la_oenb[51] la_oenb[33] la_oenb[52] la_oenb[53]
+ la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[60]
+ la_oenb[61] la_oenb[34] la_oenb[62] la_oenb[63] la_oenb[35] la_oenb[36] la_oenb[37]
+ la_oenb[38] la_oenb[39] la_oenb[40] la_oenb[41] vccd1 vssd1 wb_clk_i wb_rst_i wrapped_spell_1/wbs_ack_o
+ wrapped_spell_1/wbs_adr_i[0] wrapped_spell_1/wbs_adr_i[10] wrapped_spell_1/wbs_adr_i[11]
+ wrapped_spell_1/wbs_adr_i[12] wrapped_spell_1/wbs_adr_i[13] wrapped_spell_1/wbs_adr_i[14]
+ wrapped_spell_1/wbs_adr_i[15] wrapped_spell_1/wbs_adr_i[16] wrapped_spell_1/wbs_adr_i[17]
+ wrapped_spell_1/wbs_adr_i[18] wrapped_spell_1/wbs_adr_i[19] wrapped_spell_1/wbs_adr_i[1]
+ wrapped_spell_1/wbs_adr_i[20] wrapped_spell_1/wbs_adr_i[21] wrapped_spell_1/wbs_adr_i[22]
+ wrapped_spell_1/wbs_adr_i[23] wrapped_spell_1/wbs_adr_i[24] wrapped_spell_1/wbs_adr_i[25]
+ wrapped_spell_1/wbs_adr_i[26] wrapped_spell_1/wbs_adr_i[27] wrapped_spell_1/wbs_adr_i[28]
+ wrapped_spell_1/wbs_adr_i[29] wrapped_spell_1/wbs_adr_i[2] wrapped_spell_1/wbs_adr_i[30]
+ wrapped_spell_1/wbs_adr_i[31] wrapped_spell_1/wbs_adr_i[3] wrapped_spell_1/wbs_adr_i[4]
+ wrapped_spell_1/wbs_adr_i[5] wrapped_spell_1/wbs_adr_i[6] wrapped_spell_1/wbs_adr_i[7]
+ wrapped_spell_1/wbs_adr_i[8] wrapped_spell_1/wbs_adr_i[9] wrapped_spell_1/wbs_cyc_i
+ wrapped_spell_1/wbs_dat_i[0] wrapped_spell_1/wbs_dat_i[10] wrapped_spell_1/wbs_dat_i[11]
+ wrapped_spell_1/wbs_dat_i[12] wrapped_spell_1/wbs_dat_i[13] wrapped_spell_1/wbs_dat_i[14]
+ wrapped_spell_1/wbs_dat_i[15] wrapped_spell_1/wbs_dat_i[16] wrapped_spell_1/wbs_dat_i[17]
+ wrapped_spell_1/wbs_dat_i[18] wrapped_spell_1/wbs_dat_i[19] wrapped_spell_1/wbs_dat_i[1]
+ wrapped_spell_1/wbs_dat_i[20] wrapped_spell_1/wbs_dat_i[21] wrapped_spell_1/wbs_dat_i[22]
+ wrapped_spell_1/wbs_dat_i[23] wrapped_spell_1/wbs_dat_i[24] wrapped_spell_1/wbs_dat_i[25]
+ wrapped_spell_1/wbs_dat_i[26] wrapped_spell_1/wbs_dat_i[27] wrapped_spell_1/wbs_dat_i[28]
+ wrapped_spell_1/wbs_dat_i[29] wrapped_spell_1/wbs_dat_i[2] wrapped_spell_1/wbs_dat_i[30]
+ wrapped_spell_1/wbs_dat_i[31] wrapped_spell_1/wbs_dat_i[3] wrapped_spell_1/wbs_dat_i[4]
+ wrapped_spell_1/wbs_dat_i[5] wrapped_spell_1/wbs_dat_i[6] wrapped_spell_1/wbs_dat_i[7]
+ wrapped_spell_1/wbs_dat_i[8] wrapped_spell_1/wbs_dat_i[9] wrapped_spell_1/wbs_dat_o[0]
+ wrapped_spell_1/wbs_dat_o[10] wrapped_spell_1/wbs_dat_o[11] wrapped_spell_1/wbs_dat_o[12]
+ wrapped_spell_1/wbs_dat_o[13] wrapped_spell_1/wbs_dat_o[14] wrapped_spell_1/wbs_dat_o[15]
+ wrapped_spell_1/wbs_dat_o[16] wrapped_spell_1/wbs_dat_o[17] wrapped_spell_1/wbs_dat_o[18]
+ wrapped_spell_1/wbs_dat_o[19] wrapped_spell_1/wbs_dat_o[1] wrapped_spell_1/wbs_dat_o[20]
+ wrapped_spell_1/wbs_dat_o[21] wrapped_spell_1/wbs_dat_o[22] wrapped_spell_1/wbs_dat_o[23]
+ wrapped_spell_1/wbs_dat_o[24] wrapped_spell_1/wbs_dat_o[25] wrapped_spell_1/wbs_dat_o[26]
+ wrapped_spell_1/wbs_dat_o[27] wrapped_spell_1/wbs_dat_o[28] wrapped_spell_1/wbs_dat_o[29]
+ wrapped_spell_1/wbs_dat_o[2] wrapped_spell_1/wbs_dat_o[30] wrapped_spell_1/wbs_dat_o[31]
+ wrapped_spell_1/wbs_dat_o[3] wrapped_spell_1/wbs_dat_o[4] wrapped_spell_1/wbs_dat_o[5]
+ wrapped_spell_1/wbs_dat_o[6] wrapped_spell_1/wbs_dat_o[7] wrapped_spell_1/wbs_dat_o[8]
+ wrapped_spell_1/wbs_dat_o[9] wrapped_spell_1/wbs_sel_i[0] wrapped_spell_1/wbs_sel_i[1]
+ wrapped_spell_1/wbs_sel_i[2] wrapped_spell_1/wbs_sel_i[3] wrapped_spell_1/wbs_stb_i
+ wrapped_spell_1/wbs_we_i wrapped_keyvalue
Xwrapped_ppm_coder_2 la_data_in[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] vccd1 vssd1 wb_clk_i wrapped_ppm_coder
Xwrapped_silife_4 la_data_in[4] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[32] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46]
+ la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[50] la_data_in[51] la_data_in[33]
+ la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57]
+ la_data_in[58] la_data_in[59] la_data_in[60] la_data_in[61] la_data_in[34] la_data_in[62]
+ la_data_in[63] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39]
+ la_data_in[40] la_data_in[41] la_data_out[32] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[50] la_data_out[51] la_data_out[33] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[60] la_data_out[61] la_data_out[34] la_data_out[62]
+ la_data_out[63] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[40] la_data_out[41] la_oenb[32] la_oenb[42] la_oenb[43]
+ la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[50]
+ la_oenb[51] la_oenb[33] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56]
+ la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[60] la_oenb[61] la_oenb[34] la_oenb[62]
+ la_oenb[63] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[40]
+ la_oenb[41] vccd1 vssd1 wb_clk_i wb_rst_i wrapped_spell_1/wbs_ack_o wrapped_spell_1/wbs_adr_i[0]
+ wrapped_spell_1/wbs_adr_i[10] wrapped_spell_1/wbs_adr_i[11] wrapped_spell_1/wbs_adr_i[12]
+ wrapped_spell_1/wbs_adr_i[13] wrapped_spell_1/wbs_adr_i[14] wrapped_spell_1/wbs_adr_i[15]
+ wrapped_spell_1/wbs_adr_i[16] wrapped_spell_1/wbs_adr_i[17] wrapped_spell_1/wbs_adr_i[18]
+ wrapped_spell_1/wbs_adr_i[19] wrapped_spell_1/wbs_adr_i[1] wrapped_spell_1/wbs_adr_i[20]
+ wrapped_spell_1/wbs_adr_i[21] wrapped_spell_1/wbs_adr_i[22] wrapped_spell_1/wbs_adr_i[23]
+ wrapped_spell_1/wbs_adr_i[24] wrapped_spell_1/wbs_adr_i[25] wrapped_spell_1/wbs_adr_i[26]
+ wrapped_spell_1/wbs_adr_i[27] wrapped_spell_1/wbs_adr_i[28] wrapped_spell_1/wbs_adr_i[29]
+ wrapped_spell_1/wbs_adr_i[2] wrapped_spell_1/wbs_adr_i[30] wrapped_spell_1/wbs_adr_i[31]
+ wrapped_spell_1/wbs_adr_i[3] wrapped_spell_1/wbs_adr_i[4] wrapped_spell_1/wbs_adr_i[5]
+ wrapped_spell_1/wbs_adr_i[6] wrapped_spell_1/wbs_adr_i[7] wrapped_spell_1/wbs_adr_i[8]
+ wrapped_spell_1/wbs_adr_i[9] wrapped_spell_1/wbs_cyc_i wrapped_spell_1/wbs_dat_i[0]
+ wrapped_spell_1/wbs_dat_i[10] wrapped_spell_1/wbs_dat_i[11] wrapped_spell_1/wbs_dat_i[12]
+ wrapped_spell_1/wbs_dat_i[13] wrapped_spell_1/wbs_dat_i[14] wrapped_spell_1/wbs_dat_i[15]
+ wrapped_spell_1/wbs_dat_i[16] wrapped_spell_1/wbs_dat_i[17] wrapped_spell_1/wbs_dat_i[18]
+ wrapped_spell_1/wbs_dat_i[19] wrapped_spell_1/wbs_dat_i[1] wrapped_spell_1/wbs_dat_i[20]
+ wrapped_spell_1/wbs_dat_i[21] wrapped_spell_1/wbs_dat_i[22] wrapped_spell_1/wbs_dat_i[23]
+ wrapped_spell_1/wbs_dat_i[24] wrapped_spell_1/wbs_dat_i[25] wrapped_spell_1/wbs_dat_i[26]
+ wrapped_spell_1/wbs_dat_i[27] wrapped_spell_1/wbs_dat_i[28] wrapped_spell_1/wbs_dat_i[29]
+ wrapped_spell_1/wbs_dat_i[2] wrapped_spell_1/wbs_dat_i[30] wrapped_spell_1/wbs_dat_i[31]
+ wrapped_spell_1/wbs_dat_i[3] wrapped_spell_1/wbs_dat_i[4] wrapped_spell_1/wbs_dat_i[5]
+ wrapped_spell_1/wbs_dat_i[6] wrapped_spell_1/wbs_dat_i[7] wrapped_spell_1/wbs_dat_i[8]
+ wrapped_spell_1/wbs_dat_i[9] wrapped_spell_1/wbs_dat_o[0] wrapped_spell_1/wbs_dat_o[10]
+ wrapped_spell_1/wbs_dat_o[11] wrapped_spell_1/wbs_dat_o[12] wrapped_spell_1/wbs_dat_o[13]
+ wrapped_spell_1/wbs_dat_o[14] wrapped_spell_1/wbs_dat_o[15] wrapped_spell_1/wbs_dat_o[16]
+ wrapped_spell_1/wbs_dat_o[17] wrapped_spell_1/wbs_dat_o[18] wrapped_spell_1/wbs_dat_o[19]
+ wrapped_spell_1/wbs_dat_o[1] wrapped_spell_1/wbs_dat_o[20] wrapped_spell_1/wbs_dat_o[21]
+ wrapped_spell_1/wbs_dat_o[22] wrapped_spell_1/wbs_dat_o[23] wrapped_spell_1/wbs_dat_o[24]
+ wrapped_spell_1/wbs_dat_o[25] wrapped_spell_1/wbs_dat_o[26] wrapped_spell_1/wbs_dat_o[27]
+ wrapped_spell_1/wbs_dat_o[28] wrapped_spell_1/wbs_dat_o[29] wrapped_spell_1/wbs_dat_o[2]
+ wrapped_spell_1/wbs_dat_o[30] wrapped_spell_1/wbs_dat_o[31] wrapped_spell_1/wbs_dat_o[3]
+ wrapped_spell_1/wbs_dat_o[4] wrapped_spell_1/wbs_dat_o[5] wrapped_spell_1/wbs_dat_o[6]
+ wrapped_spell_1/wbs_dat_o[7] wrapped_spell_1/wbs_dat_o[8] wrapped_spell_1/wbs_dat_o[9]
+ wrapped_spell_1/wbs_sel_i[0] wrapped_spell_1/wbs_sel_i[1] wrapped_spell_1/wbs_sel_i[2]
+ wrapped_spell_1/wbs_sel_i[3] wrapped_spell_1/wbs_stb_i wrapped_spell_1/wbs_we_i
+ wrapped_silife
Xwrapped_spraid_6 la_data_in[6] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ vccd1 vssd1 wb_clk_i wb_rst_i wrapped_spell_1/wbs_ack_o wrapped_spell_1/wbs_adr_i[0]
+ wrapped_spell_1/wbs_adr_i[10] wrapped_spell_1/wbs_adr_i[11] wrapped_spell_1/wbs_adr_i[12]
+ wrapped_spell_1/wbs_adr_i[13] wrapped_spell_1/wbs_adr_i[14] wrapped_spell_1/wbs_adr_i[15]
+ wrapped_spell_1/wbs_adr_i[16] wrapped_spell_1/wbs_adr_i[17] wrapped_spell_1/wbs_adr_i[18]
+ wrapped_spell_1/wbs_adr_i[19] wrapped_spell_1/wbs_adr_i[1] wrapped_spell_1/wbs_adr_i[20]
+ wrapped_spell_1/wbs_adr_i[21] wrapped_spell_1/wbs_adr_i[22] wrapped_spell_1/wbs_adr_i[23]
+ wrapped_spell_1/wbs_adr_i[24] wrapped_spell_1/wbs_adr_i[25] wrapped_spell_1/wbs_adr_i[26]
+ wrapped_spell_1/wbs_adr_i[27] wrapped_spell_1/wbs_adr_i[28] wrapped_spell_1/wbs_adr_i[29]
+ wrapped_spell_1/wbs_adr_i[2] wrapped_spell_1/wbs_adr_i[30] wrapped_spell_1/wbs_adr_i[31]
+ wrapped_spell_1/wbs_adr_i[3] wrapped_spell_1/wbs_adr_i[4] wrapped_spell_1/wbs_adr_i[5]
+ wrapped_spell_1/wbs_adr_i[6] wrapped_spell_1/wbs_adr_i[7] wrapped_spell_1/wbs_adr_i[8]
+ wrapped_spell_1/wbs_adr_i[9] wrapped_spell_1/wbs_cyc_i wrapped_spell_1/wbs_dat_i[0]
+ wrapped_spell_1/wbs_dat_i[10] wrapped_spell_1/wbs_dat_i[11] wrapped_spell_1/wbs_dat_i[12]
+ wrapped_spell_1/wbs_dat_i[13] wrapped_spell_1/wbs_dat_i[14] wrapped_spell_1/wbs_dat_i[15]
+ wrapped_spell_1/wbs_dat_i[16] wrapped_spell_1/wbs_dat_i[17] wrapped_spell_1/wbs_dat_i[18]
+ wrapped_spell_1/wbs_dat_i[19] wrapped_spell_1/wbs_dat_i[1] wrapped_spell_1/wbs_dat_i[20]
+ wrapped_spell_1/wbs_dat_i[21] wrapped_spell_1/wbs_dat_i[22] wrapped_spell_1/wbs_dat_i[23]
+ wrapped_spell_1/wbs_dat_i[24] wrapped_spell_1/wbs_dat_i[25] wrapped_spell_1/wbs_dat_i[26]
+ wrapped_spell_1/wbs_dat_i[27] wrapped_spell_1/wbs_dat_i[28] wrapped_spell_1/wbs_dat_i[29]
+ wrapped_spell_1/wbs_dat_i[2] wrapped_spell_1/wbs_dat_i[30] wrapped_spell_1/wbs_dat_i[31]
+ wrapped_spell_1/wbs_dat_i[3] wrapped_spell_1/wbs_dat_i[4] wrapped_spell_1/wbs_dat_i[5]
+ wrapped_spell_1/wbs_dat_i[6] wrapped_spell_1/wbs_dat_i[7] wrapped_spell_1/wbs_dat_i[8]
+ wrapped_spell_1/wbs_dat_i[9] wrapped_spell_1/wbs_dat_o[0] wrapped_spell_1/wbs_dat_o[10]
+ wrapped_spell_1/wbs_dat_o[11] wrapped_spell_1/wbs_dat_o[12] wrapped_spell_1/wbs_dat_o[13]
+ wrapped_spell_1/wbs_dat_o[14] wrapped_spell_1/wbs_dat_o[15] wrapped_spell_1/wbs_dat_o[16]
+ wrapped_spell_1/wbs_dat_o[17] wrapped_spell_1/wbs_dat_o[18] wrapped_spell_1/wbs_dat_o[19]
+ wrapped_spell_1/wbs_dat_o[1] wrapped_spell_1/wbs_dat_o[20] wrapped_spell_1/wbs_dat_o[21]
+ wrapped_spell_1/wbs_dat_o[22] wrapped_spell_1/wbs_dat_o[23] wrapped_spell_1/wbs_dat_o[24]
+ wrapped_spell_1/wbs_dat_o[25] wrapped_spell_1/wbs_dat_o[26] wrapped_spell_1/wbs_dat_o[27]
+ wrapped_spell_1/wbs_dat_o[28] wrapped_spell_1/wbs_dat_o[29] wrapped_spell_1/wbs_dat_o[2]
+ wrapped_spell_1/wbs_dat_o[30] wrapped_spell_1/wbs_dat_o[31] wrapped_spell_1/wbs_dat_o[3]
+ wrapped_spell_1/wbs_dat_o[4] wrapped_spell_1/wbs_dat_o[5] wrapped_spell_1/wbs_dat_o[6]
+ wrapped_spell_1/wbs_dat_o[7] wrapped_spell_1/wbs_dat_o[8] wrapped_spell_1/wbs_dat_o[9]
+ wrapped_spell_1/wbs_sel_i[0] wrapped_spell_1/wbs_sel_i[1] wrapped_spell_1/wbs_sel_i[2]
+ wrapped_spell_1/wbs_sel_i[3] wrapped_spell_1/wbs_stb_i wrapped_spell_1/wbs_we_i
+ wrapped_spraid
Xwb_bridge_2way vccd1 vssd1 wb_clk_i wb_rst_i wrapped_spell_1/wbs_ack_o wrapped_spell_1/wbs_adr_i[0]
+ wrapped_spell_1/wbs_adr_i[10] wrapped_spell_1/wbs_adr_i[11] wrapped_spell_1/wbs_adr_i[12]
+ wrapped_spell_1/wbs_adr_i[13] wrapped_spell_1/wbs_adr_i[14] wrapped_spell_1/wbs_adr_i[15]
+ wrapped_spell_1/wbs_adr_i[16] wrapped_spell_1/wbs_adr_i[17] wrapped_spell_1/wbs_adr_i[18]
+ wrapped_spell_1/wbs_adr_i[19] wrapped_spell_1/wbs_adr_i[1] wrapped_spell_1/wbs_adr_i[20]
+ wrapped_spell_1/wbs_adr_i[21] wrapped_spell_1/wbs_adr_i[22] wrapped_spell_1/wbs_adr_i[23]
+ wrapped_spell_1/wbs_adr_i[24] wrapped_spell_1/wbs_adr_i[25] wrapped_spell_1/wbs_adr_i[26]
+ wrapped_spell_1/wbs_adr_i[27] wrapped_spell_1/wbs_adr_i[28] wrapped_spell_1/wbs_adr_i[29]
+ wrapped_spell_1/wbs_adr_i[2] wrapped_spell_1/wbs_adr_i[30] wrapped_spell_1/wbs_adr_i[31]
+ wrapped_spell_1/wbs_adr_i[3] wrapped_spell_1/wbs_adr_i[4] wrapped_spell_1/wbs_adr_i[5]
+ wrapped_spell_1/wbs_adr_i[6] wrapped_spell_1/wbs_adr_i[7] wrapped_spell_1/wbs_adr_i[8]
+ wrapped_spell_1/wbs_adr_i[9] wrapped_spell_1/wbs_cyc_i wrapped_spell_1/wbs_dat_o[0]
+ wrapped_spell_1/wbs_dat_o[10] wrapped_spell_1/wbs_dat_o[11] wrapped_spell_1/wbs_dat_o[12]
+ wrapped_spell_1/wbs_dat_o[13] wrapped_spell_1/wbs_dat_o[14] wrapped_spell_1/wbs_dat_o[15]
+ wrapped_spell_1/wbs_dat_o[16] wrapped_spell_1/wbs_dat_o[17] wrapped_spell_1/wbs_dat_o[18]
+ wrapped_spell_1/wbs_dat_o[19] wrapped_spell_1/wbs_dat_o[1] wrapped_spell_1/wbs_dat_o[20]
+ wrapped_spell_1/wbs_dat_o[21] wrapped_spell_1/wbs_dat_o[22] wrapped_spell_1/wbs_dat_o[23]
+ wrapped_spell_1/wbs_dat_o[24] wrapped_spell_1/wbs_dat_o[25] wrapped_spell_1/wbs_dat_o[26]
+ wrapped_spell_1/wbs_dat_o[27] wrapped_spell_1/wbs_dat_o[28] wrapped_spell_1/wbs_dat_o[29]
+ wrapped_spell_1/wbs_dat_o[2] wrapped_spell_1/wbs_dat_o[30] wrapped_spell_1/wbs_dat_o[31]
+ wrapped_spell_1/wbs_dat_o[3] wrapped_spell_1/wbs_dat_o[4] wrapped_spell_1/wbs_dat_o[5]
+ wrapped_spell_1/wbs_dat_o[6] wrapped_spell_1/wbs_dat_o[7] wrapped_spell_1/wbs_dat_o[8]
+ wrapped_spell_1/wbs_dat_o[9] wrapped_spell_1/wbs_dat_i[0] wrapped_spell_1/wbs_dat_i[10]
+ wrapped_spell_1/wbs_dat_i[11] wrapped_spell_1/wbs_dat_i[12] wrapped_spell_1/wbs_dat_i[13]
+ wrapped_spell_1/wbs_dat_i[14] wrapped_spell_1/wbs_dat_i[15] wrapped_spell_1/wbs_dat_i[16]
+ wrapped_spell_1/wbs_dat_i[17] wrapped_spell_1/wbs_dat_i[18] wrapped_spell_1/wbs_dat_i[19]
+ wrapped_spell_1/wbs_dat_i[1] wrapped_spell_1/wbs_dat_i[20] wrapped_spell_1/wbs_dat_i[21]
+ wrapped_spell_1/wbs_dat_i[22] wrapped_spell_1/wbs_dat_i[23] wrapped_spell_1/wbs_dat_i[24]
+ wrapped_spell_1/wbs_dat_i[25] wrapped_spell_1/wbs_dat_i[26] wrapped_spell_1/wbs_dat_i[27]
+ wrapped_spell_1/wbs_dat_i[28] wrapped_spell_1/wbs_dat_i[29] wrapped_spell_1/wbs_dat_i[2]
+ wrapped_spell_1/wbs_dat_i[30] wrapped_spell_1/wbs_dat_i[31] wrapped_spell_1/wbs_dat_i[3]
+ wrapped_spell_1/wbs_dat_i[4] wrapped_spell_1/wbs_dat_i[5] wrapped_spell_1/wbs_dat_i[6]
+ wrapped_spell_1/wbs_dat_i[7] wrapped_spell_1/wbs_dat_i[8] wrapped_spell_1/wbs_dat_i[9]
+ wrapped_spell_1/wbs_sel_i[0] wrapped_spell_1/wbs_sel_i[1] wrapped_spell_1/wbs_sel_i[2]
+ wrapped_spell_1/wbs_sel_i[3] wrapped_spell_1/wbs_stb_i wrapped_spell_1/wbs_we_i
+ wb_bridge_2way/wbm_b_ack_i wb_bridge_2way/wbm_b_adr_o[0] wb_bridge_2way/wbm_b_adr_o[1]
+ wb_bridge_2way/wbm_b_adr_o[2] wb_bridge_2way/wbm_b_adr_o[3] wb_bridge_2way/wbm_b_adr_o[4]
+ wb_bridge_2way/wbm_b_adr_o[5] wb_bridge_2way/wbm_b_adr_o[6] wb_bridge_2way/wbm_b_adr_o[7]
+ wb_bridge_2way/wbm_b_adr_o[8] wb_bridge_2way/wbm_b_adr_o[9] wb_bridge_2way/wbm_b_cyc_o
+ wb_bridge_2way/wbm_b_dat_i[0] wb_bridge_2way/wbm_b_dat_i[10] wb_bridge_2way/wbm_b_dat_i[11]
+ wb_bridge_2way/wbm_b_dat_i[12] wb_bridge_2way/wbm_b_dat_i[13] wb_bridge_2way/wbm_b_dat_i[14]
+ wb_bridge_2way/wbm_b_dat_i[15] wb_bridge_2way/wbm_b_dat_i[16] wb_bridge_2way/wbm_b_dat_i[17]
+ wb_bridge_2way/wbm_b_dat_i[18] wb_bridge_2way/wbm_b_dat_i[19] wb_bridge_2way/wbm_b_dat_i[1]
+ wb_bridge_2way/wbm_b_dat_i[20] wb_bridge_2way/wbm_b_dat_i[21] wb_bridge_2way/wbm_b_dat_i[22]
+ wb_bridge_2way/wbm_b_dat_i[23] wb_bridge_2way/wbm_b_dat_i[24] wb_bridge_2way/wbm_b_dat_i[25]
+ wb_bridge_2way/wbm_b_dat_i[26] wb_bridge_2way/wbm_b_dat_i[27] wb_bridge_2way/wbm_b_dat_i[28]
+ wb_bridge_2way/wbm_b_dat_i[29] wb_bridge_2way/wbm_b_dat_i[2] wb_bridge_2way/wbm_b_dat_i[30]
+ wb_bridge_2way/wbm_b_dat_i[31] wb_bridge_2way/wbm_b_dat_i[3] wb_bridge_2way/wbm_b_dat_i[4]
+ wb_bridge_2way/wbm_b_dat_i[5] wb_bridge_2way/wbm_b_dat_i[6] wb_bridge_2way/wbm_b_dat_i[7]
+ wb_bridge_2way/wbm_b_dat_i[8] wb_bridge_2way/wbm_b_dat_i[9] wb_bridge_2way/wbm_b_dat_o[0]
+ wb_bridge_2way/wbm_b_dat_o[10] wb_bridge_2way/wbm_b_dat_o[11] wb_bridge_2way/wbm_b_dat_o[12]
+ wb_bridge_2way/wbm_b_dat_o[13] wb_bridge_2way/wbm_b_dat_o[14] wb_bridge_2way/wbm_b_dat_o[15]
+ wb_bridge_2way/wbm_b_dat_o[16] wb_bridge_2way/wbm_b_dat_o[17] wb_bridge_2way/wbm_b_dat_o[18]
+ wb_bridge_2way/wbm_b_dat_o[19] wb_bridge_2way/wbm_b_dat_o[1] wb_bridge_2way/wbm_b_dat_o[20]
+ wb_bridge_2way/wbm_b_dat_o[21] wb_bridge_2way/wbm_b_dat_o[22] wb_bridge_2way/wbm_b_dat_o[23]
+ wb_bridge_2way/wbm_b_dat_o[24] wb_bridge_2way/wbm_b_dat_o[25] wb_bridge_2way/wbm_b_dat_o[26]
+ wb_bridge_2way/wbm_b_dat_o[27] wb_bridge_2way/wbm_b_dat_o[28] wb_bridge_2way/wbm_b_dat_o[29]
+ wb_bridge_2way/wbm_b_dat_o[2] wb_bridge_2way/wbm_b_dat_o[30] wb_bridge_2way/wbm_b_dat_o[31]
+ wb_bridge_2way/wbm_b_dat_o[3] wb_bridge_2way/wbm_b_dat_o[4] wb_bridge_2way/wbm_b_dat_o[5]
+ wb_bridge_2way/wbm_b_dat_o[6] wb_bridge_2way/wbm_b_dat_o[7] wb_bridge_2way/wbm_b_dat_o[8]
+ wb_bridge_2way/wbm_b_dat_o[9] wb_bridge_2way/wbm_b_sel_o[0] wb_bridge_2way/wbm_b_sel_o[1]
+ wb_bridge_2way/wbm_b_sel_o[2] wb_bridge_2way/wbm_b_sel_o[3] wb_bridge_2way/wbm_b_stb_o
+ wb_bridge_2way/wbm_b_we_o wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i wb_bridge_2way
Xopenram_1kB openram_1kB/din0[0] openram_1kB/din0[1] openram_1kB/din0[2] openram_1kB/din0[3]
+ openram_1kB/din0[4] openram_1kB/din0[5] openram_1kB/din0[6] openram_1kB/din0[7]
+ openram_1kB/din0[8] openram_1kB/din0[9] openram_1kB/din0[10] openram_1kB/din0[11]
+ openram_1kB/din0[12] openram_1kB/din0[13] openram_1kB/din0[14] openram_1kB/din0[15]
+ openram_1kB/din0[16] openram_1kB/din0[17] openram_1kB/din0[18] openram_1kB/din0[19]
+ openram_1kB/din0[20] openram_1kB/din0[21] openram_1kB/din0[22] openram_1kB/din0[23]
+ openram_1kB/din0[24] openram_1kB/din0[25] openram_1kB/din0[26] openram_1kB/din0[27]
+ openram_1kB/din0[28] openram_1kB/din0[29] openram_1kB/din0[30] openram_1kB/din0[31]
+ openram_1kB/addr0[0] openram_1kB/addr0[1] openram_1kB/addr0[2] openram_1kB/addr0[3]
+ openram_1kB/addr0[4] openram_1kB/addr0[5] openram_1kB/addr0[6] openram_1kB/addr0[7]
+ openram_1kB/addr1[0] openram_1kB/addr1[1] openram_1kB/addr1[2] openram_1kB/addr1[3]
+ openram_1kB/addr1[4] openram_1kB/addr1[5] openram_1kB/addr1[6] openram_1kB/addr1[7]
+ openram_1kB/csb0 openram_1kB/csb1 openram_1kB/web0 openram_1kB/clk0 openram_1kB/clk1
+ openram_1kB/wmask0[0] openram_1kB/wmask0[1] openram_1kB/wmask0[2] openram_1kB/wmask0[3]
+ openram_1kB/dout0[0] openram_1kB/dout0[1] openram_1kB/dout0[2] openram_1kB/dout0[3]
+ openram_1kB/dout0[4] openram_1kB/dout0[5] openram_1kB/dout0[6] openram_1kB/dout0[7]
+ openram_1kB/dout0[8] openram_1kB/dout0[9] openram_1kB/dout0[10] openram_1kB/dout0[11]
+ openram_1kB/dout0[12] openram_1kB/dout0[13] openram_1kB/dout0[14] openram_1kB/dout0[15]
+ openram_1kB/dout0[16] openram_1kB/dout0[17] openram_1kB/dout0[18] openram_1kB/dout0[19]
+ openram_1kB/dout0[20] openram_1kB/dout0[21] openram_1kB/dout0[22] openram_1kB/dout0[23]
+ openram_1kB/dout0[24] openram_1kB/dout0[25] openram_1kB/dout0[26] openram_1kB/dout0[27]
+ openram_1kB/dout0[28] openram_1kB/dout0[29] openram_1kB/dout0[30] openram_1kB/dout0[31]
+ openram_1kB/dout1[0] openram_1kB/dout1[1] openram_1kB/dout1[2] openram_1kB/dout1[3]
+ openram_1kB/dout1[4] openram_1kB/dout1[5] openram_1kB/dout1[6] openram_1kB/dout1[7]
+ openram_1kB/dout1[8] openram_1kB/dout1[9] openram_1kB/dout1[10] openram_1kB/dout1[11]
+ openram_1kB/dout1[12] openram_1kB/dout1[13] openram_1kB/dout1[14] openram_1kB/dout1[15]
+ openram_1kB/dout1[16] openram_1kB/dout1[17] openram_1kB/dout1[18] openram_1kB/dout1[19]
+ openram_1kB/dout1[20] openram_1kB/dout1[21] openram_1kB/dout1[22] openram_1kB/dout1[23]
+ openram_1kB/dout1[24] openram_1kB/dout1[25] openram_1kB/dout1[26] openram_1kB/dout1[27]
+ openram_1kB/dout1[28] openram_1kB/dout1[29] openram_1kB/dout1[30] openram_1kB/dout1[31]
+ vccd1 vssd1 sky130_sram_1kbyte_1rw1r_32x256_8
Xwrapped_skullfet_5 la_data_in[5] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] la_data_in[32] la_data_in[42] la_data_in[43] la_data_in[44]
+ la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[50]
+ la_data_in[51] la_data_in[33] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55]
+ la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[60] la_data_in[61]
+ la_data_in[34] la_data_in[62] la_data_in[63] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[40] la_data_in[41] la_data_out[32] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[50] la_data_out[51] la_data_out[33]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[60] la_data_out[61]
+ la_data_out[34] la_data_out[62] la_data_out[63] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[40] la_data_out[41]
+ la_oenb[32] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47]
+ la_oenb[48] la_oenb[49] la_oenb[50] la_oenb[51] la_oenb[33] la_oenb[52] la_oenb[53]
+ la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[60]
+ la_oenb[61] la_oenb[34] la_oenb[62] la_oenb[63] la_oenb[35] la_oenb[36] la_oenb[37]
+ la_oenb[38] la_oenb[39] la_oenb[40] la_oenb[41] vccd1 vssd1 wb_clk_i wrapped_skullfet
Xwb_openram_wrapper openram_1kB/addr0[0] openram_1kB/addr0[1] openram_1kB/addr0[2]
+ openram_1kB/addr0[3] openram_1kB/addr0[4] openram_1kB/addr0[5] openram_1kB/addr0[6]
+ openram_1kB/addr0[7] openram_1kB/addr1[0] openram_1kB/addr1[1] openram_1kB/addr1[2]
+ openram_1kB/addr1[3] openram_1kB/addr1[4] openram_1kB/addr1[5] openram_1kB/addr1[6]
+ openram_1kB/addr1[7] openram_1kB/clk0 openram_1kB/clk1 openram_1kB/csb0 openram_1kB/csb1
+ openram_1kB/din0[0] openram_1kB/din0[10] openram_1kB/din0[11] openram_1kB/din0[12]
+ openram_1kB/din0[13] openram_1kB/din0[14] openram_1kB/din0[15] openram_1kB/din0[16]
+ openram_1kB/din0[17] openram_1kB/din0[18] openram_1kB/din0[19] openram_1kB/din0[1]
+ openram_1kB/din0[20] openram_1kB/din0[21] openram_1kB/din0[22] openram_1kB/din0[23]
+ openram_1kB/din0[24] openram_1kB/din0[25] openram_1kB/din0[26] openram_1kB/din0[27]
+ openram_1kB/din0[28] openram_1kB/din0[29] openram_1kB/din0[2] openram_1kB/din0[30]
+ openram_1kB/din0[31] openram_1kB/din0[3] openram_1kB/din0[4] openram_1kB/din0[5]
+ openram_1kB/din0[6] openram_1kB/din0[7] openram_1kB/din0[8] openram_1kB/din0[9]
+ openram_1kB/dout0[0] openram_1kB/dout0[10] openram_1kB/dout0[11] openram_1kB/dout0[12]
+ openram_1kB/dout0[13] openram_1kB/dout0[14] openram_1kB/dout0[15] openram_1kB/dout0[16]
+ openram_1kB/dout0[17] openram_1kB/dout0[18] openram_1kB/dout0[19] openram_1kB/dout0[1]
+ openram_1kB/dout0[20] openram_1kB/dout0[21] openram_1kB/dout0[22] openram_1kB/dout0[23]
+ openram_1kB/dout0[24] openram_1kB/dout0[25] openram_1kB/dout0[26] openram_1kB/dout0[27]
+ openram_1kB/dout0[28] openram_1kB/dout0[29] openram_1kB/dout0[2] openram_1kB/dout0[30]
+ openram_1kB/dout0[31] openram_1kB/dout0[3] openram_1kB/dout0[4] openram_1kB/dout0[5]
+ openram_1kB/dout0[6] openram_1kB/dout0[7] openram_1kB/dout0[8] openram_1kB/dout0[9]
+ openram_1kB/dout1[0] openram_1kB/dout1[10] openram_1kB/dout1[11] openram_1kB/dout1[12]
+ openram_1kB/dout1[13] openram_1kB/dout1[14] openram_1kB/dout1[15] openram_1kB/dout1[16]
+ openram_1kB/dout1[17] openram_1kB/dout1[18] openram_1kB/dout1[19] openram_1kB/dout1[1]
+ openram_1kB/dout1[20] openram_1kB/dout1[21] openram_1kB/dout1[22] openram_1kB/dout1[23]
+ openram_1kB/dout1[24] openram_1kB/dout1[25] openram_1kB/dout1[26] openram_1kB/dout1[27]
+ openram_1kB/dout1[28] openram_1kB/dout1[29] openram_1kB/dout1[2] openram_1kB/dout1[30]
+ openram_1kB/dout1[31] openram_1kB/dout1[3] openram_1kB/dout1[4] openram_1kB/dout1[5]
+ openram_1kB/dout1[6] openram_1kB/dout1[7] openram_1kB/dout1[8] openram_1kB/dout1[9]
+ openram_1kB/web0 openram_1kB/wmask0[0] openram_1kB/wmask0[1] openram_1kB/wmask0[2]
+ openram_1kB/wmask0[3] vccd1 vssd1 wb_clk_i wb_rst_i wb_openram_wrapper/wb_b_clk_i
+ wb_openram_wrapper/wb_b_rst_i wb_bridge_2way/wbm_b_ack_i wb_bridge_2way/wbm_b_adr_o[0]
+ wb_bridge_2way/wbm_b_adr_o[1] wb_bridge_2way/wbm_b_adr_o[2] wb_bridge_2way/wbm_b_adr_o[3]
+ wb_bridge_2way/wbm_b_adr_o[4] wb_bridge_2way/wbm_b_adr_o[5] wb_bridge_2way/wbm_b_adr_o[6]
+ wb_bridge_2way/wbm_b_adr_o[7] wb_bridge_2way/wbm_b_adr_o[8] wb_bridge_2way/wbm_b_adr_o[9]
+ wb_bridge_2way/wbm_b_cyc_o wb_bridge_2way/wbm_b_dat_o[0] wb_bridge_2way/wbm_b_dat_o[10]
+ wb_bridge_2way/wbm_b_dat_o[11] wb_bridge_2way/wbm_b_dat_o[12] wb_bridge_2way/wbm_b_dat_o[13]
+ wb_bridge_2way/wbm_b_dat_o[14] wb_bridge_2way/wbm_b_dat_o[15] wb_bridge_2way/wbm_b_dat_o[16]
+ wb_bridge_2way/wbm_b_dat_o[17] wb_bridge_2way/wbm_b_dat_o[18] wb_bridge_2way/wbm_b_dat_o[19]
+ wb_bridge_2way/wbm_b_dat_o[1] wb_bridge_2way/wbm_b_dat_o[20] wb_bridge_2way/wbm_b_dat_o[21]
+ wb_bridge_2way/wbm_b_dat_o[22] wb_bridge_2way/wbm_b_dat_o[23] wb_bridge_2way/wbm_b_dat_o[24]
+ wb_bridge_2way/wbm_b_dat_o[25] wb_bridge_2way/wbm_b_dat_o[26] wb_bridge_2way/wbm_b_dat_o[27]
+ wb_bridge_2way/wbm_b_dat_o[28] wb_bridge_2way/wbm_b_dat_o[29] wb_bridge_2way/wbm_b_dat_o[2]
+ wb_bridge_2way/wbm_b_dat_o[30] wb_bridge_2way/wbm_b_dat_o[31] wb_bridge_2way/wbm_b_dat_o[3]
+ wb_bridge_2way/wbm_b_dat_o[4] wb_bridge_2way/wbm_b_dat_o[5] wb_bridge_2way/wbm_b_dat_o[6]
+ wb_bridge_2way/wbm_b_dat_o[7] wb_bridge_2way/wbm_b_dat_o[8] wb_bridge_2way/wbm_b_dat_o[9]
+ wb_bridge_2way/wbm_b_dat_i[0] wb_bridge_2way/wbm_b_dat_i[10] wb_bridge_2way/wbm_b_dat_i[11]
+ wb_bridge_2way/wbm_b_dat_i[12] wb_bridge_2way/wbm_b_dat_i[13] wb_bridge_2way/wbm_b_dat_i[14]
+ wb_bridge_2way/wbm_b_dat_i[15] wb_bridge_2way/wbm_b_dat_i[16] wb_bridge_2way/wbm_b_dat_i[17]
+ wb_bridge_2way/wbm_b_dat_i[18] wb_bridge_2way/wbm_b_dat_i[19] wb_bridge_2way/wbm_b_dat_i[1]
+ wb_bridge_2way/wbm_b_dat_i[20] wb_bridge_2way/wbm_b_dat_i[21] wb_bridge_2way/wbm_b_dat_i[22]
+ wb_bridge_2way/wbm_b_dat_i[23] wb_bridge_2way/wbm_b_dat_i[24] wb_bridge_2way/wbm_b_dat_i[25]
+ wb_bridge_2way/wbm_b_dat_i[26] wb_bridge_2way/wbm_b_dat_i[27] wb_bridge_2way/wbm_b_dat_i[28]
+ wb_bridge_2way/wbm_b_dat_i[29] wb_bridge_2way/wbm_b_dat_i[2] wb_bridge_2way/wbm_b_dat_i[30]
+ wb_bridge_2way/wbm_b_dat_i[31] wb_bridge_2way/wbm_b_dat_i[3] wb_bridge_2way/wbm_b_dat_i[4]
+ wb_bridge_2way/wbm_b_dat_i[5] wb_bridge_2way/wbm_b_dat_i[6] wb_bridge_2way/wbm_b_dat_i[7]
+ wb_bridge_2way/wbm_b_dat_i[8] wb_bridge_2way/wbm_b_dat_i[9] wb_bridge_2way/wbm_b_sel_o[0]
+ wb_bridge_2way/wbm_b_sel_o[1] wb_bridge_2way/wbm_b_sel_o[2] wb_bridge_2way/wbm_b_sel_o[3]
+ wb_bridge_2way/wbm_b_stb_o wb_bridge_2way/wbm_b_we_o wb_openram_wrapper/wbs_b_ack_o
+ wb_openram_wrapper/wbs_b_adr_i[0] wb_openram_wrapper/wbs_b_adr_i[1] wb_openram_wrapper/wbs_b_adr_i[2]
+ wb_openram_wrapper/wbs_b_adr_i[3] wb_openram_wrapper/wbs_b_adr_i[4] wb_openram_wrapper/wbs_b_adr_i[5]
+ wb_openram_wrapper/wbs_b_adr_i[6] wb_openram_wrapper/wbs_b_adr_i[7] wb_openram_wrapper/wbs_b_adr_i[8]
+ wb_openram_wrapper/wbs_b_adr_i[9] wb_openram_wrapper/wbs_b_cyc_i wb_openram_wrapper/wbs_b_dat_i[0]
+ wb_openram_wrapper/wbs_b_dat_i[10] wb_openram_wrapper/wbs_b_dat_i[11] wb_openram_wrapper/wbs_b_dat_i[12]
+ wb_openram_wrapper/wbs_b_dat_i[13] wb_openram_wrapper/wbs_b_dat_i[14] wb_openram_wrapper/wbs_b_dat_i[15]
+ wb_openram_wrapper/wbs_b_dat_i[16] wb_openram_wrapper/wbs_b_dat_i[17] wb_openram_wrapper/wbs_b_dat_i[18]
+ wb_openram_wrapper/wbs_b_dat_i[19] wb_openram_wrapper/wbs_b_dat_i[1] wb_openram_wrapper/wbs_b_dat_i[20]
+ wb_openram_wrapper/wbs_b_dat_i[21] wb_openram_wrapper/wbs_b_dat_i[22] wb_openram_wrapper/wbs_b_dat_i[23]
+ wb_openram_wrapper/wbs_b_dat_i[24] wb_openram_wrapper/wbs_b_dat_i[25] wb_openram_wrapper/wbs_b_dat_i[26]
+ wb_openram_wrapper/wbs_b_dat_i[27] wb_openram_wrapper/wbs_b_dat_i[28] wb_openram_wrapper/wbs_b_dat_i[29]
+ wb_openram_wrapper/wbs_b_dat_i[2] wb_openram_wrapper/wbs_b_dat_i[30] wb_openram_wrapper/wbs_b_dat_i[31]
+ wb_openram_wrapper/wbs_b_dat_i[3] wb_openram_wrapper/wbs_b_dat_i[4] wb_openram_wrapper/wbs_b_dat_i[5]
+ wb_openram_wrapper/wbs_b_dat_i[6] wb_openram_wrapper/wbs_b_dat_i[7] wb_openram_wrapper/wbs_b_dat_i[8]
+ wb_openram_wrapper/wbs_b_dat_i[9] wb_openram_wrapper/wbs_b_dat_o[0] wb_openram_wrapper/wbs_b_dat_o[10]
+ wb_openram_wrapper/wbs_b_dat_o[11] wb_openram_wrapper/wbs_b_dat_o[12] wb_openram_wrapper/wbs_b_dat_o[13]
+ wb_openram_wrapper/wbs_b_dat_o[14] wb_openram_wrapper/wbs_b_dat_o[15] wb_openram_wrapper/wbs_b_dat_o[16]
+ wb_openram_wrapper/wbs_b_dat_o[17] wb_openram_wrapper/wbs_b_dat_o[18] wb_openram_wrapper/wbs_b_dat_o[19]
+ wb_openram_wrapper/wbs_b_dat_o[1] wb_openram_wrapper/wbs_b_dat_o[20] wb_openram_wrapper/wbs_b_dat_o[21]
+ wb_openram_wrapper/wbs_b_dat_o[22] wb_openram_wrapper/wbs_b_dat_o[23] wb_openram_wrapper/wbs_b_dat_o[24]
+ wb_openram_wrapper/wbs_b_dat_o[25] wb_openram_wrapper/wbs_b_dat_o[26] wb_openram_wrapper/wbs_b_dat_o[27]
+ wb_openram_wrapper/wbs_b_dat_o[28] wb_openram_wrapper/wbs_b_dat_o[29] wb_openram_wrapper/wbs_b_dat_o[2]
+ wb_openram_wrapper/wbs_b_dat_o[30] wb_openram_wrapper/wbs_b_dat_o[31] wb_openram_wrapper/wbs_b_dat_o[3]
+ wb_openram_wrapper/wbs_b_dat_o[4] wb_openram_wrapper/wbs_b_dat_o[5] wb_openram_wrapper/wbs_b_dat_o[6]
+ wb_openram_wrapper/wbs_b_dat_o[7] wb_openram_wrapper/wbs_b_dat_o[8] wb_openram_wrapper/wbs_b_dat_o[9]
+ wb_openram_wrapper/wbs_b_sel_i[0] wb_openram_wrapper/wbs_b_sel_i[1] wb_openram_wrapper/wbs_b_sel_i[2]
+ wb_openram_wrapper/wbs_b_sel_i[3] wb_openram_wrapper/wbs_b_stb_i wb_openram_wrapper/wbs_b_we_i
+ la_data_in[31] wb_openram_wrapper
Xwrapped_ppm_decoder_3 la_data_in[3] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] vccd1 vssd1 wb_clk_i wrapped_ppm_decoder
Xwrapped_function_generator_0 la_data_in[0] io_in[0] io_in[10] io_in[11] io_in[12]
+ io_in[13] io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20]
+ io_in[21] io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28]
+ io_in[29] io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36]
+ io_in[37] io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0]
+ io_oeb[10] io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17]
+ io_oeb[18] io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24]
+ io_oeb[25] io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31]
+ io_oeb[32] io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4]
+ io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11]
+ io_out[12] io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19]
+ io_out[1] io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26]
+ io_out[27] io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33]
+ io_out[34] io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6]
+ io_out[7] io_out[8] io_out[9] wb_openram_wrapper/wbs_b_ack_o wb_openram_wrapper/wbs_b_adr_i[0]
+ wb_openram_wrapper/wbs_b_adr_i[1] wb_openram_wrapper/wbs_b_adr_i[2] wb_openram_wrapper/wbs_b_adr_i[3]
+ wb_openram_wrapper/wbs_b_adr_i[4] wb_openram_wrapper/wbs_b_adr_i[5] wb_openram_wrapper/wbs_b_adr_i[6]
+ wb_openram_wrapper/wbs_b_adr_i[7] wb_openram_wrapper/wbs_b_adr_i[8] wb_openram_wrapper/wbs_b_adr_i[9]
+ wb_openram_wrapper/wb_b_clk_i wb_openram_wrapper/wbs_b_cyc_i wb_openram_wrapper/wbs_b_dat_o[0]
+ wb_openram_wrapper/wbs_b_dat_o[10] wb_openram_wrapper/wbs_b_dat_o[11] wb_openram_wrapper/wbs_b_dat_o[12]
+ wb_openram_wrapper/wbs_b_dat_o[13] wb_openram_wrapper/wbs_b_dat_o[14] wb_openram_wrapper/wbs_b_dat_o[15]
+ wb_openram_wrapper/wbs_b_dat_o[16] wb_openram_wrapper/wbs_b_dat_o[17] wb_openram_wrapper/wbs_b_dat_o[18]
+ wb_openram_wrapper/wbs_b_dat_o[19] wb_openram_wrapper/wbs_b_dat_o[1] wb_openram_wrapper/wbs_b_dat_o[20]
+ wb_openram_wrapper/wbs_b_dat_o[21] wb_openram_wrapper/wbs_b_dat_o[22] wb_openram_wrapper/wbs_b_dat_o[23]
+ wb_openram_wrapper/wbs_b_dat_o[24] wb_openram_wrapper/wbs_b_dat_o[25] wb_openram_wrapper/wbs_b_dat_o[26]
+ wb_openram_wrapper/wbs_b_dat_o[27] wb_openram_wrapper/wbs_b_dat_o[28] wb_openram_wrapper/wbs_b_dat_o[29]
+ wb_openram_wrapper/wbs_b_dat_o[2] wb_openram_wrapper/wbs_b_dat_o[30] wb_openram_wrapper/wbs_b_dat_o[31]
+ wb_openram_wrapper/wbs_b_dat_o[3] wb_openram_wrapper/wbs_b_dat_o[4] wb_openram_wrapper/wbs_b_dat_o[5]
+ wb_openram_wrapper/wbs_b_dat_o[6] wb_openram_wrapper/wbs_b_dat_o[7] wb_openram_wrapper/wbs_b_dat_o[8]
+ wb_openram_wrapper/wbs_b_dat_o[9] wb_openram_wrapper/wbs_b_dat_i[0] wb_openram_wrapper/wbs_b_dat_i[10]
+ wb_openram_wrapper/wbs_b_dat_i[11] wb_openram_wrapper/wbs_b_dat_i[12] wb_openram_wrapper/wbs_b_dat_i[13]
+ wb_openram_wrapper/wbs_b_dat_i[14] wb_openram_wrapper/wbs_b_dat_i[15] wb_openram_wrapper/wbs_b_dat_i[16]
+ wb_openram_wrapper/wbs_b_dat_i[17] wb_openram_wrapper/wbs_b_dat_i[18] wb_openram_wrapper/wbs_b_dat_i[19]
+ wb_openram_wrapper/wbs_b_dat_i[1] wb_openram_wrapper/wbs_b_dat_i[20] wb_openram_wrapper/wbs_b_dat_i[21]
+ wb_openram_wrapper/wbs_b_dat_i[22] wb_openram_wrapper/wbs_b_dat_i[23] wb_openram_wrapper/wbs_b_dat_i[24]
+ wb_openram_wrapper/wbs_b_dat_i[25] wb_openram_wrapper/wbs_b_dat_i[26] wb_openram_wrapper/wbs_b_dat_i[27]
+ wb_openram_wrapper/wbs_b_dat_i[28] wb_openram_wrapper/wbs_b_dat_i[29] wb_openram_wrapper/wbs_b_dat_i[2]
+ wb_openram_wrapper/wbs_b_dat_i[30] wb_openram_wrapper/wbs_b_dat_i[31] wb_openram_wrapper/wbs_b_dat_i[3]
+ wb_openram_wrapper/wbs_b_dat_i[4] wb_openram_wrapper/wbs_b_dat_i[5] wb_openram_wrapper/wbs_b_dat_i[6]
+ wb_openram_wrapper/wbs_b_dat_i[7] wb_openram_wrapper/wbs_b_dat_i[8] wb_openram_wrapper/wbs_b_dat_i[9]
+ wb_openram_wrapper/wb_b_rst_i wb_openram_wrapper/wbs_b_sel_i[0] wb_openram_wrapper/wbs_b_sel_i[1]
+ wb_openram_wrapper/wbs_b_sel_i[2] wb_openram_wrapper/wbs_b_sel_i[3] wb_openram_wrapper/wbs_b_stb_i
+ wb_openram_wrapper/wbs_b_we_i vccd1 vssd1 wb_clk_i wb_rst_i wrapped_spell_1/wbs_ack_o
+ wrapped_spell_1/wbs_adr_i[0] wrapped_spell_1/wbs_adr_i[10] wrapped_spell_1/wbs_adr_i[11]
+ wrapped_spell_1/wbs_adr_i[12] wrapped_spell_1/wbs_adr_i[13] wrapped_spell_1/wbs_adr_i[14]
+ wrapped_spell_1/wbs_adr_i[15] wrapped_spell_1/wbs_adr_i[16] wrapped_spell_1/wbs_adr_i[17]
+ wrapped_spell_1/wbs_adr_i[18] wrapped_spell_1/wbs_adr_i[19] wrapped_spell_1/wbs_adr_i[1]
+ wrapped_spell_1/wbs_adr_i[20] wrapped_spell_1/wbs_adr_i[21] wrapped_spell_1/wbs_adr_i[22]
+ wrapped_spell_1/wbs_adr_i[23] wrapped_spell_1/wbs_adr_i[24] wrapped_spell_1/wbs_adr_i[25]
+ wrapped_spell_1/wbs_adr_i[26] wrapped_spell_1/wbs_adr_i[27] wrapped_spell_1/wbs_adr_i[28]
+ wrapped_spell_1/wbs_adr_i[29] wrapped_spell_1/wbs_adr_i[2] wrapped_spell_1/wbs_adr_i[30]
+ wrapped_spell_1/wbs_adr_i[31] wrapped_spell_1/wbs_adr_i[3] wrapped_spell_1/wbs_adr_i[4]
+ wrapped_spell_1/wbs_adr_i[5] wrapped_spell_1/wbs_adr_i[6] wrapped_spell_1/wbs_adr_i[7]
+ wrapped_spell_1/wbs_adr_i[8] wrapped_spell_1/wbs_adr_i[9] wrapped_spell_1/wbs_cyc_i
+ wrapped_spell_1/wbs_dat_i[0] wrapped_spell_1/wbs_dat_i[10] wrapped_spell_1/wbs_dat_i[11]
+ wrapped_spell_1/wbs_dat_i[12] wrapped_spell_1/wbs_dat_i[13] wrapped_spell_1/wbs_dat_i[14]
+ wrapped_spell_1/wbs_dat_i[15] wrapped_spell_1/wbs_dat_i[16] wrapped_spell_1/wbs_dat_i[17]
+ wrapped_spell_1/wbs_dat_i[18] wrapped_spell_1/wbs_dat_i[19] wrapped_spell_1/wbs_dat_i[1]
+ wrapped_spell_1/wbs_dat_i[20] wrapped_spell_1/wbs_dat_i[21] wrapped_spell_1/wbs_dat_i[22]
+ wrapped_spell_1/wbs_dat_i[23] wrapped_spell_1/wbs_dat_i[24] wrapped_spell_1/wbs_dat_i[25]
+ wrapped_spell_1/wbs_dat_i[26] wrapped_spell_1/wbs_dat_i[27] wrapped_spell_1/wbs_dat_i[28]
+ wrapped_spell_1/wbs_dat_i[29] wrapped_spell_1/wbs_dat_i[2] wrapped_spell_1/wbs_dat_i[30]
+ wrapped_spell_1/wbs_dat_i[31] wrapped_spell_1/wbs_dat_i[3] wrapped_spell_1/wbs_dat_i[4]
+ wrapped_spell_1/wbs_dat_i[5] wrapped_spell_1/wbs_dat_i[6] wrapped_spell_1/wbs_dat_i[7]
+ wrapped_spell_1/wbs_dat_i[8] wrapped_spell_1/wbs_dat_i[9] wrapped_spell_1/wbs_dat_o[0]
+ wrapped_spell_1/wbs_dat_o[10] wrapped_spell_1/wbs_dat_o[11] wrapped_spell_1/wbs_dat_o[12]
+ wrapped_spell_1/wbs_dat_o[13] wrapped_spell_1/wbs_dat_o[14] wrapped_spell_1/wbs_dat_o[15]
+ wrapped_spell_1/wbs_dat_o[16] wrapped_spell_1/wbs_dat_o[17] wrapped_spell_1/wbs_dat_o[18]
+ wrapped_spell_1/wbs_dat_o[19] wrapped_spell_1/wbs_dat_o[1] wrapped_spell_1/wbs_dat_o[20]
+ wrapped_spell_1/wbs_dat_o[21] wrapped_spell_1/wbs_dat_o[22] wrapped_spell_1/wbs_dat_o[23]
+ wrapped_spell_1/wbs_dat_o[24] wrapped_spell_1/wbs_dat_o[25] wrapped_spell_1/wbs_dat_o[26]
+ wrapped_spell_1/wbs_dat_o[27] wrapped_spell_1/wbs_dat_o[28] wrapped_spell_1/wbs_dat_o[29]
+ wrapped_spell_1/wbs_dat_o[2] wrapped_spell_1/wbs_dat_o[30] wrapped_spell_1/wbs_dat_o[31]
+ wrapped_spell_1/wbs_dat_o[3] wrapped_spell_1/wbs_dat_o[4] wrapped_spell_1/wbs_dat_o[5]
+ wrapped_spell_1/wbs_dat_o[6] wrapped_spell_1/wbs_dat_o[7] wrapped_spell_1/wbs_dat_o[8]
+ wrapped_spell_1/wbs_dat_o[9] wrapped_spell_1/wbs_sel_i[0] wrapped_spell_1/wbs_sel_i[1]
+ wrapped_spell_1/wbs_sel_i[2] wrapped_spell_1/wbs_sel_i[3] wrapped_spell_1/wbs_stb_i
+ wrapped_spell_1/wbs_we_i wrapped_function_generator
Xwrapped_spell_1 la_data_in[1] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[32] la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46]
+ la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[50] la_data_in[51] la_data_in[33]
+ la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57]
+ la_data_in[58] la_data_in[59] la_data_in[60] la_data_in[61] la_data_in[34] la_data_in[62]
+ la_data_in[63] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39]
+ la_data_in[40] la_data_in[41] la_data_out[32] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[50] la_data_out[51] la_data_out[33] la_data_out[52] la_data_out[53]
+ la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58]
+ la_data_out[59] la_data_out[60] la_data_out[61] la_data_out[34] la_data_out[62]
+ la_data_out[63] la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38]
+ la_data_out[39] la_data_out[40] la_data_out[41] la_oenb[32] la_oenb[42] la_oenb[43]
+ la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[50]
+ la_oenb[51] la_oenb[33] la_oenb[52] la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56]
+ la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[60] la_oenb[61] la_oenb[34] la_oenb[62]
+ la_oenb[63] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[40]
+ la_oenb[41] wb_openram_wrapper/wbs_b_ack_o wb_openram_wrapper/wbs_b_adr_i[0] wb_openram_wrapper/wbs_b_adr_i[1]
+ wb_openram_wrapper/wbs_b_adr_i[2] wb_openram_wrapper/wbs_b_adr_i[3] wb_openram_wrapper/wbs_b_adr_i[4]
+ wb_openram_wrapper/wbs_b_adr_i[5] wb_openram_wrapper/wbs_b_adr_i[6] wb_openram_wrapper/wbs_b_adr_i[7]
+ wb_openram_wrapper/wbs_b_adr_i[8] wb_openram_wrapper/wbs_b_adr_i[9] wb_openram_wrapper/wb_b_clk_i
+ wb_openram_wrapper/wbs_b_cyc_i wb_openram_wrapper/wbs_b_dat_o[0] wb_openram_wrapper/wbs_b_dat_o[10]
+ wb_openram_wrapper/wbs_b_dat_o[11] wb_openram_wrapper/wbs_b_dat_o[12] wb_openram_wrapper/wbs_b_dat_o[13]
+ wb_openram_wrapper/wbs_b_dat_o[14] wb_openram_wrapper/wbs_b_dat_o[15] wb_openram_wrapper/wbs_b_dat_o[16]
+ wb_openram_wrapper/wbs_b_dat_o[17] wb_openram_wrapper/wbs_b_dat_o[18] wb_openram_wrapper/wbs_b_dat_o[19]
+ wb_openram_wrapper/wbs_b_dat_o[1] wb_openram_wrapper/wbs_b_dat_o[20] wb_openram_wrapper/wbs_b_dat_o[21]
+ wb_openram_wrapper/wbs_b_dat_o[22] wb_openram_wrapper/wbs_b_dat_o[23] wb_openram_wrapper/wbs_b_dat_o[24]
+ wb_openram_wrapper/wbs_b_dat_o[25] wb_openram_wrapper/wbs_b_dat_o[26] wb_openram_wrapper/wbs_b_dat_o[27]
+ wb_openram_wrapper/wbs_b_dat_o[28] wb_openram_wrapper/wbs_b_dat_o[29] wb_openram_wrapper/wbs_b_dat_o[2]
+ wb_openram_wrapper/wbs_b_dat_o[30] wb_openram_wrapper/wbs_b_dat_o[31] wb_openram_wrapper/wbs_b_dat_o[3]
+ wb_openram_wrapper/wbs_b_dat_o[4] wb_openram_wrapper/wbs_b_dat_o[5] wb_openram_wrapper/wbs_b_dat_o[6]
+ wb_openram_wrapper/wbs_b_dat_o[7] wb_openram_wrapper/wbs_b_dat_o[8] wb_openram_wrapper/wbs_b_dat_o[9]
+ wb_openram_wrapper/wbs_b_dat_i[0] wb_openram_wrapper/wbs_b_dat_i[10] wb_openram_wrapper/wbs_b_dat_i[11]
+ wb_openram_wrapper/wbs_b_dat_i[12] wb_openram_wrapper/wbs_b_dat_i[13] wb_openram_wrapper/wbs_b_dat_i[14]
+ wb_openram_wrapper/wbs_b_dat_i[15] wb_openram_wrapper/wbs_b_dat_i[16] wb_openram_wrapper/wbs_b_dat_i[17]
+ wb_openram_wrapper/wbs_b_dat_i[18] wb_openram_wrapper/wbs_b_dat_i[19] wb_openram_wrapper/wbs_b_dat_i[1]
+ wb_openram_wrapper/wbs_b_dat_i[20] wb_openram_wrapper/wbs_b_dat_i[21] wb_openram_wrapper/wbs_b_dat_i[22]
+ wb_openram_wrapper/wbs_b_dat_i[23] wb_openram_wrapper/wbs_b_dat_i[24] wb_openram_wrapper/wbs_b_dat_i[25]
+ wb_openram_wrapper/wbs_b_dat_i[26] wb_openram_wrapper/wbs_b_dat_i[27] wb_openram_wrapper/wbs_b_dat_i[28]
+ wb_openram_wrapper/wbs_b_dat_i[29] wb_openram_wrapper/wbs_b_dat_i[2] wb_openram_wrapper/wbs_b_dat_i[30]
+ wb_openram_wrapper/wbs_b_dat_i[31] wb_openram_wrapper/wbs_b_dat_i[3] wb_openram_wrapper/wbs_b_dat_i[4]
+ wb_openram_wrapper/wbs_b_dat_i[5] wb_openram_wrapper/wbs_b_dat_i[6] wb_openram_wrapper/wbs_b_dat_i[7]
+ wb_openram_wrapper/wbs_b_dat_i[8] wb_openram_wrapper/wbs_b_dat_i[9] wb_openram_wrapper/wb_b_rst_i
+ wb_openram_wrapper/wbs_b_sel_i[0] wb_openram_wrapper/wbs_b_sel_i[1] wb_openram_wrapper/wbs_b_sel_i[2]
+ wb_openram_wrapper/wbs_b_sel_i[3] wb_openram_wrapper/wbs_b_stb_i wb_openram_wrapper/wbs_b_we_i
+ user_irq[0] user_irq[1] user_irq[2] vccd1 vssd1 wb_clk_i wb_rst_i wrapped_spell_1/wbs_ack_o
+ wrapped_spell_1/wbs_adr_i[0] wrapped_spell_1/wbs_adr_i[10] wrapped_spell_1/wbs_adr_i[11]
+ wrapped_spell_1/wbs_adr_i[12] wrapped_spell_1/wbs_adr_i[13] wrapped_spell_1/wbs_adr_i[14]
+ wrapped_spell_1/wbs_adr_i[15] wrapped_spell_1/wbs_adr_i[16] wrapped_spell_1/wbs_adr_i[17]
+ wrapped_spell_1/wbs_adr_i[18] wrapped_spell_1/wbs_adr_i[19] wrapped_spell_1/wbs_adr_i[1]
+ wrapped_spell_1/wbs_adr_i[20] wrapped_spell_1/wbs_adr_i[21] wrapped_spell_1/wbs_adr_i[22]
+ wrapped_spell_1/wbs_adr_i[23] wrapped_spell_1/wbs_adr_i[24] wrapped_spell_1/wbs_adr_i[25]
+ wrapped_spell_1/wbs_adr_i[26] wrapped_spell_1/wbs_adr_i[27] wrapped_spell_1/wbs_adr_i[28]
+ wrapped_spell_1/wbs_adr_i[29] wrapped_spell_1/wbs_adr_i[2] wrapped_spell_1/wbs_adr_i[30]
+ wrapped_spell_1/wbs_adr_i[31] wrapped_spell_1/wbs_adr_i[3] wrapped_spell_1/wbs_adr_i[4]
+ wrapped_spell_1/wbs_adr_i[5] wrapped_spell_1/wbs_adr_i[6] wrapped_spell_1/wbs_adr_i[7]
+ wrapped_spell_1/wbs_adr_i[8] wrapped_spell_1/wbs_adr_i[9] wrapped_spell_1/wbs_cyc_i
+ wrapped_spell_1/wbs_dat_i[0] wrapped_spell_1/wbs_dat_i[10] wrapped_spell_1/wbs_dat_i[11]
+ wrapped_spell_1/wbs_dat_i[12] wrapped_spell_1/wbs_dat_i[13] wrapped_spell_1/wbs_dat_i[14]
+ wrapped_spell_1/wbs_dat_i[15] wrapped_spell_1/wbs_dat_i[16] wrapped_spell_1/wbs_dat_i[17]
+ wrapped_spell_1/wbs_dat_i[18] wrapped_spell_1/wbs_dat_i[19] wrapped_spell_1/wbs_dat_i[1]
+ wrapped_spell_1/wbs_dat_i[20] wrapped_spell_1/wbs_dat_i[21] wrapped_spell_1/wbs_dat_i[22]
+ wrapped_spell_1/wbs_dat_i[23] wrapped_spell_1/wbs_dat_i[24] wrapped_spell_1/wbs_dat_i[25]
+ wrapped_spell_1/wbs_dat_i[26] wrapped_spell_1/wbs_dat_i[27] wrapped_spell_1/wbs_dat_i[28]
+ wrapped_spell_1/wbs_dat_i[29] wrapped_spell_1/wbs_dat_i[2] wrapped_spell_1/wbs_dat_i[30]
+ wrapped_spell_1/wbs_dat_i[31] wrapped_spell_1/wbs_dat_i[3] wrapped_spell_1/wbs_dat_i[4]
+ wrapped_spell_1/wbs_dat_i[5] wrapped_spell_1/wbs_dat_i[6] wrapped_spell_1/wbs_dat_i[7]
+ wrapped_spell_1/wbs_dat_i[8] wrapped_spell_1/wbs_dat_i[9] wrapped_spell_1/wbs_dat_o[0]
+ wrapped_spell_1/wbs_dat_o[10] wrapped_spell_1/wbs_dat_o[11] wrapped_spell_1/wbs_dat_o[12]
+ wrapped_spell_1/wbs_dat_o[13] wrapped_spell_1/wbs_dat_o[14] wrapped_spell_1/wbs_dat_o[15]
+ wrapped_spell_1/wbs_dat_o[16] wrapped_spell_1/wbs_dat_o[17] wrapped_spell_1/wbs_dat_o[18]
+ wrapped_spell_1/wbs_dat_o[19] wrapped_spell_1/wbs_dat_o[1] wrapped_spell_1/wbs_dat_o[20]
+ wrapped_spell_1/wbs_dat_o[21] wrapped_spell_1/wbs_dat_o[22] wrapped_spell_1/wbs_dat_o[23]
+ wrapped_spell_1/wbs_dat_o[24] wrapped_spell_1/wbs_dat_o[25] wrapped_spell_1/wbs_dat_o[26]
+ wrapped_spell_1/wbs_dat_o[27] wrapped_spell_1/wbs_dat_o[28] wrapped_spell_1/wbs_dat_o[29]
+ wrapped_spell_1/wbs_dat_o[2] wrapped_spell_1/wbs_dat_o[30] wrapped_spell_1/wbs_dat_o[31]
+ wrapped_spell_1/wbs_dat_o[3] wrapped_spell_1/wbs_dat_o[4] wrapped_spell_1/wbs_dat_o[5]
+ wrapped_spell_1/wbs_dat_o[6] wrapped_spell_1/wbs_dat_o[7] wrapped_spell_1/wbs_dat_o[8]
+ wrapped_spell_1/wbs_dat_o[9] wrapped_spell_1/wbs_sel_i[0] wrapped_spell_1/wbs_sel_i[1]
+ wrapped_spell_1/wbs_sel_i[2] wrapped_spell_1/wbs_sel_i[3] wrapped_spell_1/wbs_stb_i
+ wrapped_spell_1/wbs_we_i wrapped_spell
Xwrapped_bin_mult_7 la_data_in[7] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] vccd1 vssd1 wb_clk_i wb_rst_i wrapped_spell_1/wbs_ack_o wrapped_spell_1/wbs_adr_i[0]
+ wrapped_spell_1/wbs_adr_i[10] wrapped_spell_1/wbs_adr_i[11] wrapped_spell_1/wbs_adr_i[12]
+ wrapped_spell_1/wbs_adr_i[13] wrapped_spell_1/wbs_adr_i[14] wrapped_spell_1/wbs_adr_i[15]
+ wrapped_spell_1/wbs_adr_i[16] wrapped_spell_1/wbs_adr_i[17] wrapped_spell_1/wbs_adr_i[18]
+ wrapped_spell_1/wbs_adr_i[19] wrapped_spell_1/wbs_adr_i[1] wrapped_spell_1/wbs_adr_i[20]
+ wrapped_spell_1/wbs_adr_i[21] wrapped_spell_1/wbs_adr_i[22] wrapped_spell_1/wbs_adr_i[23]
+ wrapped_spell_1/wbs_adr_i[24] wrapped_spell_1/wbs_adr_i[25] wrapped_spell_1/wbs_adr_i[26]
+ wrapped_spell_1/wbs_adr_i[27] wrapped_spell_1/wbs_adr_i[28] wrapped_spell_1/wbs_adr_i[29]
+ wrapped_spell_1/wbs_adr_i[2] wrapped_spell_1/wbs_adr_i[30] wrapped_spell_1/wbs_adr_i[31]
+ wrapped_spell_1/wbs_adr_i[3] wrapped_spell_1/wbs_adr_i[4] wrapped_spell_1/wbs_adr_i[5]
+ wrapped_spell_1/wbs_adr_i[6] wrapped_spell_1/wbs_adr_i[7] wrapped_spell_1/wbs_adr_i[8]
+ wrapped_spell_1/wbs_adr_i[9] wrapped_spell_1/wbs_cyc_i wrapped_spell_1/wbs_dat_i[0]
+ wrapped_spell_1/wbs_dat_i[10] wrapped_spell_1/wbs_dat_i[11] wrapped_spell_1/wbs_dat_i[12]
+ wrapped_spell_1/wbs_dat_i[13] wrapped_spell_1/wbs_dat_i[14] wrapped_spell_1/wbs_dat_i[15]
+ wrapped_spell_1/wbs_dat_i[16] wrapped_spell_1/wbs_dat_i[17] wrapped_spell_1/wbs_dat_i[18]
+ wrapped_spell_1/wbs_dat_i[19] wrapped_spell_1/wbs_dat_i[1] wrapped_spell_1/wbs_dat_i[20]
+ wrapped_spell_1/wbs_dat_i[21] wrapped_spell_1/wbs_dat_i[22] wrapped_spell_1/wbs_dat_i[23]
+ wrapped_spell_1/wbs_dat_i[24] wrapped_spell_1/wbs_dat_i[25] wrapped_spell_1/wbs_dat_i[26]
+ wrapped_spell_1/wbs_dat_i[27] wrapped_spell_1/wbs_dat_i[28] wrapped_spell_1/wbs_dat_i[29]
+ wrapped_spell_1/wbs_dat_i[2] wrapped_spell_1/wbs_dat_i[30] wrapped_spell_1/wbs_dat_i[31]
+ wrapped_spell_1/wbs_dat_i[3] wrapped_spell_1/wbs_dat_i[4] wrapped_spell_1/wbs_dat_i[5]
+ wrapped_spell_1/wbs_dat_i[6] wrapped_spell_1/wbs_dat_i[7] wrapped_spell_1/wbs_dat_i[8]
+ wrapped_spell_1/wbs_dat_i[9] wrapped_spell_1/wbs_dat_o[0] wrapped_spell_1/wbs_dat_o[10]
+ wrapped_spell_1/wbs_dat_o[11] wrapped_spell_1/wbs_dat_o[12] wrapped_spell_1/wbs_dat_o[13]
+ wrapped_spell_1/wbs_dat_o[14] wrapped_spell_1/wbs_dat_o[15] wrapped_spell_1/wbs_dat_o[16]
+ wrapped_spell_1/wbs_dat_o[17] wrapped_spell_1/wbs_dat_o[18] wrapped_spell_1/wbs_dat_o[19]
+ wrapped_spell_1/wbs_dat_o[1] wrapped_spell_1/wbs_dat_o[20] wrapped_spell_1/wbs_dat_o[21]
+ wrapped_spell_1/wbs_dat_o[22] wrapped_spell_1/wbs_dat_o[23] wrapped_spell_1/wbs_dat_o[24]
+ wrapped_spell_1/wbs_dat_o[25] wrapped_spell_1/wbs_dat_o[26] wrapped_spell_1/wbs_dat_o[27]
+ wrapped_spell_1/wbs_dat_o[28] wrapped_spell_1/wbs_dat_o[29] wrapped_spell_1/wbs_dat_o[2]
+ wrapped_spell_1/wbs_dat_o[30] wrapped_spell_1/wbs_dat_o[31] wrapped_spell_1/wbs_dat_o[3]
+ wrapped_spell_1/wbs_dat_o[4] wrapped_spell_1/wbs_dat_o[5] wrapped_spell_1/wbs_dat_o[6]
+ wrapped_spell_1/wbs_dat_o[7] wrapped_spell_1/wbs_dat_o[8] wrapped_spell_1/wbs_dat_o[9]
+ wrapped_spell_1/wbs_sel_i[0] wrapped_spell_1/wbs_sel_i[1] wrapped_spell_1/wbs_sel_i[2]
+ wrapped_spell_1/wbs_sel_i[3] wrapped_spell_1/wbs_stb_i wrapped_spell_1/wbs_we_i
+ wrapped_bin_mult
Xwrapped_asic_watch_8 la_data_in[8] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29]
+ io_in[2] io_in[30] io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37]
+ io_in[3] io_in[4] io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[27] io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32]
+ io_oeb[33] io_oeb[34] io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5]
+ io_oeb[6] io_oeb[7] io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12]
+ io_out[13] io_out[14] io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1]
+ io_out[20] io_out[21] io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27]
+ io_out[28] io_out[29] io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34]
+ io_out[35] io_out[36] io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7]
+ io_out[8] io_out[9] la_data_in[32] la_data_in[42] la_data_in[43] la_data_in[44]
+ la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[50]
+ la_data_in[51] la_data_in[33] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55]
+ la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[60] la_data_in[61]
+ la_data_in[34] la_data_in[62] la_data_in[63] la_data_in[35] la_data_in[36] la_data_in[37]
+ la_data_in[38] la_data_in[39] la_data_in[40] la_data_in[41] la_data_out[32] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[50] la_data_out[51] la_data_out[33]
+ la_data_out[52] la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56]
+ la_data_out[57] la_data_out[58] la_data_out[59] la_data_out[60] la_data_out[61]
+ la_data_out[34] la_data_out[62] la_data_out[63] la_data_out[35] la_data_out[36]
+ la_data_out[37] la_data_out[38] la_data_out[39] la_data_out[40] la_data_out[41]
+ la_oenb[32] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46] la_oenb[47]
+ la_oenb[48] la_oenb[49] la_oenb[50] la_oenb[51] la_oenb[33] la_oenb[52] la_oenb[53]
+ la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59] la_oenb[60]
+ la_oenb[61] la_oenb[34] la_oenb[62] la_oenb[63] la_oenb[35] la_oenb[36] la_oenb[37]
+ la_oenb[38] la_oenb[39] la_oenb[40] la_oenb[41] vccd1 vssd1 wb_clk_i wb_rst_i wrapped_spell_1/wbs_ack_o
+ wrapped_spell_1/wbs_adr_i[0] wrapped_spell_1/wbs_adr_i[10] wrapped_spell_1/wbs_adr_i[11]
+ wrapped_spell_1/wbs_adr_i[12] wrapped_spell_1/wbs_adr_i[13] wrapped_spell_1/wbs_adr_i[14]
+ wrapped_spell_1/wbs_adr_i[15] wrapped_spell_1/wbs_adr_i[16] wrapped_spell_1/wbs_adr_i[17]
+ wrapped_spell_1/wbs_adr_i[18] wrapped_spell_1/wbs_adr_i[19] wrapped_spell_1/wbs_adr_i[1]
+ wrapped_spell_1/wbs_adr_i[20] wrapped_spell_1/wbs_adr_i[21] wrapped_spell_1/wbs_adr_i[22]
+ wrapped_spell_1/wbs_adr_i[23] wrapped_spell_1/wbs_adr_i[24] wrapped_spell_1/wbs_adr_i[25]
+ wrapped_spell_1/wbs_adr_i[26] wrapped_spell_1/wbs_adr_i[27] wrapped_spell_1/wbs_adr_i[28]
+ wrapped_spell_1/wbs_adr_i[29] wrapped_spell_1/wbs_adr_i[2] wrapped_spell_1/wbs_adr_i[30]
+ wrapped_spell_1/wbs_adr_i[31] wrapped_spell_1/wbs_adr_i[3] wrapped_spell_1/wbs_adr_i[4]
+ wrapped_spell_1/wbs_adr_i[5] wrapped_spell_1/wbs_adr_i[6] wrapped_spell_1/wbs_adr_i[7]
+ wrapped_spell_1/wbs_adr_i[8] wrapped_spell_1/wbs_adr_i[9] wrapped_spell_1/wbs_cyc_i
+ wrapped_spell_1/wbs_dat_i[0] wrapped_spell_1/wbs_dat_i[10] wrapped_spell_1/wbs_dat_i[11]
+ wrapped_spell_1/wbs_dat_i[12] wrapped_spell_1/wbs_dat_i[13] wrapped_spell_1/wbs_dat_i[14]
+ wrapped_spell_1/wbs_dat_i[15] wrapped_spell_1/wbs_dat_i[16] wrapped_spell_1/wbs_dat_i[17]
+ wrapped_spell_1/wbs_dat_i[18] wrapped_spell_1/wbs_dat_i[19] wrapped_spell_1/wbs_dat_i[1]
+ wrapped_spell_1/wbs_dat_i[20] wrapped_spell_1/wbs_dat_i[21] wrapped_spell_1/wbs_dat_i[22]
+ wrapped_spell_1/wbs_dat_i[23] wrapped_spell_1/wbs_dat_i[24] wrapped_spell_1/wbs_dat_i[25]
+ wrapped_spell_1/wbs_dat_i[26] wrapped_spell_1/wbs_dat_i[27] wrapped_spell_1/wbs_dat_i[28]
+ wrapped_spell_1/wbs_dat_i[29] wrapped_spell_1/wbs_dat_i[2] wrapped_spell_1/wbs_dat_i[30]
+ wrapped_spell_1/wbs_dat_i[31] wrapped_spell_1/wbs_dat_i[3] wrapped_spell_1/wbs_dat_i[4]
+ wrapped_spell_1/wbs_dat_i[5] wrapped_spell_1/wbs_dat_i[6] wrapped_spell_1/wbs_dat_i[7]
+ wrapped_spell_1/wbs_dat_i[8] wrapped_spell_1/wbs_dat_i[9] wrapped_spell_1/wbs_dat_o[0]
+ wrapped_spell_1/wbs_dat_o[10] wrapped_spell_1/wbs_dat_o[11] wrapped_spell_1/wbs_dat_o[12]
+ wrapped_spell_1/wbs_dat_o[13] wrapped_spell_1/wbs_dat_o[14] wrapped_spell_1/wbs_dat_o[15]
+ wrapped_spell_1/wbs_dat_o[16] wrapped_spell_1/wbs_dat_o[17] wrapped_spell_1/wbs_dat_o[18]
+ wrapped_spell_1/wbs_dat_o[19] wrapped_spell_1/wbs_dat_o[1] wrapped_spell_1/wbs_dat_o[20]
+ wrapped_spell_1/wbs_dat_o[21] wrapped_spell_1/wbs_dat_o[22] wrapped_spell_1/wbs_dat_o[23]
+ wrapped_spell_1/wbs_dat_o[24] wrapped_spell_1/wbs_dat_o[25] wrapped_spell_1/wbs_dat_o[26]
+ wrapped_spell_1/wbs_dat_o[27] wrapped_spell_1/wbs_dat_o[28] wrapped_spell_1/wbs_dat_o[29]
+ wrapped_spell_1/wbs_dat_o[2] wrapped_spell_1/wbs_dat_o[30] wrapped_spell_1/wbs_dat_o[31]
+ wrapped_spell_1/wbs_dat_o[3] wrapped_spell_1/wbs_dat_o[4] wrapped_spell_1/wbs_dat_o[5]
+ wrapped_spell_1/wbs_dat_o[6] wrapped_spell_1/wbs_dat_o[7] wrapped_spell_1/wbs_dat_o[8]
+ wrapped_spell_1/wbs_dat_o[9] wrapped_spell_1/wbs_sel_i[0] wrapped_spell_1/wbs_sel_i[1]
+ wrapped_spell_1/wbs_sel_i[2] wrapped_spell_1/wbs_sel_i[3] wrapped_spell_1/wbs_stb_i
+ wrapped_spell_1/wbs_we_i wrapped_asic_watch
.ends

