magic
tech sky130A
magscale 1 2
timestamp 1640170089
<< metal1 >>
rect 122098 703604 122104 703656
rect 122156 703644 122162 703656
rect 234982 703644 234988 703656
rect 122156 703616 234988 703644
rect 122156 703604 122162 703616
rect 234982 703604 234988 703616
rect 235040 703604 235046 703656
rect 75822 703536 75828 703588
rect 75880 703576 75886 703588
rect 202598 703576 202604 703588
rect 75880 703548 202604 703576
rect 75880 703536 75886 703548
rect 202598 703536 202604 703548
rect 202656 703536 202662 703588
rect 67634 703468 67640 703520
rect 67692 703508 67698 703520
rect 267458 703508 267464 703520
rect 67692 703480 267464 703508
rect 67692 703468 67698 703480
rect 267458 703468 267464 703480
rect 267516 703468 267522 703520
rect 93762 703400 93768 703452
rect 93820 703440 93826 703452
rect 300118 703440 300124 703452
rect 93820 703412 300124 703440
rect 93820 703400 93826 703412
rect 300118 703400 300124 703412
rect 300176 703400 300182 703452
rect 59262 703332 59268 703384
rect 59320 703372 59326 703384
rect 283834 703372 283840 703384
rect 59320 703344 283840 703372
rect 59320 703332 59326 703344
rect 283834 703332 283840 703344
rect 283892 703332 283898 703384
rect 73062 703264 73068 703316
rect 73120 703304 73126 703316
rect 332502 703304 332508 703316
rect 73120 703276 332508 703304
rect 73120 703264 73126 703276
rect 332502 703264 332508 703276
rect 332560 703264 332566 703316
rect 130378 703196 130384 703248
rect 130436 703236 130442 703248
rect 413646 703236 413652 703248
rect 130436 703208 413652 703236
rect 130436 703196 130442 703208
rect 413646 703196 413652 703208
rect 413704 703196 413710 703248
rect 61838 703128 61844 703180
rect 61896 703168 61902 703180
rect 348786 703168 348792 703180
rect 61896 703140 348792 703168
rect 61896 703128 61902 703140
rect 348786 703128 348792 703140
rect 348844 703128 348850 703180
rect 101490 703060 101496 703112
rect 101548 703100 101554 703112
rect 397454 703100 397460 703112
rect 101548 703072 397460 703100
rect 101548 703060 101554 703072
rect 397454 703060 397460 703072
rect 397512 703060 397518 703112
rect 124858 702992 124864 703044
rect 124916 703032 124922 703044
rect 429838 703032 429844 703044
rect 124916 703004 429844 703032
rect 124916 702992 124922 703004
rect 429838 702992 429844 703004
rect 429896 702992 429902 703044
rect 57882 702924 57888 702976
rect 57940 702964 57946 702976
rect 364978 702964 364984 702976
rect 57940 702936 364984 702964
rect 57940 702924 57946 702936
rect 364978 702924 364984 702936
rect 365036 702924 365042 702976
rect 126238 702856 126244 702908
rect 126296 702896 126302 702908
rect 462314 702896 462320 702908
rect 126296 702868 462320 702896
rect 126296 702856 126302 702868
rect 462314 702856 462320 702868
rect 462372 702856 462378 702908
rect 71038 702788 71044 702840
rect 71096 702828 71102 702840
rect 494790 702828 494796 702840
rect 71096 702800 494796 702828
rect 71096 702788 71102 702800
rect 494790 702788 494796 702800
rect 494848 702788 494854 702840
rect 97902 702720 97908 702772
rect 97960 702760 97966 702772
rect 478506 702760 478512 702772
rect 97960 702732 478512 702760
rect 97960 702720 97966 702732
rect 478506 702720 478512 702732
rect 478564 702720 478570 702772
rect 128998 702652 129004 702704
rect 129056 702692 129062 702704
rect 543458 702692 543464 702704
rect 129056 702664 543464 702692
rect 129056 702652 129062 702664
rect 543458 702652 543464 702664
rect 543516 702652 543522 702704
rect 8110 702584 8116 702636
rect 8168 702624 8174 702636
rect 89806 702624 89812 702636
rect 8168 702596 89812 702624
rect 8168 702584 8174 702596
rect 89806 702584 89812 702596
rect 89864 702584 89870 702636
rect 94498 702584 94504 702636
rect 94556 702624 94562 702636
rect 527174 702624 527180 702636
rect 94556 702596 527180 702624
rect 94556 702584 94562 702596
rect 527174 702584 527180 702596
rect 527232 702584 527238 702636
rect 53742 702516 53748 702568
rect 53800 702556 53806 702568
rect 580258 702556 580264 702568
rect 53800 702528 580264 702556
rect 53800 702516 53806 702528
rect 580258 702516 580264 702528
rect 580316 702516 580322 702568
rect 66162 702448 66168 702500
rect 66220 702488 66226 702500
rect 559650 702488 559656 702500
rect 66220 702460 559656 702488
rect 66220 702448 66226 702460
rect 559650 702448 559656 702460
rect 559708 702448 559714 702500
rect 83458 700340 83464 700392
rect 83516 700380 83522 700392
rect 89162 700380 89168 700392
rect 83516 700352 89168 700380
rect 83516 700340 83522 700352
rect 89162 700340 89168 700352
rect 89220 700340 89226 700392
rect 40494 700272 40500 700324
rect 40552 700312 40558 700324
rect 89070 700312 89076 700324
rect 40552 700284 89076 700312
rect 40552 700272 40558 700284
rect 89070 700272 89076 700284
rect 89128 700272 89134 700324
rect 133138 700272 133144 700324
rect 133196 700312 133202 700324
rect 218974 700312 218980 700324
rect 133196 700284 218980 700312
rect 133196 700272 133202 700284
rect 218974 700272 218980 700284
rect 219032 700272 219038 700324
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 25498 699700 25504 699712
rect 24360 699672 25504 699700
rect 24360 699660 24366 699672
rect 25498 699660 25504 699672
rect 25556 699660 25562 699712
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 11698 683176 11704 683188
rect 3476 683148 11704 683176
rect 3476 683136 3482 683148
rect 11698 683136 11704 683148
rect 11756 683136 11762 683188
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 14458 670732 14464 670744
rect 3568 670704 14464 670732
rect 3568 670692 3574 670704
rect 14458 670692 14464 670704
rect 14516 670692 14522 670744
rect 3418 658112 3424 658164
rect 3476 658152 3482 658164
rect 7558 658152 7564 658164
rect 3476 658124 7564 658152
rect 3476 658112 3482 658124
rect 7558 658112 7564 658124
rect 7616 658112 7622 658164
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 17218 632108 17224 632120
rect 3476 632080 17224 632108
rect 3476 632068 3482 632080
rect 17218 632068 17224 632080
rect 17276 632068 17282 632120
rect 2774 619080 2780 619132
rect 2832 619120 2838 619132
rect 4798 619120 4804 619132
rect 2832 619092 4804 619120
rect 2832 619080 2838 619092
rect 4798 619080 4804 619092
rect 4856 619080 4862 619132
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 87598 605860 87604 605872
rect 3292 605832 87604 605860
rect 3292 605820 3298 605832
rect 87598 605820 87604 605832
rect 87656 605820 87662 605872
rect 67450 599564 67456 599616
rect 67508 599604 67514 599616
rect 104894 599604 104900 599616
rect 67508 599576 104900 599604
rect 67508 599564 67514 599576
rect 104894 599564 104900 599576
rect 104952 599564 104958 599616
rect 79962 597524 79968 597576
rect 80020 597564 80026 597576
rect 106918 597564 106924 597576
rect 80020 597536 106924 597564
rect 80020 597524 80026 597536
rect 106918 597524 106924 597536
rect 106976 597524 106982 597576
rect 67542 596776 67548 596828
rect 67600 596816 67606 596828
rect 169754 596816 169760 596828
rect 67600 596788 169760 596816
rect 67600 596776 67606 596788
rect 169754 596776 169760 596788
rect 169812 596776 169818 596828
rect 25498 596096 25504 596148
rect 25556 596136 25562 596148
rect 79962 596136 79968 596148
rect 25556 596108 79968 596136
rect 25556 596096 25562 596108
rect 79962 596096 79968 596108
rect 80020 596096 80026 596148
rect 108298 595416 108304 595468
rect 108356 595456 108362 595468
rect 582742 595456 582748 595468
rect 108356 595428 582748 595456
rect 108356 595416 108362 595428
rect 582742 595416 582748 595428
rect 582800 595416 582806 595468
rect 77018 594804 77024 594856
rect 77076 594844 77082 594856
rect 101398 594844 101404 594856
rect 77076 594816 101404 594844
rect 77076 594804 77082 594816
rect 101398 594804 101404 594816
rect 101456 594804 101462 594856
rect 87598 594532 87604 594584
rect 87656 594572 87662 594584
rect 91186 594572 91192 594584
rect 87656 594544 91192 594572
rect 87656 594532 87662 594544
rect 91186 594532 91192 594544
rect 91244 594532 91250 594584
rect 83458 593376 83464 593428
rect 83516 593416 83522 593428
rect 110414 593416 110420 593428
rect 83516 593388 110420 593416
rect 83516 593376 83522 593388
rect 110414 593376 110420 593388
rect 110472 593376 110478 593428
rect 7558 592628 7564 592680
rect 7616 592668 7622 592680
rect 69014 592668 69020 592680
rect 7616 592640 69020 592668
rect 7616 592628 7622 592640
rect 69014 592628 69020 592640
rect 69072 592628 69078 592680
rect 75730 592084 75736 592136
rect 75788 592124 75794 592136
rect 96614 592124 96620 592136
rect 75788 592096 96620 592124
rect 75788 592084 75794 592096
rect 96614 592084 96620 592096
rect 96672 592084 96678 592136
rect 79778 592016 79784 592068
rect 79836 592056 79842 592068
rect 105538 592056 105544 592068
rect 79836 592028 105544 592056
rect 79836 592016 79842 592028
rect 105538 592016 105544 592028
rect 105596 592016 105602 592068
rect 78398 590792 78404 590844
rect 78456 590832 78462 590844
rect 103514 590832 103520 590844
rect 78456 590804 103520 590832
rect 78456 590792 78462 590804
rect 103514 590792 103520 590804
rect 103572 590792 103578 590844
rect 61930 590656 61936 590708
rect 61988 590696 61994 590708
rect 70854 590696 70860 590708
rect 61988 590668 70860 590696
rect 61988 590656 61994 590668
rect 70854 590656 70860 590668
rect 70912 590656 70918 590708
rect 71682 590656 71688 590708
rect 71740 590696 71746 590708
rect 74994 590696 75000 590708
rect 71740 590668 75000 590696
rect 71740 590656 71746 590668
rect 74994 590656 75000 590668
rect 75052 590696 75058 590708
rect 75730 590696 75736 590708
rect 75052 590668 75736 590696
rect 75052 590656 75058 590668
rect 75730 590656 75736 590668
rect 75788 590656 75794 590708
rect 3418 589908 3424 589960
rect 3476 589948 3482 589960
rect 71682 589948 71688 589960
rect 3476 589920 71688 589948
rect 3476 589908 3482 589920
rect 71682 589908 71688 589920
rect 71740 589908 71746 589960
rect 81342 589432 81348 589484
rect 81400 589472 81406 589484
rect 81400 589444 93854 589472
rect 81400 589432 81406 589444
rect 70302 589364 70308 589416
rect 70360 589404 70366 589416
rect 89714 589404 89720 589416
rect 70360 589376 89720 589404
rect 70360 589364 70366 589376
rect 89714 589364 89720 589376
rect 89772 589364 89778 589416
rect 93826 589336 93854 589444
rect 108298 589336 108304 589348
rect 93826 589308 108304 589336
rect 108298 589296 108304 589308
rect 108356 589296 108362 589348
rect 69474 588616 69480 588668
rect 69532 588656 69538 588668
rect 88978 588656 88984 588668
rect 69532 588628 88984 588656
rect 69532 588616 69538 588628
rect 88978 588616 88984 588628
rect 89036 588616 89042 588668
rect 85574 588548 85580 588600
rect 85632 588588 85638 588600
rect 114462 588588 114468 588600
rect 85632 588560 114468 588588
rect 85632 588548 85638 588560
rect 114462 588548 114468 588560
rect 114520 588548 114526 588600
rect 84378 588412 84384 588464
rect 84436 588412 84442 588464
rect 86218 588412 86224 588464
rect 86276 588452 86282 588464
rect 89162 588452 89168 588464
rect 86276 588424 89168 588452
rect 86276 588412 86282 588424
rect 89162 588412 89168 588424
rect 89220 588412 89226 588464
rect 63310 587868 63316 587920
rect 63368 587908 63374 587920
rect 66806 587908 66812 587920
rect 63368 587880 66812 587908
rect 63368 587868 63374 587880
rect 66806 587868 66812 587880
rect 66864 587868 66870 587920
rect 84396 587840 84424 588412
rect 92474 587840 92480 587852
rect 84396 587812 92480 587840
rect 92474 587800 92480 587812
rect 92532 587800 92538 587852
rect 114462 587800 114468 587852
rect 114520 587840 114526 587852
rect 122098 587840 122104 587852
rect 114520 587812 122104 587840
rect 114520 587800 114526 587812
rect 122098 587800 122104 587812
rect 122156 587800 122162 587852
rect 59170 586508 59176 586560
rect 59228 586548 59234 586560
rect 66254 586548 66260 586560
rect 59228 586520 66260 586548
rect 59228 586508 59234 586520
rect 66254 586508 66260 586520
rect 66312 586508 66318 586560
rect 89162 585760 89168 585812
rect 89220 585800 89226 585812
rect 116578 585800 116584 585812
rect 89220 585772 116584 585800
rect 89220 585760 89226 585772
rect 116578 585760 116584 585772
rect 116636 585760 116642 585812
rect 50890 585148 50896 585200
rect 50948 585188 50954 585200
rect 67726 585188 67732 585200
rect 50948 585160 67732 585188
rect 50948 585148 50954 585160
rect 67726 585148 67732 585160
rect 67784 585148 67790 585200
rect 91922 584400 91928 584452
rect 91980 584440 91986 584452
rect 93762 584440 93768 584452
rect 91980 584412 93768 584440
rect 91980 584400 91986 584412
rect 93762 584400 93768 584412
rect 93820 584440 93826 584452
rect 115198 584440 115204 584452
rect 93820 584412 115204 584440
rect 93820 584400 93826 584412
rect 115198 584400 115204 584412
rect 115256 584400 115262 584452
rect 91922 583652 91928 583704
rect 91980 583692 91986 583704
rect 93762 583692 93768 583704
rect 91980 583664 93768 583692
rect 91980 583652 91986 583664
rect 93762 583652 93768 583664
rect 93820 583692 93826 583704
rect 94498 583692 94504 583704
rect 93820 583664 94504 583692
rect 93820 583652 93826 583664
rect 94498 583652 94504 583664
rect 94556 583652 94562 583704
rect 48130 582360 48136 582412
rect 48188 582400 48194 582412
rect 66806 582400 66812 582412
rect 48188 582372 66812 582400
rect 48188 582360 48194 582372
rect 66806 582360 66812 582372
rect 66864 582360 66870 582412
rect 64690 581000 64696 581052
rect 64748 581040 64754 581052
rect 66990 581040 66996 581052
rect 64748 581012 66996 581040
rect 64748 581000 64754 581012
rect 66990 581000 66996 581012
rect 67048 581000 67054 581052
rect 91094 581000 91100 581052
rect 91152 581040 91158 581052
rect 102778 581040 102784 581052
rect 91152 581012 102784 581040
rect 91152 581000 91158 581012
rect 102778 581000 102784 581012
rect 102836 581000 102842 581052
rect 91094 578212 91100 578264
rect 91152 578252 91158 578264
rect 121546 578252 121552 578264
rect 91152 578224 121552 578252
rect 91152 578212 91158 578224
rect 121546 578212 121552 578224
rect 121604 578212 121610 578264
rect 100662 577464 100668 577516
rect 100720 577504 100726 577516
rect 582466 577504 582472 577516
rect 100720 577476 582472 577504
rect 100720 577464 100726 577476
rect 582466 577464 582472 577476
rect 582524 577464 582530 577516
rect 91094 576852 91100 576904
rect 91152 576892 91158 576904
rect 100662 576892 100668 576904
rect 91152 576864 100668 576892
rect 91152 576852 91158 576864
rect 100662 576852 100668 576864
rect 100720 576852 100726 576904
rect 17218 576104 17224 576156
rect 17276 576144 17282 576156
rect 34514 576144 34520 576156
rect 17276 576116 34520 576144
rect 17276 576104 17282 576116
rect 34514 576104 34520 576116
rect 34572 576104 34578 576156
rect 91186 576104 91192 576156
rect 91244 576144 91250 576156
rect 105630 576144 105636 576156
rect 91244 576116 105636 576144
rect 91244 576104 91250 576116
rect 105630 576104 105636 576116
rect 105688 576104 105694 576156
rect 34514 575492 34520 575544
rect 34572 575532 34578 575544
rect 35802 575532 35808 575544
rect 34572 575504 35808 575532
rect 34572 575492 34578 575504
rect 35802 575492 35808 575504
rect 35860 575532 35866 575544
rect 66898 575532 66904 575544
rect 35860 575504 66904 575532
rect 35860 575492 35866 575504
rect 66898 575492 66904 575504
rect 66956 575492 66962 575544
rect 89070 575492 89076 575544
rect 89128 575532 89134 575544
rect 91278 575532 91284 575544
rect 89128 575504 91284 575532
rect 89128 575492 89134 575504
rect 91278 575492 91284 575504
rect 91336 575492 91342 575544
rect 55030 574744 55036 574796
rect 55088 574784 55094 574796
rect 67450 574784 67456 574796
rect 55088 574756 67456 574784
rect 55088 574744 55094 574756
rect 67450 574744 67456 574756
rect 67508 574744 67514 574796
rect 91922 574744 91928 574796
rect 91980 574784 91986 574796
rect 93762 574784 93768 574796
rect 91980 574756 93768 574784
rect 91980 574744 91986 574756
rect 93762 574744 93768 574756
rect 93820 574784 93826 574796
rect 101490 574784 101496 574796
rect 93820 574756 101496 574784
rect 93820 574744 93826 574756
rect 101490 574744 101496 574756
rect 101548 574744 101554 574796
rect 41322 572704 41328 572756
rect 41380 572744 41386 572756
rect 66438 572744 66444 572756
rect 41380 572716 66444 572744
rect 41380 572704 41386 572716
rect 66438 572704 66444 572716
rect 66496 572704 66502 572756
rect 91094 572704 91100 572756
rect 91152 572744 91158 572756
rect 120718 572744 120724 572756
rect 91152 572716 120724 572744
rect 91152 572704 91158 572716
rect 120718 572704 120724 572716
rect 120776 572704 120782 572756
rect 91094 571412 91100 571464
rect 91152 571452 91158 571464
rect 94498 571452 94504 571464
rect 91152 571424 94504 571452
rect 91152 571412 91158 571424
rect 94498 571412 94504 571424
rect 94556 571412 94562 571464
rect 49602 571344 49608 571396
rect 49660 571384 49666 571396
rect 66438 571384 66444 571396
rect 49660 571356 66444 571384
rect 49660 571344 49666 571356
rect 66438 571344 66444 571356
rect 66496 571344 66502 571396
rect 91186 571344 91192 571396
rect 91244 571384 91250 571396
rect 126974 571384 126980 571396
rect 91244 571356 126980 571384
rect 91244 571344 91250 571356
rect 126974 571344 126980 571356
rect 127032 571344 127038 571396
rect 91094 569916 91100 569968
rect 91152 569956 91158 569968
rect 128354 569956 128360 569968
rect 91152 569928 128360 569956
rect 91152 569916 91158 569928
rect 128354 569916 128360 569928
rect 128412 569916 128418 569968
rect 93762 569168 93768 569220
rect 93820 569208 93826 569220
rect 123478 569208 123484 569220
rect 93820 569180 123484 569208
rect 93820 569168 93826 569180
rect 123478 569168 123484 569180
rect 123536 569168 123542 569220
rect 64782 568556 64788 568608
rect 64840 568596 64846 568608
rect 66806 568596 66812 568608
rect 64840 568568 66812 568596
rect 64840 568556 64846 568568
rect 66806 568556 66812 568568
rect 66864 568556 66870 568608
rect 91278 567808 91284 567860
rect 91336 567848 91342 567860
rect 124214 567848 124220 567860
rect 91336 567820 124220 567848
rect 91336 567808 91342 567820
rect 124214 567808 124220 567820
rect 124272 567808 124278 567860
rect 57698 567196 57704 567248
rect 57756 567236 57762 567248
rect 66898 567236 66904 567248
rect 57756 567208 66904 567236
rect 57756 567196 57762 567208
rect 66898 567196 66904 567208
rect 66956 567196 66962 567248
rect 53650 566448 53656 566500
rect 53708 566488 53714 566500
rect 67542 566488 67548 566500
rect 53708 566460 67548 566488
rect 53708 566448 53714 566460
rect 67542 566448 67548 566460
rect 67600 566448 67606 566500
rect 91094 565836 91100 565888
rect 91152 565876 91158 565888
rect 101490 565876 101496 565888
rect 91152 565848 101496 565876
rect 91152 565836 91158 565848
rect 101490 565836 101496 565848
rect 101548 565836 101554 565888
rect 60642 564408 60648 564460
rect 60700 564448 60706 564460
rect 66622 564448 66628 564460
rect 60700 564420 66628 564448
rect 60700 564408 60706 564420
rect 66622 564408 66628 564420
rect 66680 564408 66686 564460
rect 91094 564408 91100 564460
rect 91152 564448 91158 564460
rect 120626 564448 120632 564460
rect 91152 564420 120632 564448
rect 91152 564408 91158 564420
rect 120626 564408 120632 564420
rect 120684 564408 120690 564460
rect 50982 564340 50988 564392
rect 51040 564380 51046 564392
rect 53742 564380 53748 564392
rect 51040 564352 53748 564380
rect 51040 564340 51046 564352
rect 53742 564340 53748 564352
rect 53800 564380 53806 564392
rect 66438 564380 66444 564392
rect 53800 564352 66444 564380
rect 53800 564340 53806 564352
rect 66438 564340 66444 564352
rect 66496 564340 66502 564392
rect 91094 563048 91100 563100
rect 91152 563088 91158 563100
rect 129734 563088 129740 563100
rect 91152 563060 129740 563088
rect 91152 563048 91158 563060
rect 129734 563048 129740 563060
rect 129792 563048 129798 563100
rect 37182 561688 37188 561740
rect 37240 561728 37246 561740
rect 66438 561728 66444 561740
rect 37240 561700 66444 561728
rect 37240 561688 37246 561700
rect 66438 561688 66444 561700
rect 66496 561688 66502 561740
rect 44082 560260 44088 560312
rect 44140 560300 44146 560312
rect 66622 560300 66628 560312
rect 44140 560272 66628 560300
rect 44140 560260 44146 560272
rect 66622 560260 66628 560272
rect 66680 560260 66686 560312
rect 56502 558900 56508 558952
rect 56560 558940 56566 558952
rect 66622 558940 66628 558952
rect 56560 558912 66628 558940
rect 56560 558900 56566 558912
rect 66622 558900 66628 558912
rect 66680 558900 66686 558952
rect 48222 557540 48228 557592
rect 48280 557580 48286 557592
rect 67634 557580 67640 557592
rect 48280 557552 67640 557580
rect 48280 557540 48286 557552
rect 67634 557540 67640 557552
rect 67692 557540 67698 557592
rect 91186 557540 91192 557592
rect 91244 557580 91250 557592
rect 125594 557580 125600 557592
rect 91244 557552 125600 557580
rect 91244 557540 91250 557552
rect 125594 557540 125600 557552
rect 125652 557540 125658 557592
rect 91186 556180 91192 556232
rect 91244 556220 91250 556232
rect 122098 556220 122104 556232
rect 91244 556192 122104 556220
rect 91244 556180 91250 556192
rect 122098 556180 122104 556192
rect 122156 556180 122162 556232
rect 58986 554752 58992 554804
rect 59044 554792 59050 554804
rect 66346 554792 66352 554804
rect 59044 554764 66352 554792
rect 59044 554752 59050 554764
rect 66346 554752 66352 554764
rect 66404 554752 66410 554804
rect 91186 554752 91192 554804
rect 91244 554792 91250 554804
rect 108942 554792 108948 554804
rect 91244 554764 108948 554792
rect 91244 554752 91250 554764
rect 108942 554752 108948 554764
rect 109000 554792 109006 554804
rect 582466 554792 582472 554804
rect 109000 554764 582472 554792
rect 109000 554752 109006 554764
rect 582466 554752 582472 554764
rect 582524 554752 582530 554804
rect 59262 554684 59268 554736
rect 59320 554724 59326 554736
rect 65518 554724 65524 554736
rect 59320 554696 65524 554724
rect 59320 554684 59326 554696
rect 65518 554684 65524 554696
rect 65576 554724 65582 554736
rect 66254 554724 66260 554736
rect 65576 554696 66260 554724
rect 65576 554684 65582 554696
rect 66254 554684 66260 554696
rect 66312 554684 66318 554736
rect 3326 553392 3332 553444
rect 3384 553432 3390 553444
rect 32398 553432 32404 553444
rect 3384 553404 32404 553432
rect 3384 553392 3390 553404
rect 32398 553392 32404 553404
rect 32456 553392 32462 553444
rect 107102 553052 107108 553104
rect 107160 553092 107166 553104
rect 109034 553092 109040 553104
rect 107160 553064 109040 553092
rect 107160 553052 107166 553064
rect 109034 553052 109040 553064
rect 109092 553052 109098 553104
rect 91186 552100 91192 552152
rect 91244 552140 91250 552152
rect 107010 552140 107016 552152
rect 91244 552112 107016 552140
rect 91244 552100 91250 552112
rect 107010 552100 107016 552112
rect 107068 552100 107074 552152
rect 91278 552032 91284 552084
rect 91336 552072 91342 552084
rect 134518 552072 134524 552084
rect 91336 552044 134524 552072
rect 91336 552032 91342 552044
rect 134518 552032 134524 552044
rect 134576 552032 134582 552084
rect 63402 549244 63408 549296
rect 63460 549284 63466 549296
rect 66530 549284 66536 549296
rect 63460 549256 66536 549284
rect 63460 549244 63466 549256
rect 66530 549244 66536 549256
rect 66588 549244 66594 549296
rect 91186 549244 91192 549296
rect 91244 549284 91250 549296
rect 104250 549284 104256 549296
rect 91244 549256 104256 549284
rect 91244 549244 91250 549256
rect 104250 549244 104256 549256
rect 104308 549244 104314 549296
rect 91830 548496 91836 548548
rect 91888 548536 91894 548548
rect 121454 548536 121460 548548
rect 91888 548508 121460 548536
rect 91888 548496 91894 548508
rect 121454 548496 121460 548508
rect 121512 548496 121518 548548
rect 62022 547884 62028 547936
rect 62080 547924 62086 547936
rect 66530 547924 66536 547936
rect 62080 547896 66536 547924
rect 62080 547884 62086 547896
rect 66530 547884 66536 547896
rect 66588 547884 66594 547936
rect 61838 547748 61844 547800
rect 61896 547788 61902 547800
rect 66806 547788 66812 547800
rect 61896 547760 66812 547788
rect 61896 547748 61902 547760
rect 66806 547748 66812 547760
rect 66864 547748 66870 547800
rect 53742 547136 53748 547188
rect 53800 547176 53806 547188
rect 61838 547176 61844 547188
rect 53800 547148 61844 547176
rect 53800 547136 53806 547148
rect 61838 547136 61844 547148
rect 61896 547136 61902 547188
rect 91278 546456 91284 546508
rect 91336 546496 91342 546508
rect 104158 546496 104164 546508
rect 91336 546468 104164 546496
rect 91336 546456 91342 546468
rect 104158 546456 104164 546468
rect 104216 546456 104222 546508
rect 57790 545708 57796 545760
rect 57848 545748 57854 545760
rect 66162 545748 66168 545760
rect 57848 545720 66168 545748
rect 57848 545708 57854 545720
rect 66162 545708 66168 545720
rect 66220 545708 66226 545760
rect 91278 545708 91284 545760
rect 91336 545748 91342 545760
rect 96430 545748 96436 545760
rect 91336 545720 96436 545748
rect 91336 545708 91342 545720
rect 96430 545708 96436 545720
rect 96488 545748 96494 545760
rect 126238 545748 126244 545760
rect 96488 545720 126244 545748
rect 96488 545708 96494 545720
rect 126238 545708 126244 545720
rect 126296 545708 126302 545760
rect 52362 545028 52368 545080
rect 52420 545068 52426 545080
rect 57882 545068 57888 545080
rect 52420 545040 57888 545068
rect 52420 545028 52426 545040
rect 57882 545028 57888 545040
rect 57940 545068 57946 545080
rect 66806 545068 66812 545080
rect 57940 545040 66812 545068
rect 57940 545028 57946 545040
rect 66806 545028 66812 545040
rect 66864 545028 66870 545080
rect 91278 544348 91284 544400
rect 91336 544388 91342 544400
rect 96522 544388 96528 544400
rect 91336 544360 96528 544388
rect 91336 544348 91342 544360
rect 96522 544348 96528 544360
rect 96580 544388 96586 544400
rect 128998 544388 129004 544400
rect 96580 544360 129004 544388
rect 96580 544348 96586 544360
rect 128998 544348 129004 544360
rect 129056 544348 129062 544400
rect 11698 542988 11704 543040
rect 11756 543028 11762 543040
rect 39942 543028 39948 543040
rect 11756 543000 39948 543028
rect 11756 542988 11762 543000
rect 39942 542988 39948 543000
rect 40000 542988 40006 543040
rect 95878 542988 95884 543040
rect 95936 543028 95942 543040
rect 117314 543028 117320 543040
rect 95936 543000 117320 543028
rect 95936 542988 95942 543000
rect 117314 542988 117320 543000
rect 117372 542988 117378 543040
rect 39942 542376 39948 542428
rect 40000 542416 40006 542428
rect 66806 542416 66812 542428
rect 40000 542388 66812 542416
rect 40000 542376 40006 542388
rect 66806 542376 66812 542388
rect 66864 542376 66870 542428
rect 91278 542376 91284 542428
rect 91336 542416 91342 542428
rect 97258 542416 97264 542428
rect 91336 542388 97264 542416
rect 91336 542376 91342 542388
rect 97258 542376 97264 542388
rect 97316 542376 97322 542428
rect 14458 541628 14464 541680
rect 14516 541668 14522 541680
rect 67082 541668 67088 541680
rect 14516 541640 67088 541668
rect 14516 541628 14522 541640
rect 67082 541628 67088 541640
rect 67140 541628 67146 541680
rect 91278 541628 91284 541680
rect 91336 541668 91342 541680
rect 136634 541668 136640 541680
rect 91336 541640 136640 541668
rect 91336 541628 91342 541640
rect 136634 541628 136640 541640
rect 136692 541628 136698 541680
rect 67542 540880 67548 540932
rect 67600 540920 67606 540932
rect 68646 540920 68652 540932
rect 67600 540892 68652 540920
rect 67600 540880 67606 540892
rect 68646 540880 68652 540892
rect 68704 540920 68710 540932
rect 582650 540920 582656 540932
rect 68704 540892 582656 540920
rect 68704 540880 68710 540892
rect 582650 540880 582656 540892
rect 582708 540880 582714 540932
rect 3418 540200 3424 540252
rect 3476 540240 3482 540252
rect 3476 540212 64874 540240
rect 3476 540200 3482 540212
rect 64846 539696 64874 540212
rect 64846 539668 69888 539696
rect 69860 539640 69888 539668
rect 91278 539656 91284 539708
rect 91336 539696 91342 539708
rect 93118 539696 93124 539708
rect 91336 539668 93124 539696
rect 91336 539656 91342 539668
rect 93118 539656 93124 539668
rect 93176 539656 93182 539708
rect 55122 539588 55128 539640
rect 55180 539628 55186 539640
rect 67542 539628 67548 539640
rect 55180 539600 67548 539628
rect 55180 539588 55186 539600
rect 67542 539588 67548 539600
rect 67600 539588 67606 539640
rect 69842 539588 69848 539640
rect 69900 539588 69906 539640
rect 67082 539452 67088 539504
rect 67140 539492 67146 539504
rect 67542 539492 67548 539504
rect 67140 539464 67548 539492
rect 67140 539452 67146 539464
rect 67542 539452 67548 539464
rect 67600 539452 67606 539504
rect 67818 538908 67824 538960
rect 67876 538948 67882 538960
rect 74718 538948 74724 538960
rect 67876 538920 74724 538948
rect 67876 538908 67882 538920
rect 74718 538908 74724 538920
rect 74776 538908 74782 538960
rect 3418 538840 3424 538892
rect 3476 538880 3482 538892
rect 89898 538880 89904 538892
rect 3476 538852 89904 538880
rect 3476 538840 3482 538852
rect 89898 538840 89904 538852
rect 89956 538840 89962 538892
rect 80330 538228 80336 538280
rect 80388 538268 80394 538280
rect 80790 538268 80796 538280
rect 80388 538240 80796 538268
rect 80388 538228 80394 538240
rect 80790 538228 80796 538240
rect 80848 538268 80854 538280
rect 582558 538268 582564 538280
rect 80848 538240 582564 538268
rect 80848 538228 80854 538240
rect 582558 538228 582564 538240
rect 582616 538228 582622 538280
rect 32398 538160 32404 538212
rect 32456 538200 32462 538212
rect 70670 538200 70676 538212
rect 32456 538172 70676 538200
rect 32456 538160 32462 538172
rect 70670 538160 70676 538172
rect 70728 538160 70734 538212
rect 86862 538160 86868 538212
rect 86920 538200 86926 538212
rect 133138 538200 133144 538212
rect 86920 538172 133144 538200
rect 86920 538160 86926 538172
rect 133138 538160 133144 538172
rect 133196 538160 133202 538212
rect 72418 537480 72424 537532
rect 72476 537520 72482 537532
rect 579798 537520 579804 537532
rect 72476 537492 579804 537520
rect 72476 537480 72482 537492
rect 579798 537480 579804 537492
rect 579856 537480 579862 537532
rect 76006 536732 76012 536784
rect 76064 536772 76070 536784
rect 124858 536772 124864 536784
rect 76064 536744 124864 536772
rect 76064 536732 76070 536744
rect 124858 536732 124864 536744
rect 124916 536732 124922 536784
rect 85482 536188 85488 536240
rect 85540 536228 85546 536240
rect 86218 536228 86224 536240
rect 85540 536200 86224 536228
rect 85540 536188 85546 536200
rect 86218 536188 86224 536200
rect 86276 536188 86282 536240
rect 66162 536120 66168 536172
rect 66220 536160 66226 536172
rect 76006 536160 76012 536172
rect 66220 536132 76012 536160
rect 66220 536120 66226 536132
rect 76006 536120 76012 536132
rect 76064 536120 76070 536172
rect 4798 536052 4804 536104
rect 4856 536092 4862 536104
rect 45462 536092 45468 536104
rect 4856 536064 45468 536092
rect 4856 536052 4862 536064
rect 45462 536052 45468 536064
rect 45520 536092 45526 536104
rect 73154 536092 73160 536104
rect 45520 536064 73160 536092
rect 45520 536052 45526 536064
rect 73154 536052 73160 536064
rect 73212 536052 73218 536104
rect 73154 535440 73160 535492
rect 73212 535480 73218 535492
rect 73982 535480 73988 535492
rect 73212 535452 73988 535480
rect 73212 535440 73218 535452
rect 73982 535440 73988 535452
rect 74040 535440 74046 535492
rect 7558 534692 7564 534744
rect 7616 534732 7622 534744
rect 91370 534732 91376 534744
rect 7616 534704 91376 534732
rect 7616 534692 7622 534704
rect 91370 534692 91376 534704
rect 91428 534692 91434 534744
rect 56410 534012 56416 534064
rect 56468 534052 56474 534064
rect 580258 534052 580264 534064
rect 56468 534024 580264 534052
rect 56468 534012 56474 534024
rect 580258 534012 580264 534024
rect 580316 534012 580322 534064
rect 78674 533400 78680 533452
rect 78732 533440 78738 533452
rect 79502 533440 79508 533452
rect 78732 533412 79508 533440
rect 78732 533400 78738 533412
rect 79502 533400 79508 533412
rect 79560 533400 79566 533452
rect 5442 533332 5448 533384
rect 5500 533372 5506 533384
rect 91186 533372 91192 533384
rect 5500 533344 91192 533372
rect 5500 533332 5506 533344
rect 91186 533332 91192 533344
rect 91244 533332 91250 533384
rect 66070 531972 66076 532024
rect 66128 532012 66134 532024
rect 77938 532012 77944 532024
rect 66128 531984 77944 532012
rect 66128 531972 66134 531984
rect 77938 531972 77944 531984
rect 77996 531972 78002 532024
rect 15838 530544 15844 530596
rect 15896 530584 15902 530596
rect 91094 530584 91100 530596
rect 15896 530556 91100 530584
rect 15896 530544 15902 530556
rect 91094 530544 91100 530556
rect 91152 530544 91158 530596
rect 3510 514768 3516 514820
rect 3568 514808 3574 514820
rect 14458 514808 14464 514820
rect 3568 514780 14464 514808
rect 3568 514768 3574 514780
rect 14458 514768 14464 514780
rect 14516 514768 14522 514820
rect 102778 512592 102784 512644
rect 102836 512632 102842 512644
rect 122926 512632 122932 512644
rect 102836 512604 122932 512632
rect 102836 512592 102842 512604
rect 122926 512592 122932 512604
rect 122984 512592 122990 512644
rect 44082 511232 44088 511284
rect 44140 511272 44146 511284
rect 580166 511272 580172 511284
rect 44140 511244 580172 511272
rect 44140 511232 44146 511244
rect 580166 511232 580172 511244
rect 580224 511232 580230 511284
rect 3326 502052 3332 502104
rect 3384 502092 3390 502104
rect 7558 502092 7564 502104
rect 3384 502064 7564 502092
rect 3384 502052 3390 502064
rect 7558 502052 7564 502064
rect 7616 502052 7622 502104
rect 4062 475328 4068 475380
rect 4120 475368 4126 475380
rect 5442 475368 5448 475380
rect 4120 475340 5448 475368
rect 4120 475328 4126 475340
rect 5442 475328 5448 475340
rect 5500 475368 5506 475380
rect 11698 475368 11704 475380
rect 5500 475340 11704 475368
rect 5500 475328 5506 475340
rect 11698 475328 11704 475340
rect 11756 475328 11762 475380
rect 54846 468460 54852 468512
rect 54904 468500 54910 468512
rect 77294 468500 77300 468512
rect 54904 468472 77300 468500
rect 54904 468460 54910 468472
rect 77294 468460 77300 468472
rect 77352 468460 77358 468512
rect 52270 465672 52276 465724
rect 52328 465712 52334 465724
rect 95878 465712 95884 465724
rect 52328 465684 95884 465712
rect 52328 465672 52334 465684
rect 95878 465672 95884 465684
rect 95936 465672 95942 465724
rect 59078 464312 59084 464364
rect 59136 464352 59142 464364
rect 80054 464352 80060 464364
rect 59136 464324 80060 464352
rect 59136 464312 59142 464324
rect 80054 464312 80060 464324
rect 80112 464312 80118 464364
rect 50798 462952 50804 463004
rect 50856 462992 50862 463004
rect 75914 462992 75920 463004
rect 50856 462964 75920 462992
rect 50856 462952 50862 462964
rect 75914 462952 75920 462964
rect 75972 462952 75978 463004
rect 94498 462952 94504 463004
rect 94556 462992 94562 463004
rect 125686 462992 125692 463004
rect 94556 462964 125692 462992
rect 94556 462952 94562 462964
rect 125686 462952 125692 462964
rect 125744 462952 125750 463004
rect 2774 462544 2780 462596
rect 2832 462584 2838 462596
rect 4798 462584 4804 462596
rect 2832 462556 4804 462584
rect 2832 462544 2838 462556
rect 4798 462544 4804 462556
rect 4856 462544 4862 462596
rect 52270 461592 52276 461644
rect 52328 461632 52334 461644
rect 78674 461632 78680 461644
rect 52328 461604 78680 461632
rect 52328 461592 52334 461604
rect 78674 461592 78680 461604
rect 78732 461592 78738 461644
rect 63310 460912 63316 460964
rect 63368 460952 63374 460964
rect 86954 460952 86960 460964
rect 63368 460924 86960 460952
rect 63368 460912 63374 460924
rect 86954 460912 86960 460924
rect 87012 460912 87018 460964
rect 64690 460164 64696 460216
rect 64748 460204 64754 460216
rect 78674 460204 78680 460216
rect 64748 460176 78680 460204
rect 64748 460164 64754 460176
rect 78674 460164 78680 460176
rect 78732 460164 78738 460216
rect 64690 458872 64696 458924
rect 64748 458912 64754 458924
rect 70486 458912 70492 458924
rect 64748 458884 70492 458912
rect 64748 458872 64754 458884
rect 70486 458872 70492 458884
rect 70544 458872 70550 458924
rect 59170 458804 59176 458856
rect 59228 458844 59234 458856
rect 85574 458844 85580 458856
rect 59228 458816 85580 458844
rect 59228 458804 59234 458816
rect 85574 458804 85580 458816
rect 85632 458804 85638 458856
rect 77294 458192 77300 458244
rect 77352 458232 77358 458244
rect 77938 458232 77944 458244
rect 77352 458204 77944 458232
rect 77352 458192 77358 458204
rect 77938 458192 77944 458204
rect 77996 458232 78002 458244
rect 124858 458232 124864 458244
rect 77996 458204 124864 458232
rect 77996 458192 78002 458204
rect 124858 458192 124864 458204
rect 124916 458192 124922 458244
rect 61746 457512 61752 457564
rect 61804 457552 61810 457564
rect 73154 457552 73160 457564
rect 61804 457524 73160 457552
rect 61804 457512 61810 457524
rect 73154 457512 73160 457524
rect 73212 457512 73218 457564
rect 50890 457444 50896 457496
rect 50948 457484 50954 457496
rect 83458 457484 83464 457496
rect 50948 457456 83464 457484
rect 50948 457444 50954 457456
rect 83458 457444 83464 457456
rect 83516 457444 83522 457496
rect 105630 457444 105636 457496
rect 105688 457484 105694 457496
rect 123018 457484 123024 457496
rect 105688 457456 123024 457484
rect 105688 457444 105694 457456
rect 123018 457444 123024 457456
rect 123076 457444 123082 457496
rect 98546 456764 98552 456816
rect 98604 456804 98610 456816
rect 98730 456804 98736 456816
rect 98604 456776 98736 456804
rect 98604 456764 98610 456776
rect 98730 456764 98736 456776
rect 98788 456804 98794 456816
rect 151078 456804 151084 456816
rect 98788 456776 151084 456804
rect 98788 456764 98794 456776
rect 151078 456764 151084 456776
rect 151136 456764 151142 456816
rect 61930 456016 61936 456068
rect 61988 456056 61994 456068
rect 91094 456056 91100 456068
rect 61988 456028 91100 456056
rect 61988 456016 61994 456028
rect 91094 456016 91100 456028
rect 91152 456016 91158 456068
rect 101490 456016 101496 456068
rect 101548 456056 101554 456068
rect 123202 456056 123208 456068
rect 101548 456028 123208 456056
rect 101548 456016 101554 456028
rect 123202 456016 123208 456028
rect 123260 456016 123266 456068
rect 112438 455404 112444 455456
rect 112496 455444 112502 455456
rect 152458 455444 152464 455456
rect 112496 455416 152464 455444
rect 112496 455404 112502 455416
rect 152458 455404 152464 455416
rect 152516 455404 152522 455456
rect 55030 454724 55036 454776
rect 55088 454764 55094 454776
rect 72050 454764 72056 454776
rect 55088 454736 72056 454764
rect 55088 454724 55094 454736
rect 72050 454724 72056 454736
rect 72108 454724 72114 454776
rect 35802 454656 35808 454708
rect 35860 454696 35866 454708
rect 71038 454696 71044 454708
rect 35860 454668 71044 454696
rect 35860 454656 35866 454668
rect 71038 454656 71044 454668
rect 71096 454656 71102 454708
rect 91094 454044 91100 454096
rect 91152 454084 91158 454096
rect 158714 454084 158720 454096
rect 91152 454056 158720 454084
rect 91152 454044 91158 454056
rect 158714 454044 158720 454056
rect 158772 454044 158778 454096
rect 67726 453976 67732 454028
rect 67784 454016 67790 454028
rect 68278 454016 68284 454028
rect 67784 453988 68284 454016
rect 67784 453976 67790 453988
rect 68278 453976 68284 453988
rect 68336 453976 68342 454028
rect 49602 453296 49608 453348
rect 49660 453336 49666 453348
rect 68738 453336 68744 453348
rect 49660 453308 68744 453336
rect 49660 453296 49666 453308
rect 68738 453296 68744 453308
rect 68796 453296 68802 453348
rect 91738 453296 91744 453348
rect 91796 453336 91802 453348
rect 121638 453336 121644 453348
rect 91796 453308 121644 453336
rect 91796 453296 91802 453308
rect 121638 453296 121644 453308
rect 121696 453296 121702 453348
rect 68278 452684 68284 452736
rect 68336 452724 68342 452736
rect 82078 452724 82084 452736
rect 68336 452696 82084 452724
rect 68336 452684 68342 452696
rect 82078 452684 82084 452696
rect 82136 452684 82142 452736
rect 72050 452616 72056 452668
rect 72108 452656 72114 452668
rect 127618 452656 127624 452668
rect 72108 452628 127624 452656
rect 72108 452616 72114 452628
rect 127618 452616 127624 452628
rect 127676 452616 127682 452668
rect 61838 451936 61844 451988
rect 61896 451976 61902 451988
rect 72418 451976 72424 451988
rect 61896 451948 72424 451976
rect 61896 451936 61902 451948
rect 72418 451936 72424 451948
rect 72476 451936 72482 451988
rect 3418 451868 3424 451920
rect 3476 451908 3482 451920
rect 120810 451908 120816 451920
rect 3476 451880 120816 451908
rect 3476 451868 3482 451880
rect 120810 451868 120816 451880
rect 120868 451868 120874 451920
rect 14458 451188 14464 451240
rect 14516 451228 14522 451240
rect 112438 451228 112444 451240
rect 14516 451200 112444 451228
rect 14516 451188 14522 451200
rect 112438 451188 112444 451200
rect 112496 451188 112502 451240
rect 116578 449964 116584 450016
rect 116636 450004 116642 450016
rect 161566 450004 161572 450016
rect 116636 449976 161572 450004
rect 116636 449964 116642 449976
rect 161566 449964 161572 449976
rect 161624 449964 161630 450016
rect 71038 449896 71044 449948
rect 71096 449936 71102 449948
rect 73246 449936 73252 449948
rect 71096 449908 73252 449936
rect 71096 449896 71102 449908
rect 73246 449896 73252 449908
rect 73304 449936 73310 449948
rect 144178 449936 144184 449948
rect 73304 449908 144184 449936
rect 73304 449896 73310 449908
rect 144178 449896 144184 449908
rect 144236 449896 144242 449948
rect 64598 449216 64604 449268
rect 64656 449256 64662 449268
rect 74626 449256 74632 449268
rect 64656 449228 74632 449256
rect 64656 449216 64662 449228
rect 74626 449216 74632 449228
rect 74684 449216 74690 449268
rect 48130 449148 48136 449200
rect 48188 449188 48194 449200
rect 80054 449188 80060 449200
rect 48188 449160 80060 449188
rect 48188 449148 48194 449160
rect 80054 449148 80060 449160
rect 80112 449148 80118 449200
rect 169018 449148 169024 449200
rect 169076 449188 169082 449200
rect 169662 449188 169668 449200
rect 169076 449160 169668 449188
rect 169076 449148 169082 449160
rect 169662 449148 169668 449160
rect 169720 449188 169726 449200
rect 582466 449188 582472 449200
rect 169720 449160 582472 449188
rect 169720 449148 169726 449160
rect 582466 449148 582472 449160
rect 582524 449148 582530 449200
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 14458 448576 14464 448588
rect 3200 448548 14464 448576
rect 3200 448536 3206 448548
rect 14458 448536 14464 448548
rect 14516 448536 14522 448588
rect 80054 448536 80060 448588
rect 80112 448576 80118 448588
rect 80882 448576 80888 448588
rect 80112 448548 80888 448576
rect 80112 448536 80118 448548
rect 80882 448536 80888 448548
rect 80940 448576 80946 448588
rect 169018 448576 169024 448588
rect 80940 448548 169024 448576
rect 80940 448536 80946 448548
rect 169018 448536 169024 448548
rect 169076 448536 169082 448588
rect 4798 447788 4804 447840
rect 4856 447828 4862 447840
rect 68462 447828 68468 447840
rect 4856 447800 68468 447828
rect 4856 447788 4862 447800
rect 68462 447788 68468 447800
rect 68520 447788 68526 447840
rect 115198 447788 115204 447840
rect 115256 447828 115262 447840
rect 124306 447828 124312 447840
rect 115256 447800 124312 447828
rect 115256 447788 115262 447800
rect 124306 447788 124312 447800
rect 124364 447788 124370 447840
rect 68462 447176 68468 447228
rect 68520 447216 68526 447228
rect 68646 447216 68652 447228
rect 68520 447188 68652 447216
rect 68520 447176 68526 447188
rect 68646 447176 68652 447188
rect 68704 447216 68710 447228
rect 103514 447216 103520 447228
rect 68704 447188 103520 447216
rect 68704 447176 68710 447188
rect 103514 447176 103520 447188
rect 103572 447176 103578 447228
rect 49602 447108 49608 447160
rect 49660 447148 49666 447160
rect 74718 447148 74724 447160
rect 49660 447120 74724 447148
rect 49660 447108 49666 447120
rect 74718 447108 74724 447120
rect 74776 447108 74782 447160
rect 95878 447108 95884 447160
rect 95936 447148 95942 447160
rect 171134 447148 171140 447160
rect 95936 447120 171140 447148
rect 95936 447108 95942 447120
rect 171134 447108 171140 447120
rect 171192 447108 171198 447160
rect 78674 446904 78680 446956
rect 78732 446944 78738 446956
rect 79134 446944 79140 446956
rect 78732 446916 79140 446944
rect 78732 446904 78738 446916
rect 79134 446904 79140 446916
rect 79192 446904 79198 446956
rect 41322 445816 41328 445868
rect 41380 445856 41386 445868
rect 79134 445856 79140 445868
rect 41380 445828 79140 445856
rect 41380 445816 41386 445828
rect 79134 445816 79140 445828
rect 79192 445816 79198 445868
rect 106918 445816 106924 445868
rect 106976 445856 106982 445868
rect 124950 445856 124956 445868
rect 106976 445828 124956 445856
rect 106976 445816 106982 445828
rect 124950 445816 124956 445828
rect 125008 445816 125014 445868
rect 76558 445748 76564 445800
rect 76616 445788 76622 445800
rect 155218 445788 155224 445800
rect 76616 445760 155224 445788
rect 76616 445748 76622 445760
rect 155218 445748 155224 445760
rect 155276 445748 155282 445800
rect 54938 444456 54944 444508
rect 54996 444496 55002 444508
rect 92474 444496 92480 444508
rect 54996 444468 92480 444496
rect 54996 444456 55002 444468
rect 92474 444456 92480 444468
rect 92532 444496 92538 444508
rect 93072 444496 93078 444508
rect 92532 444468 93078 444496
rect 92532 444456 92538 444468
rect 93072 444456 93078 444468
rect 93130 444456 93136 444508
rect 101398 444456 101404 444508
rect 101456 444496 101462 444508
rect 126238 444496 126244 444508
rect 101456 444468 126244 444496
rect 101456 444456 101462 444468
rect 126238 444456 126244 444468
rect 126296 444456 126302 444508
rect 4798 444388 4804 444440
rect 4856 444428 4862 444440
rect 118694 444428 118700 444440
rect 4856 444400 118700 444428
rect 4856 444388 4862 444400
rect 118694 444388 118700 444400
rect 118752 444388 118758 444440
rect 124122 444320 124128 444372
rect 124180 444360 124186 444372
rect 132494 444360 132500 444372
rect 124180 444332 132500 444360
rect 124180 444320 124186 444332
rect 132494 444320 132500 444332
rect 132552 444360 132558 444372
rect 133782 444360 133788 444372
rect 132552 444332 133788 444360
rect 132552 444320 132558 444332
rect 133782 444320 133788 444332
rect 133840 444320 133846 444372
rect 133782 443640 133788 443692
rect 133840 443680 133846 443692
rect 165614 443680 165620 443692
rect 133840 443652 165620 443680
rect 133840 443640 133846 443652
rect 165614 443640 165620 443652
rect 165672 443640 165678 443692
rect 67266 442892 67272 442944
rect 67324 442932 67330 442944
rect 67726 442932 67732 442944
rect 67324 442904 67732 442932
rect 67324 442892 67330 442904
rect 67726 442892 67732 442904
rect 67784 442892 67790 442944
rect 124122 441600 124128 441652
rect 124180 441640 124186 441652
rect 133138 441640 133144 441652
rect 124180 441612 133144 441640
rect 124180 441600 124186 441612
rect 133138 441600 133144 441612
rect 133196 441600 133202 441652
rect 56502 440852 56508 440904
rect 56560 440892 56566 440904
rect 68278 440892 68284 440904
rect 56560 440864 68284 440892
rect 56560 440852 56566 440864
rect 68278 440852 68284 440864
rect 68336 440852 68342 440904
rect 64782 439016 64788 439068
rect 64840 439056 64846 439068
rect 66990 439056 66996 439068
rect 64840 439028 66996 439056
rect 64840 439016 64846 439028
rect 66990 439016 66996 439028
rect 67048 439056 67054 439068
rect 67266 439056 67272 439068
rect 67048 439028 67272 439056
rect 67048 439016 67054 439028
rect 67266 439016 67272 439028
rect 67324 439016 67330 439068
rect 124122 438880 124128 438932
rect 124180 438920 124186 438932
rect 186958 438920 186964 438932
rect 124180 438892 186964 438920
rect 124180 438880 124186 438892
rect 186958 438880 186964 438892
rect 187016 438880 187022 438932
rect 124122 438132 124128 438184
rect 124180 438172 124186 438184
rect 124306 438172 124312 438184
rect 124180 438144 124312 438172
rect 124180 438132 124186 438144
rect 124306 438132 124312 438144
rect 124364 438172 124370 438184
rect 157978 438172 157984 438184
rect 124364 438144 157984 438172
rect 124364 438132 124370 438144
rect 157978 438132 157984 438144
rect 158036 438132 158042 438184
rect 57698 437452 57704 437504
rect 57756 437492 57762 437504
rect 60550 437492 60556 437504
rect 57756 437464 60556 437492
rect 57756 437452 57762 437464
rect 60550 437452 60556 437464
rect 60608 437492 60614 437504
rect 66806 437492 66812 437504
rect 60608 437464 66812 437492
rect 60608 437452 60614 437464
rect 66806 437452 66812 437464
rect 66864 437452 66870 437504
rect 53650 435344 53656 435396
rect 53708 435384 53714 435396
rect 66806 435384 66812 435396
rect 53708 435356 66812 435384
rect 53708 435344 53714 435356
rect 66806 435344 66812 435356
rect 66864 435344 66870 435396
rect 124122 432556 124128 432608
rect 124180 432596 124186 432608
rect 135162 432596 135168 432608
rect 124180 432568 135168 432596
rect 124180 432556 124186 432568
rect 135162 432556 135168 432568
rect 135220 432596 135226 432608
rect 582374 432596 582380 432608
rect 135220 432568 582380 432596
rect 135220 432556 135226 432568
rect 582374 432556 582380 432568
rect 582432 432556 582438 432608
rect 60642 432012 60648 432064
rect 60700 432052 60706 432064
rect 66898 432052 66904 432064
rect 60700 432024 66904 432052
rect 60700 432012 60706 432024
rect 66898 432012 66904 432024
rect 66956 432012 66962 432064
rect 50982 431876 50988 431928
rect 51040 431916 51046 431928
rect 66898 431916 66904 431928
rect 51040 431888 66904 431916
rect 51040 431876 51046 431888
rect 66898 431876 66904 431888
rect 66956 431876 66962 431928
rect 48130 430584 48136 430636
rect 48188 430624 48194 430636
rect 50982 430624 50988 430636
rect 48188 430596 50988 430624
rect 48188 430584 48194 430596
rect 50982 430584 50988 430596
rect 51040 430584 51046 430636
rect 36722 429088 36728 429140
rect 36780 429128 36786 429140
rect 37182 429128 37188 429140
rect 36780 429100 37188 429128
rect 36780 429088 36786 429100
rect 37182 429088 37188 429100
rect 37240 429128 37246 429140
rect 66806 429128 66812 429140
rect 37240 429100 66812 429128
rect 37240 429088 37246 429100
rect 66806 429088 66812 429100
rect 66864 429088 66870 429140
rect 22738 428408 22744 428460
rect 22796 428448 22802 428460
rect 36722 428448 36728 428460
rect 22796 428420 36728 428448
rect 22796 428408 22802 428420
rect 36722 428408 36728 428420
rect 36780 428408 36786 428460
rect 44082 425688 44088 425740
rect 44140 425728 44146 425740
rect 57882 425728 57888 425740
rect 44140 425700 57888 425728
rect 44140 425688 44146 425700
rect 57882 425688 57888 425700
rect 57940 425688 57946 425740
rect 57698 425076 57704 425128
rect 57756 425116 57762 425128
rect 57882 425116 57888 425128
rect 57756 425088 57888 425116
rect 57756 425076 57762 425088
rect 57882 425076 57888 425088
rect 57940 425116 57946 425128
rect 66254 425116 66260 425128
rect 57940 425088 66260 425116
rect 57940 425076 57946 425088
rect 66254 425076 66260 425088
rect 66312 425076 66318 425128
rect 56410 424328 56416 424380
rect 56468 424368 56474 424380
rect 66070 424368 66076 424380
rect 56468 424340 66076 424368
rect 56468 424328 56474 424340
rect 66070 424328 66076 424340
rect 66128 424368 66134 424380
rect 66254 424368 66260 424380
rect 66128 424340 66260 424368
rect 66128 424328 66134 424340
rect 66254 424328 66260 424340
rect 66312 424328 66318 424380
rect 3142 422900 3148 422952
rect 3200 422940 3206 422952
rect 15838 422940 15844 422952
rect 3200 422912 15844 422940
rect 3200 422900 3206 422912
rect 15838 422900 15844 422912
rect 15896 422900 15902 422952
rect 123018 422288 123024 422340
rect 123076 422328 123082 422340
rect 123478 422328 123484 422340
rect 123076 422300 123484 422328
rect 123076 422288 123082 422300
rect 123478 422288 123484 422300
rect 123536 422328 123542 422340
rect 172514 422328 172520 422340
rect 123536 422300 172520 422328
rect 123536 422288 123542 422300
rect 172514 422288 172520 422300
rect 172572 422288 172578 422340
rect 48222 421540 48228 421592
rect 48280 421580 48286 421592
rect 61378 421580 61384 421592
rect 48280 421552 61384 421580
rect 48280 421540 48286 421552
rect 61378 421540 61384 421552
rect 61436 421580 61442 421592
rect 66254 421580 66260 421592
rect 61436 421552 66260 421580
rect 61436 421540 61442 421552
rect 66254 421540 66260 421552
rect 66312 421540 66318 421592
rect 121546 418072 121552 418124
rect 121604 418112 121610 418124
rect 126974 418112 126980 418124
rect 121604 418084 126980 418112
rect 121604 418072 121610 418084
rect 126974 418072 126980 418084
rect 127032 418072 127038 418124
rect 58986 416780 58992 416832
rect 59044 416820 59050 416832
rect 63310 416820 63316 416832
rect 59044 416792 63316 416820
rect 59044 416780 59050 416792
rect 63310 416780 63316 416792
rect 63368 416820 63374 416832
rect 66898 416820 66904 416832
rect 63368 416792 66904 416820
rect 63368 416780 63374 416792
rect 66898 416780 66904 416792
rect 66956 416780 66962 416832
rect 65518 415148 65524 415200
rect 65576 415188 65582 415200
rect 66438 415188 66444 415200
rect 65576 415160 66444 415188
rect 65576 415148 65582 415160
rect 66438 415148 66444 415160
rect 66496 415148 66502 415200
rect 124122 415148 124128 415200
rect 124180 415188 124186 415200
rect 125686 415188 125692 415200
rect 124180 415160 125692 415188
rect 124180 415148 124186 415160
rect 125686 415148 125692 415160
rect 125744 415148 125750 415200
rect 57882 414672 57888 414724
rect 57940 414712 57946 414724
rect 65518 414712 65524 414724
rect 57940 414684 65524 414712
rect 57940 414672 57946 414684
rect 65518 414672 65524 414684
rect 65576 414672 65582 414724
rect 123110 413924 123116 413976
rect 123168 413964 123174 413976
rect 128354 413964 128360 413976
rect 123168 413936 128360 413964
rect 123168 413924 123174 413936
rect 128354 413924 128360 413936
rect 128412 413924 128418 413976
rect 121638 409844 121644 409896
rect 121696 409884 121702 409896
rect 129090 409884 129096 409896
rect 121696 409856 129096 409884
rect 121696 409844 121702 409856
rect 129090 409844 129096 409856
rect 129148 409844 129154 409896
rect 63402 408416 63408 408468
rect 63460 408456 63466 408468
rect 65886 408456 65892 408468
rect 63460 408428 65892 408456
rect 63460 408416 63466 408428
rect 65886 408416 65892 408428
rect 65944 408456 65950 408468
rect 66530 408456 66536 408468
rect 65944 408428 66536 408456
rect 65944 408416 65950 408428
rect 66530 408416 66536 408428
rect 66588 408416 66594 408468
rect 124122 407736 124128 407788
rect 124180 407776 124186 407788
rect 135898 407776 135904 407788
rect 124180 407748 135904 407776
rect 124180 407736 124186 407748
rect 135898 407736 135904 407748
rect 135956 407736 135962 407788
rect 122098 407056 122104 407108
rect 122156 407096 122162 407108
rect 122926 407096 122932 407108
rect 122156 407068 122932 407096
rect 122156 407056 122162 407068
rect 122926 407056 122932 407068
rect 122984 407056 122990 407108
rect 57606 406512 57612 406564
rect 57664 406552 57670 406564
rect 57790 406552 57796 406564
rect 57664 406524 57796 406552
rect 57664 406512 57670 406524
rect 57790 406512 57796 406524
rect 57848 406512 57854 406564
rect 123202 406104 123208 406156
rect 123260 406144 123266 406156
rect 125042 406144 125048 406156
rect 123260 406116 125048 406144
rect 123260 406104 123266 406116
rect 125042 406104 125048 406116
rect 125100 406104 125106 406156
rect 62022 405764 62028 405816
rect 62080 405804 62086 405816
rect 64782 405804 64788 405816
rect 62080 405776 64788 405804
rect 62080 405764 62086 405776
rect 64782 405764 64788 405776
rect 64840 405804 64846 405816
rect 66622 405804 66628 405816
rect 64840 405776 66628 405804
rect 64840 405764 64846 405776
rect 66622 405764 66628 405776
rect 66680 405764 66686 405816
rect 57974 403588 57980 403640
rect 58032 403628 58038 403640
rect 66346 403628 66352 403640
rect 58032 403600 66352 403628
rect 58032 403588 58038 403600
rect 66346 403588 66352 403600
rect 66404 403588 66410 403640
rect 163498 403588 163504 403640
rect 163556 403628 163562 403640
rect 582374 403628 582380 403640
rect 163556 403600 582380 403628
rect 163556 403588 163562 403600
rect 582374 403588 582380 403600
rect 582432 403588 582438 403640
rect 120626 402976 120632 403028
rect 120684 403016 120690 403028
rect 163498 403016 163504 403028
rect 120684 402988 163504 403016
rect 120684 402976 120690 402988
rect 163498 402976 163504 402988
rect 163556 402976 163562 403028
rect 53650 402228 53656 402280
rect 53708 402268 53714 402280
rect 57974 402268 57980 402280
rect 53708 402240 57980 402268
rect 53708 402228 53714 402240
rect 57974 402228 57980 402240
rect 58032 402228 58038 402280
rect 50890 401548 50896 401600
rect 50948 401588 50954 401600
rect 57606 401588 57612 401600
rect 50948 401560 57612 401588
rect 50948 401548 50954 401560
rect 57606 401548 57612 401560
rect 57664 401588 57670 401600
rect 66806 401588 66812 401600
rect 57664 401560 66812 401588
rect 57664 401548 57670 401560
rect 66806 401548 66812 401560
rect 66864 401548 66870 401600
rect 124122 401480 124128 401532
rect 124180 401520 124186 401532
rect 129734 401520 129740 401532
rect 124180 401492 129740 401520
rect 124180 401480 124186 401492
rect 129734 401480 129740 401492
rect 129792 401480 129798 401532
rect 129734 400188 129740 400240
rect 129792 400228 129798 400240
rect 130378 400228 130384 400240
rect 129792 400200 130384 400228
rect 129792 400188 129798 400200
rect 130378 400188 130384 400200
rect 130436 400188 130442 400240
rect 59998 399440 60004 399492
rect 60056 399480 60062 399492
rect 66346 399480 66352 399492
rect 60056 399452 66352 399480
rect 60056 399440 60062 399452
rect 66346 399440 66352 399452
rect 66404 399440 66410 399492
rect 123478 398828 123484 398880
rect 123536 398868 123542 398880
rect 124950 398868 124956 398880
rect 123536 398840 124956 398868
rect 123536 398828 123542 398840
rect 124950 398828 124956 398840
rect 125008 398828 125014 398880
rect 2774 398692 2780 398744
rect 2832 398732 2838 398744
rect 4798 398732 4804 398744
rect 2832 398704 4804 398732
rect 2832 398692 2838 398704
rect 4798 398692 4804 398704
rect 4856 398692 4862 398744
rect 43990 398080 43996 398132
rect 44048 398120 44054 398132
rect 52362 398120 52368 398132
rect 44048 398092 52368 398120
rect 44048 398080 44054 398092
rect 52362 398080 52368 398092
rect 52420 398120 52426 398132
rect 59998 398120 60004 398132
rect 52420 398092 60004 398120
rect 52420 398080 52426 398092
rect 59998 398080 60004 398092
rect 60056 398080 60062 398132
rect 39942 396720 39948 396772
rect 40000 396760 40006 396772
rect 66990 396760 66996 396772
rect 40000 396732 66996 396760
rect 40000 396720 40006 396732
rect 66990 396720 66996 396732
rect 67048 396720 67054 396772
rect 121454 396040 121460 396092
rect 121512 396080 121518 396092
rect 180058 396080 180064 396092
rect 121512 396052 180064 396080
rect 121512 396040 121518 396052
rect 180058 396040 180064 396052
rect 180116 396040 180122 396092
rect 123662 395496 123668 395548
rect 123720 395536 123726 395548
rect 125594 395536 125600 395548
rect 123720 395508 125600 395536
rect 123720 395496 123726 395508
rect 125594 395496 125600 395508
rect 125652 395496 125658 395548
rect 55122 393252 55128 393304
rect 55180 393292 55186 393304
rect 66254 393292 66260 393304
rect 55180 393264 66260 393292
rect 55180 393252 55186 393264
rect 66254 393252 66260 393264
rect 66312 393252 66318 393304
rect 124950 391960 124956 392012
rect 125008 392000 125014 392012
rect 172606 392000 172612 392012
rect 125008 391972 172612 392000
rect 125008 391960 125014 391972
rect 172606 391960 172612 391972
rect 172664 391960 172670 392012
rect 15838 391348 15844 391400
rect 15896 391388 15902 391400
rect 124950 391388 124956 391400
rect 15896 391360 124956 391388
rect 15896 391348 15902 391360
rect 124950 391348 124956 391360
rect 125008 391348 125014 391400
rect 111702 389784 111708 389836
rect 111760 389824 111766 389836
rect 121546 389824 121552 389836
rect 111760 389796 121552 389824
rect 111760 389784 111766 389796
rect 121546 389784 121552 389796
rect 121604 389784 121610 389836
rect 61746 389240 61752 389292
rect 61804 389280 61810 389292
rect 77386 389280 77392 389292
rect 61804 389252 77392 389280
rect 61804 389240 61810 389252
rect 77386 389240 77392 389252
rect 77444 389240 77450 389292
rect 11698 389172 11704 389224
rect 11756 389212 11762 389224
rect 111610 389212 111616 389224
rect 11756 389184 111616 389212
rect 11756 389172 11762 389184
rect 111610 389172 111616 389184
rect 111668 389172 111674 389224
rect 169754 389212 169760 389224
rect 135180 389184 169760 389212
rect 102594 389104 102600 389156
rect 102652 389144 102658 389156
rect 105538 389144 105544 389156
rect 102652 389116 105544 389144
rect 102652 389104 102658 389116
rect 105538 389104 105544 389116
rect 105596 389104 105602 389156
rect 117866 389104 117872 389156
rect 117924 389144 117930 389156
rect 134518 389144 134524 389156
rect 117924 389116 134524 389144
rect 117924 389104 117930 389116
rect 134518 389104 134524 389116
rect 134576 389144 134582 389156
rect 135180 389144 135208 389184
rect 169754 389172 169760 389184
rect 169812 389172 169818 389224
rect 134576 389116 135208 389144
rect 134576 389104 134582 389116
rect 64690 388424 64696 388476
rect 64748 388464 64754 388476
rect 71774 388464 71780 388476
rect 64748 388436 71780 388464
rect 64748 388424 64754 388436
rect 71774 388424 71780 388436
rect 71832 388424 71838 388476
rect 93394 388424 93400 388476
rect 93452 388464 93458 388476
rect 100018 388464 100024 388476
rect 93452 388436 100024 388464
rect 93452 388424 93458 388436
rect 100018 388424 100024 388436
rect 100076 388424 100082 388476
rect 101398 388424 101404 388476
rect 101456 388464 101462 388476
rect 120166 388464 120172 388476
rect 101456 388436 120172 388464
rect 101456 388424 101462 388436
rect 120166 388424 120172 388436
rect 120224 388424 120230 388476
rect 93762 388356 93768 388408
rect 93820 388396 93826 388408
rect 94222 388396 94228 388408
rect 93820 388368 94228 388396
rect 93820 388356 93826 388368
rect 94222 388356 94228 388368
rect 94280 388356 94286 388408
rect 71774 387812 71780 387864
rect 71832 387852 71838 387864
rect 73154 387852 73160 387864
rect 71832 387824 73160 387852
rect 71832 387812 71838 387824
rect 73154 387812 73160 387824
rect 73212 387812 73218 387864
rect 111610 387812 111616 387864
rect 111668 387852 111674 387864
rect 112438 387852 112444 387864
rect 111668 387824 112444 387852
rect 111668 387812 111674 387824
rect 112438 387812 112444 387824
rect 112496 387812 112502 387864
rect 45462 387744 45468 387796
rect 45520 387784 45526 387796
rect 76558 387784 76564 387796
rect 45520 387756 76564 387784
rect 45520 387744 45526 387756
rect 76558 387744 76564 387756
rect 76616 387744 76622 387796
rect 3418 387064 3424 387116
rect 3476 387104 3482 387116
rect 89714 387104 89720 387116
rect 3476 387076 89720 387104
rect 3476 387064 3482 387076
rect 89714 387064 89720 387076
rect 89772 387064 89778 387116
rect 104066 387064 104072 387116
rect 104124 387104 104130 387116
rect 135070 387104 135076 387116
rect 104124 387076 135076 387104
rect 104124 387064 104130 387076
rect 135070 387064 135076 387076
rect 135128 387104 135134 387116
rect 136634 387104 136640 387116
rect 135128 387076 136640 387104
rect 135128 387064 135134 387076
rect 136634 387064 136640 387076
rect 136692 387064 136698 387116
rect 61838 386316 61844 386368
rect 61896 386356 61902 386368
rect 74626 386356 74632 386368
rect 61896 386328 74632 386356
rect 61896 386316 61902 386328
rect 74626 386316 74632 386328
rect 74684 386316 74690 386368
rect 77202 385636 77208 385688
rect 77260 385676 77266 385688
rect 113174 385676 113180 385688
rect 77260 385648 113180 385676
rect 77260 385636 77266 385648
rect 113174 385636 113180 385648
rect 113232 385636 113238 385688
rect 65978 384956 65984 385008
rect 66036 384996 66042 385008
rect 85574 384996 85580 385008
rect 66036 384968 85580 384996
rect 66036 384956 66042 384968
rect 85574 384956 85580 384968
rect 85632 384996 85638 385008
rect 86218 384996 86224 385008
rect 85632 384968 86224 384996
rect 85632 384956 85638 384968
rect 86218 384956 86224 384968
rect 86276 384956 86282 385008
rect 15838 384276 15844 384328
rect 15896 384316 15902 384328
rect 123110 384316 123116 384328
rect 15896 384288 123116 384316
rect 15896 384276 15902 384288
rect 123110 384276 123116 384288
rect 123168 384276 123174 384328
rect 110230 382916 110236 382968
rect 110288 382956 110294 382968
rect 177482 382956 177488 382968
rect 110288 382928 177488 382956
rect 110288 382916 110294 382928
rect 177482 382916 177488 382928
rect 177540 382916 177546 382968
rect 7558 382236 7564 382288
rect 7616 382276 7622 382288
rect 118694 382276 118700 382288
rect 7616 382248 118700 382276
rect 7616 382236 7622 382248
rect 118694 382236 118700 382248
rect 118752 382276 118758 382288
rect 119430 382276 119436 382288
rect 118752 382248 119436 382276
rect 118752 382236 118758 382248
rect 119430 382236 119436 382248
rect 119488 382236 119494 382288
rect 4798 381488 4804 381540
rect 4856 381528 4862 381540
rect 105630 381528 105636 381540
rect 4856 381500 105636 381528
rect 4856 381488 4862 381500
rect 105630 381488 105636 381500
rect 105688 381528 105694 381540
rect 175274 381528 175280 381540
rect 105688 381500 175280 381528
rect 105688 381488 105694 381500
rect 175274 381488 175280 381500
rect 175332 381488 175338 381540
rect 50798 380808 50804 380860
rect 50856 380848 50862 380860
rect 81434 380848 81440 380860
rect 50856 380820 81440 380848
rect 50856 380808 50862 380820
rect 81434 380808 81440 380820
rect 81492 380808 81498 380860
rect 81434 379584 81440 379636
rect 81492 379624 81498 379636
rect 82078 379624 82084 379636
rect 81492 379596 82084 379624
rect 81492 379584 81498 379596
rect 82078 379584 82084 379596
rect 82136 379584 82142 379636
rect 72418 379516 72424 379568
rect 72476 379556 72482 379568
rect 73062 379556 73068 379568
rect 72476 379528 73068 379556
rect 72476 379516 72482 379528
rect 73062 379516 73068 379528
rect 73120 379556 73126 379568
rect 188338 379556 188344 379568
rect 73120 379528 188344 379556
rect 73120 379516 73126 379528
rect 188338 379516 188344 379528
rect 188396 379516 188402 379568
rect 64782 378836 64788 378888
rect 64840 378876 64846 378888
rect 108298 378876 108304 378888
rect 64840 378848 108304 378876
rect 64840 378836 64846 378848
rect 108298 378836 108304 378848
rect 108356 378836 108362 378888
rect 99282 378768 99288 378820
rect 99340 378808 99346 378820
rect 165706 378808 165712 378820
rect 99340 378780 165712 378808
rect 99340 378768 99346 378780
rect 165706 378768 165712 378780
rect 165764 378768 165770 378820
rect 52270 378088 52276 378140
rect 52328 378128 52334 378140
rect 86954 378128 86960 378140
rect 52328 378100 86960 378128
rect 52328 378088 52334 378100
rect 86954 378088 86960 378100
rect 87012 378088 87018 378140
rect 53558 376728 53564 376780
rect 53616 376768 53622 376780
rect 53742 376768 53748 376780
rect 53616 376740 53748 376768
rect 53616 376728 53622 376740
rect 53742 376728 53748 376740
rect 53800 376768 53806 376780
rect 185578 376768 185584 376780
rect 53800 376740 185584 376768
rect 53800 376728 53806 376740
rect 185578 376728 185584 376740
rect 185636 376728 185642 376780
rect 67726 374620 67732 374672
rect 67784 374660 67790 374672
rect 124950 374660 124956 374672
rect 67784 374632 124956 374660
rect 67784 374620 67790 374632
rect 124950 374620 124956 374632
rect 125008 374620 125014 374672
rect 86218 374008 86224 374060
rect 86276 374048 86282 374060
rect 211798 374048 211804 374060
rect 86276 374020 211804 374048
rect 86276 374008 86282 374020
rect 211798 374008 211804 374020
rect 211856 374008 211862 374060
rect 60642 373260 60648 373312
rect 60700 373300 60706 373312
rect 164878 373300 164884 373312
rect 60700 373272 164884 373300
rect 60700 373260 60706 373272
rect 164878 373260 164884 373272
rect 164936 373260 164942 373312
rect 122098 372580 122104 372632
rect 122156 372620 122162 372632
rect 122742 372620 122748 372632
rect 122156 372592 122748 372620
rect 122156 372580 122162 372592
rect 122742 372580 122748 372592
rect 122800 372620 122806 372632
rect 204898 372620 204904 372632
rect 122800 372592 204904 372620
rect 122800 372580 122806 372592
rect 204898 372580 204904 372592
rect 204956 372580 204962 372632
rect 70302 371832 70308 371884
rect 70360 371872 70366 371884
rect 166994 371872 167000 371884
rect 70360 371844 167000 371872
rect 70360 371832 70366 371844
rect 166994 371832 167000 371844
rect 167052 371832 167058 371884
rect 125042 371220 125048 371272
rect 125100 371260 125106 371272
rect 125502 371260 125508 371272
rect 125100 371232 125508 371260
rect 125100 371220 125106 371232
rect 125502 371220 125508 371232
rect 125560 371260 125566 371272
rect 258074 371260 258080 371272
rect 125560 371232 258080 371260
rect 125560 371220 125566 371232
rect 258074 371220 258080 371232
rect 258132 371220 258138 371272
rect 139302 369928 139308 369980
rect 139360 369968 139366 369980
rect 242158 369968 242164 369980
rect 139360 369940 242164 369968
rect 139360 369928 139366 369940
rect 242158 369928 242164 369940
rect 242216 369928 242222 369980
rect 125594 369860 125600 369912
rect 125652 369900 125658 369912
rect 126238 369900 126244 369912
rect 125652 369872 126244 369900
rect 125652 369860 125658 369872
rect 126238 369860 126244 369872
rect 126296 369900 126302 369912
rect 231118 369900 231124 369912
rect 126296 369872 231124 369900
rect 126296 369860 126302 369872
rect 231118 369860 231124 369872
rect 231176 369860 231182 369912
rect 142798 369112 142804 369164
rect 142856 369152 142862 369164
rect 174630 369152 174636 369164
rect 142856 369124 174636 369152
rect 142856 369112 142862 369124
rect 174630 369112 174636 369124
rect 174688 369112 174694 369164
rect 121362 368500 121368 368552
rect 121420 368540 121426 368552
rect 182818 368540 182824 368552
rect 121420 368512 182824 368540
rect 121420 368500 121426 368512
rect 182818 368500 182824 368512
rect 182876 368500 182882 368552
rect 119430 367752 119436 367804
rect 119488 367792 119494 367804
rect 171226 367792 171232 367804
rect 119488 367764 171232 367792
rect 119488 367752 119494 367764
rect 171226 367752 171232 367764
rect 171284 367752 171290 367804
rect 137922 367072 137928 367124
rect 137980 367112 137986 367124
rect 327074 367112 327080 367124
rect 137980 367084 327080 367112
rect 137980 367072 137986 367084
rect 327074 367072 327080 367084
rect 327132 367072 327138 367124
rect 81342 366324 81348 366376
rect 81400 366364 81406 366376
rect 96430 366364 96436 366376
rect 81400 366336 96436 366364
rect 81400 366324 81406 366336
rect 96430 366324 96436 366336
rect 96488 366324 96494 366376
rect 124858 365780 124864 365832
rect 124916 365820 124922 365832
rect 214558 365820 214564 365832
rect 124916 365792 214564 365820
rect 124916 365780 124922 365792
rect 214558 365780 214564 365792
rect 214616 365780 214622 365832
rect 104894 365712 104900 365764
rect 104952 365752 104958 365764
rect 224218 365752 224224 365764
rect 104952 365724 224224 365752
rect 104952 365712 104958 365724
rect 224218 365712 224224 365724
rect 224276 365712 224282 365764
rect 81434 365644 81440 365696
rect 81492 365684 81498 365696
rect 82078 365684 82084 365696
rect 81492 365656 82084 365684
rect 81492 365644 81498 365656
rect 82078 365644 82084 365656
rect 82136 365644 82142 365696
rect 143442 364420 143448 364472
rect 143500 364460 143506 364472
rect 238018 364460 238024 364472
rect 143500 364432 238024 364460
rect 143500 364420 143506 364432
rect 238018 364420 238024 364432
rect 238076 364420 238082 364472
rect 81434 364352 81440 364404
rect 81492 364392 81498 364404
rect 238110 364392 238116 364404
rect 81492 364364 238116 364392
rect 81492 364352 81498 364364
rect 238110 364352 238116 364364
rect 238168 364352 238174 364404
rect 131114 362992 131120 363044
rect 131172 363032 131178 363044
rect 214650 363032 214656 363044
rect 131172 363004 214656 363032
rect 131172 362992 131178 363004
rect 214650 362992 214656 363004
rect 214708 362992 214714 363044
rect 90358 362924 90364 362976
rect 90416 362964 90422 362976
rect 188430 362964 188436 362976
rect 90416 362936 188436 362964
rect 90416 362924 90422 362936
rect 188430 362924 188436 362936
rect 188488 362924 188494 362976
rect 137278 362652 137284 362704
rect 137336 362692 137342 362704
rect 137830 362692 137836 362704
rect 137336 362664 137836 362692
rect 137336 362652 137342 362664
rect 137830 362652 137836 362664
rect 137888 362652 137894 362704
rect 63218 362176 63224 362228
rect 63276 362216 63282 362228
rect 87046 362216 87052 362228
rect 63276 362188 87052 362216
rect 63276 362176 63282 362188
rect 87046 362176 87052 362188
rect 87104 362216 87110 362228
rect 87966 362216 87972 362228
rect 87104 362188 87972 362216
rect 87104 362176 87110 362188
rect 87966 362176 87972 362188
rect 88024 362176 88030 362228
rect 137830 361632 137836 361684
rect 137888 361672 137894 361684
rect 164234 361672 164240 361684
rect 137888 361644 164240 361672
rect 137888 361632 137894 361644
rect 164234 361632 164240 361644
rect 164292 361632 164298 361684
rect 87966 361564 87972 361616
rect 88024 361604 88030 361616
rect 240226 361604 240232 361616
rect 88024 361576 240232 361604
rect 88024 361564 88030 361576
rect 240226 361564 240232 361576
rect 240284 361564 240290 361616
rect 50798 361496 50804 361548
rect 50856 361536 50862 361548
rect 54846 361536 54852 361548
rect 50856 361508 54852 361536
rect 50856 361496 50862 361508
rect 54846 361496 54852 361508
rect 54904 361536 54910 361548
rect 82814 361536 82820 361548
rect 54904 361508 82820 361536
rect 54904 361496 54910 361508
rect 82814 361496 82820 361508
rect 82872 361496 82878 361548
rect 92290 360816 92296 360868
rect 92348 360856 92354 360868
rect 118694 360856 118700 360868
rect 92348 360828 118700 360856
rect 92348 360816 92354 360828
rect 118694 360816 118700 360828
rect 118752 360816 118758 360868
rect 124950 360272 124956 360324
rect 125008 360312 125014 360324
rect 178678 360312 178684 360324
rect 125008 360284 178684 360312
rect 125008 360272 125014 360284
rect 178678 360272 178684 360284
rect 178736 360272 178742 360324
rect 99282 360204 99288 360256
rect 99340 360244 99346 360256
rect 226978 360244 226984 360256
rect 99340 360216 226984 360244
rect 99340 360204 99346 360216
rect 226978 360204 226984 360216
rect 227036 360204 227042 360256
rect 66070 359456 66076 359508
rect 66128 359496 66134 359508
rect 127710 359496 127716 359508
rect 66128 359468 127716 359496
rect 66128 359456 66134 359468
rect 127710 359456 127716 359468
rect 127768 359456 127774 359508
rect 128354 358844 128360 358896
rect 128412 358884 128418 358896
rect 181530 358884 181536 358896
rect 128412 358856 181536 358884
rect 128412 358844 128418 358856
rect 181530 358844 181536 358856
rect 181588 358844 181594 358896
rect 136634 358776 136640 358828
rect 136692 358816 136698 358828
rect 238754 358816 238760 358828
rect 136692 358788 238760 358816
rect 136692 358776 136698 358788
rect 238754 358776 238760 358788
rect 238812 358776 238818 358828
rect 3510 358572 3516 358624
rect 3568 358612 3574 358624
rect 7558 358612 7564 358624
rect 3568 358584 7564 358612
rect 3568 358572 3574 358584
rect 7558 358572 7564 358584
rect 7616 358572 7622 358624
rect 93762 358028 93768 358080
rect 93820 358068 93826 358080
rect 131114 358068 131120 358080
rect 93820 358040 131120 358068
rect 93820 358028 93826 358040
rect 131114 358028 131120 358040
rect 131172 358028 131178 358080
rect 118694 357416 118700 357468
rect 118752 357456 118758 357468
rect 225598 357456 225604 357468
rect 118752 357428 225604 357456
rect 118752 357416 118758 357428
rect 225598 357416 225604 357428
rect 225656 357416 225662 357468
rect 64782 356668 64788 356720
rect 64840 356708 64846 356720
rect 111794 356708 111800 356720
rect 64840 356680 111800 356708
rect 64840 356668 64846 356680
rect 111794 356668 111800 356680
rect 111852 356668 111858 356720
rect 70394 356600 70400 356652
rect 70452 356640 70458 356652
rect 71682 356640 71688 356652
rect 70452 356612 71688 356640
rect 70452 356600 70458 356612
rect 71682 356600 71688 356612
rect 71740 356600 71746 356652
rect 141418 356124 141424 356176
rect 141476 356164 141482 356176
rect 231210 356164 231216 356176
rect 141476 356136 231216 356164
rect 141476 356124 141482 356136
rect 231210 356124 231216 356136
rect 231268 356124 231274 356176
rect 71682 356056 71688 356108
rect 71740 356096 71746 356108
rect 255406 356096 255412 356108
rect 71740 356068 255412 356096
rect 71740 356056 71746 356068
rect 255406 356056 255412 356068
rect 255464 356056 255470 356108
rect 155218 355988 155224 356040
rect 155276 356028 155282 356040
rect 155954 356028 155960 356040
rect 155276 356000 155960 356028
rect 155276 355988 155282 356000
rect 155954 355988 155960 356000
rect 156012 355988 156018 356040
rect 97810 355308 97816 355360
rect 97868 355348 97874 355360
rect 155310 355348 155316 355360
rect 97868 355320 155316 355348
rect 97868 355308 97874 355320
rect 155310 355308 155316 355320
rect 155368 355308 155374 355360
rect 120074 354696 120080 354748
rect 120132 354736 120138 354748
rect 203518 354736 203524 354748
rect 120132 354708 203524 354736
rect 120132 354696 120138 354708
rect 203518 354696 203524 354708
rect 203576 354696 203582 354748
rect 122650 353948 122656 354000
rect 122708 353988 122714 354000
rect 127618 353988 127624 354000
rect 122708 353960 127624 353988
rect 122708 353948 122714 353960
rect 127618 353948 127624 353960
rect 127676 353948 127682 354000
rect 60550 353336 60556 353388
rect 60608 353376 60614 353388
rect 162118 353376 162124 353388
rect 60608 353348 162124 353376
rect 60608 353336 60614 353348
rect 162118 353336 162124 353348
rect 162176 353336 162182 353388
rect 132402 353268 132408 353320
rect 132460 353308 132466 353320
rect 320174 353308 320180 353320
rect 132460 353280 320180 353308
rect 132460 353268 132466 353280
rect 320174 353268 320180 353280
rect 320232 353268 320238 353320
rect 54846 352520 54852 352572
rect 54904 352560 54910 352572
rect 86954 352560 86960 352572
rect 54904 352532 86960 352560
rect 54904 352520 54910 352532
rect 86954 352520 86960 352532
rect 87012 352520 87018 352572
rect 104802 352520 104808 352572
rect 104860 352560 104866 352572
rect 120718 352560 120724 352572
rect 104860 352532 120724 352560
rect 104860 352520 104866 352532
rect 120718 352520 120724 352532
rect 120776 352520 120782 352572
rect 89070 351976 89076 352028
rect 89128 352016 89134 352028
rect 92658 352016 92664 352028
rect 89128 351988 92664 352016
rect 89128 351976 89134 351988
rect 92658 351976 92664 351988
rect 92716 352016 92722 352028
rect 92716 351988 93854 352016
rect 92716 351976 92722 351988
rect 85482 351908 85488 351960
rect 85540 351948 85546 351960
rect 90358 351948 90364 351960
rect 85540 351920 90364 351948
rect 85540 351908 85546 351920
rect 90358 351908 90364 351920
rect 90416 351908 90422 351960
rect 93826 351948 93854 351988
rect 125502 351976 125508 352028
rect 125560 352016 125566 352028
rect 125686 352016 125692 352028
rect 125560 351988 125692 352016
rect 125560 351976 125566 351988
rect 125686 351976 125692 351988
rect 125744 351976 125750 352028
rect 144178 351976 144184 352028
rect 144236 352016 144242 352028
rect 146294 352016 146300 352028
rect 144236 351988 146300 352016
rect 144236 351976 144242 351988
rect 146294 351976 146300 351988
rect 146352 352016 146358 352028
rect 195238 352016 195244 352028
rect 146352 351988 195244 352016
rect 146352 351976 146358 351988
rect 195238 351976 195244 351988
rect 195296 351976 195302 352028
rect 251266 351948 251272 351960
rect 93826 351920 251272 351948
rect 251266 351908 251272 351920
rect 251324 351908 251330 351960
rect 88978 351840 88984 351892
rect 89036 351880 89042 351892
rect 129642 351880 129648 351892
rect 89036 351852 129648 351880
rect 89036 351840 89042 351852
rect 129642 351840 129648 351852
rect 129700 351840 129706 351892
rect 118786 350548 118792 350600
rect 118844 350588 118850 350600
rect 119338 350588 119344 350600
rect 118844 350560 119344 350588
rect 118844 350548 118850 350560
rect 119338 350548 119344 350560
rect 119396 350588 119402 350600
rect 249886 350588 249892 350600
rect 119396 350560 249892 350588
rect 119396 350548 119402 350560
rect 249886 350548 249892 350560
rect 249944 350548 249950 350600
rect 79962 349800 79968 349852
rect 80020 349840 80026 349852
rect 111334 349840 111340 349852
rect 80020 349812 111340 349840
rect 80020 349800 80026 349812
rect 111334 349800 111340 349812
rect 111392 349800 111398 349852
rect 112438 349800 112444 349852
rect 112496 349840 112502 349852
rect 156046 349840 156052 349852
rect 112496 349812 156052 349840
rect 112496 349800 112502 349812
rect 156046 349800 156052 349812
rect 156104 349800 156110 349852
rect 133874 349120 133880 349172
rect 133932 349160 133938 349172
rect 236638 349160 236644 349172
rect 133932 349132 236644 349160
rect 133932 349120 133938 349132
rect 236638 349120 236644 349132
rect 236696 349120 236702 349172
rect 83458 348372 83464 348424
rect 83516 348412 83522 348424
rect 109678 348412 109684 348424
rect 83516 348384 109684 348412
rect 83516 348372 83522 348384
rect 109678 348372 109684 348384
rect 109736 348372 109742 348424
rect 121638 347828 121644 347880
rect 121696 347868 121702 347880
rect 122742 347868 122748 347880
rect 121696 347840 122748 347868
rect 121696 347828 121702 347840
rect 122742 347828 122748 347840
rect 122800 347868 122806 347880
rect 196618 347868 196624 347880
rect 122800 347840 196624 347868
rect 122800 347828 122806 347840
rect 196618 347828 196624 347840
rect 196676 347828 196682 347880
rect 77202 347760 77208 347812
rect 77260 347800 77266 347812
rect 204346 347800 204352 347812
rect 77260 347772 204352 347800
rect 77260 347760 77266 347772
rect 204346 347760 204352 347772
rect 204404 347760 204410 347812
rect 79318 347692 79324 347744
rect 79376 347732 79382 347744
rect 121638 347732 121644 347744
rect 79376 347704 121644 347732
rect 79376 347692 79382 347704
rect 121638 347692 121644 347704
rect 121696 347692 121702 347744
rect 204162 347692 204168 347744
rect 204220 347732 204226 347744
rect 582374 347732 582380 347744
rect 204220 347704 582380 347732
rect 204220 347692 204226 347704
rect 582374 347692 582380 347704
rect 582432 347692 582438 347744
rect 152458 347080 152464 347132
rect 152516 347120 152522 347132
rect 161658 347120 161664 347132
rect 152516 347092 161664 347120
rect 152516 347080 152522 347092
rect 161658 347080 161664 347092
rect 161716 347080 161722 347132
rect 203058 347052 203064 347064
rect 93826 347024 203064 347052
rect 85574 346944 85580 346996
rect 85632 346984 85638 346996
rect 86310 346984 86316 346996
rect 85632 346956 86316 346984
rect 85632 346944 85638 346956
rect 86310 346944 86316 346956
rect 86368 346984 86374 346996
rect 93826 346984 93854 347024
rect 203058 347012 203064 347024
rect 203116 347052 203122 347064
rect 204162 347052 204168 347064
rect 203116 347024 204168 347052
rect 203116 347012 203122 347024
rect 204162 347012 204168 347024
rect 204220 347012 204226 347064
rect 86368 346956 93854 346984
rect 86368 346944 86374 346956
rect 2774 346264 2780 346316
rect 2832 346304 2838 346316
rect 4798 346304 4804 346316
rect 2832 346276 4804 346304
rect 2832 346264 2838 346276
rect 4798 346264 4804 346276
rect 4856 346264 4862 346316
rect 115198 345108 115204 345160
rect 115256 345148 115262 345160
rect 229186 345148 229192 345160
rect 115256 345120 229192 345148
rect 115256 345108 115262 345120
rect 229186 345108 229192 345120
rect 229244 345108 229250 345160
rect 91002 345040 91008 345092
rect 91060 345080 91066 345092
rect 210418 345080 210424 345092
rect 91060 345052 210424 345080
rect 91060 345040 91066 345052
rect 210418 345040 210424 345052
rect 210476 345040 210482 345092
rect 87966 343680 87972 343732
rect 88024 343720 88030 343732
rect 216030 343720 216036 343732
rect 88024 343692 216036 343720
rect 88024 343680 88030 343692
rect 216030 343680 216036 343692
rect 216088 343680 216094 343732
rect 73798 343612 73804 343664
rect 73856 343652 73862 343664
rect 209130 343652 209136 343664
rect 73856 343624 209136 343652
rect 73856 343612 73862 343624
rect 209130 343612 209136 343624
rect 209188 343612 209194 343664
rect 62022 342320 62028 342372
rect 62080 342360 62086 342372
rect 163682 342360 163688 342372
rect 62080 342332 163688 342360
rect 62080 342320 62086 342332
rect 163682 342320 163688 342332
rect 163740 342320 163746 342372
rect 93670 342252 93676 342304
rect 93728 342292 93734 342304
rect 252646 342292 252652 342304
rect 93728 342264 252652 342292
rect 93728 342252 93734 342264
rect 252646 342252 252652 342264
rect 252704 342252 252710 342304
rect 130010 340960 130016 341012
rect 130068 341000 130074 341012
rect 166258 341000 166264 341012
rect 130068 340972 166264 341000
rect 130068 340960 130074 340972
rect 166258 340960 166264 340972
rect 166316 340960 166322 341012
rect 102778 340892 102784 340944
rect 102836 340932 102842 340944
rect 258166 340932 258172 340944
rect 102836 340904 258172 340932
rect 102836 340892 102842 340904
rect 258166 340892 258172 340904
rect 258224 340892 258230 340944
rect 78490 340144 78496 340196
rect 78548 340184 78554 340196
rect 93118 340184 93124 340196
rect 78548 340156 93124 340184
rect 78548 340144 78554 340156
rect 93118 340144 93124 340156
rect 93176 340144 93182 340196
rect 114462 339532 114468 339584
rect 114520 339572 114526 339584
rect 169018 339572 169024 339584
rect 114520 339544 169024 339572
rect 114520 339532 114526 339544
rect 169018 339532 169024 339544
rect 169076 339532 169082 339584
rect 64690 339464 64696 339516
rect 64748 339504 64754 339516
rect 122190 339504 122196 339516
rect 64748 339476 122196 339504
rect 64748 339464 64754 339476
rect 122190 339464 122196 339476
rect 122248 339464 122254 339516
rect 132770 339464 132776 339516
rect 132828 339504 132834 339516
rect 259454 339504 259460 339516
rect 132828 339476 259460 339504
rect 132828 339464 132834 339476
rect 259454 339464 259460 339476
rect 259512 339464 259518 339516
rect 79870 338716 79876 338768
rect 79928 338756 79934 338768
rect 89070 338756 89076 338768
rect 79928 338728 89076 338756
rect 79928 338716 79934 338728
rect 89070 338716 89076 338728
rect 89128 338716 89134 338768
rect 67726 338512 67732 338564
rect 67784 338552 67790 338564
rect 72418 338552 72424 338564
rect 67784 338524 72424 338552
rect 67784 338512 67790 338524
rect 72418 338512 72424 338524
rect 72476 338512 72482 338564
rect 148410 338172 148416 338224
rect 148468 338212 148474 338224
rect 155218 338212 155224 338224
rect 148468 338184 155224 338212
rect 148468 338172 148474 338184
rect 155218 338172 155224 338184
rect 155276 338172 155282 338224
rect 106458 338104 106464 338156
rect 106516 338144 106522 338156
rect 184290 338144 184296 338156
rect 106516 338116 184296 338144
rect 106516 338104 106522 338116
rect 184290 338104 184296 338116
rect 184348 338104 184354 338156
rect 115934 336812 115940 336864
rect 115992 336852 115998 336864
rect 247034 336852 247040 336864
rect 115992 336824 247040 336852
rect 115992 336812 115998 336824
rect 247034 336812 247040 336824
rect 247092 336812 247098 336864
rect 67266 336744 67272 336796
rect 67324 336784 67330 336796
rect 206370 336784 206376 336796
rect 67324 336756 206376 336784
rect 67324 336744 67330 336756
rect 206370 336744 206376 336756
rect 206428 336744 206434 336796
rect 61838 335384 61844 335436
rect 61896 335424 61902 335436
rect 115290 335424 115296 335436
rect 61896 335396 115296 335424
rect 61896 335384 61902 335396
rect 115290 335384 115296 335396
rect 115348 335384 115354 335436
rect 127066 335384 127072 335436
rect 127124 335424 127130 335436
rect 182910 335424 182916 335436
rect 127124 335396 182916 335424
rect 127124 335384 127130 335396
rect 182910 335384 182916 335396
rect 182968 335384 182974 335436
rect 73154 335316 73160 335368
rect 73212 335356 73218 335368
rect 192478 335356 192484 335368
rect 73212 335328 192484 335356
rect 73212 335316 73218 335328
rect 192478 335316 192484 335328
rect 192536 335316 192542 335368
rect 76466 334636 76472 334688
rect 76524 334676 76530 334688
rect 87046 334676 87052 334688
rect 76524 334648 87052 334676
rect 76524 334636 76530 334648
rect 87046 334636 87052 334648
rect 87104 334636 87110 334688
rect 3418 334568 3424 334620
rect 3476 334608 3482 334620
rect 11698 334608 11704 334620
rect 3476 334580 11704 334608
rect 3476 334568 3482 334580
rect 11698 334568 11704 334580
rect 11756 334568 11762 334620
rect 67818 334568 67824 334620
rect 67876 334608 67882 334620
rect 115198 334608 115204 334620
rect 67876 334580 115204 334608
rect 67876 334568 67882 334580
rect 115198 334568 115204 334580
rect 115256 334568 115262 334620
rect 141326 334024 141332 334076
rect 141384 334064 141390 334076
rect 171778 334064 171784 334076
rect 141384 334036 171784 334064
rect 141384 334024 141390 334036
rect 171778 334024 171784 334036
rect 171836 334024 171842 334076
rect 101490 333956 101496 334008
rect 101548 333996 101554 334008
rect 159542 333996 159548 334008
rect 101548 333968 159548 333996
rect 101548 333956 101554 333968
rect 159542 333956 159548 333968
rect 159600 333956 159606 334008
rect 66162 333344 66168 333396
rect 66220 333384 66226 333396
rect 74534 333384 74540 333396
rect 66220 333356 74540 333384
rect 66220 333344 66226 333356
rect 74534 333344 74540 333356
rect 74592 333344 74598 333396
rect 75730 333208 75736 333260
rect 75788 333248 75794 333260
rect 101398 333248 101404 333260
rect 75788 333220 101404 333248
rect 75788 333208 75794 333220
rect 101398 333208 101404 333220
rect 101456 333208 101462 333260
rect 97258 332664 97264 332716
rect 97316 332704 97322 332716
rect 170398 332704 170404 332716
rect 97316 332676 170404 332704
rect 97316 332664 97322 332676
rect 170398 332664 170404 332676
rect 170456 332664 170462 332716
rect 115658 332596 115664 332648
rect 115716 332636 115722 332648
rect 198090 332636 198096 332648
rect 115716 332608 198096 332636
rect 115716 332596 115722 332608
rect 198090 332596 198096 332608
rect 198148 332596 198154 332648
rect 60458 331848 60464 331900
rect 60516 331888 60522 331900
rect 122098 331888 122104 331900
rect 60516 331860 122104 331888
rect 60516 331848 60522 331860
rect 122098 331848 122104 331860
rect 122156 331848 122162 331900
rect 133782 331304 133788 331356
rect 133840 331344 133846 331356
rect 195422 331344 195428 331356
rect 133840 331316 195428 331344
rect 133840 331304 133846 331316
rect 195422 331304 195428 331316
rect 195480 331304 195486 331356
rect 72234 331236 72240 331288
rect 72292 331276 72298 331288
rect 215938 331276 215944 331288
rect 72292 331248 215944 331276
rect 72292 331236 72298 331248
rect 215938 331236 215944 331248
rect 215996 331236 216002 331288
rect 59262 331168 59268 331220
rect 59320 331208 59326 331220
rect 99374 331208 99380 331220
rect 59320 331180 99380 331208
rect 59320 331168 59326 331180
rect 99374 331168 99380 331180
rect 99432 331168 99438 331220
rect 80698 331100 80704 331152
rect 80756 331140 80762 331152
rect 81342 331140 81348 331152
rect 80756 331112 81348 331140
rect 80756 331100 80762 331112
rect 81342 331100 81348 331112
rect 81400 331100 81406 331152
rect 82722 331100 82728 331152
rect 82780 331140 82786 331152
rect 83458 331140 83464 331152
rect 82780 331112 83464 331140
rect 82780 331100 82786 331112
rect 83458 331100 83464 331112
rect 83516 331100 83522 331152
rect 85574 331100 85580 331152
rect 85632 331140 85638 331152
rect 86586 331140 86592 331152
rect 85632 331112 86592 331140
rect 85632 331100 85638 331112
rect 86586 331100 86592 331112
rect 86644 331100 86650 331152
rect 114370 331100 114376 331152
rect 114428 331140 114434 331152
rect 114738 331140 114744 331152
rect 114428 331112 114744 331140
rect 114428 331100 114434 331112
rect 114738 331100 114744 331112
rect 114796 331100 114802 331152
rect 126974 331100 126980 331152
rect 127032 331140 127038 331152
rect 127894 331140 127900 331152
rect 127032 331112 127900 331140
rect 127032 331100 127038 331112
rect 127894 331100 127900 331112
rect 127952 331100 127958 331152
rect 137830 331100 137836 331152
rect 137888 331140 137894 331152
rect 139394 331140 139400 331152
rect 137888 331112 139400 331140
rect 137888 331100 137894 331112
rect 139394 331100 139400 331112
rect 139452 331100 139458 331152
rect 70670 330760 70676 330812
rect 70728 330800 70734 330812
rect 73798 330800 73804 330812
rect 70728 330772 73804 330800
rect 70728 330760 70734 330772
rect 73798 330760 73804 330772
rect 73856 330760 73862 330812
rect 122098 330556 122104 330608
rect 122156 330596 122162 330608
rect 137278 330596 137284 330608
rect 122156 330568 137284 330596
rect 122156 330556 122162 330568
rect 137278 330556 137284 330568
rect 137336 330556 137342 330608
rect 17218 330488 17224 330540
rect 17276 330528 17282 330540
rect 59262 330528 59268 330540
rect 17276 330500 59268 330528
rect 17276 330488 17282 330500
rect 59262 330488 59268 330500
rect 59320 330488 59326 330540
rect 96430 330488 96436 330540
rect 96488 330528 96494 330540
rect 124858 330528 124864 330540
rect 96488 330500 124864 330528
rect 96488 330488 96494 330500
rect 124858 330488 124864 330500
rect 124916 330488 124922 330540
rect 178770 330488 178776 330540
rect 178828 330528 178834 330540
rect 228358 330528 228364 330540
rect 178828 330500 228364 330528
rect 178828 330488 178834 330500
rect 228358 330488 228364 330500
rect 228416 330488 228422 330540
rect 98546 330352 98552 330404
rect 98604 330392 98610 330404
rect 99282 330392 99288 330404
rect 98604 330364 99288 330392
rect 98604 330352 98610 330364
rect 99282 330352 99288 330364
rect 99340 330352 99346 330404
rect 77938 330216 77944 330268
rect 77996 330256 78002 330268
rect 78582 330256 78588 330268
rect 77996 330228 78588 330256
rect 77996 330216 78002 330228
rect 78582 330216 78588 330228
rect 78640 330216 78646 330268
rect 79410 330216 79416 330268
rect 79468 330256 79474 330268
rect 79962 330256 79968 330268
rect 79468 330228 79968 330256
rect 79468 330216 79474 330228
rect 79962 330216 79968 330228
rect 80020 330216 80026 330268
rect 117774 330216 117780 330268
rect 117832 330256 117838 330268
rect 118602 330256 118608 330268
rect 117832 330228 118608 330256
rect 117832 330216 117838 330228
rect 118602 330216 118608 330228
rect 118660 330216 118666 330268
rect 110598 330080 110604 330132
rect 110656 330120 110662 330132
rect 111702 330120 111708 330132
rect 110656 330092 111708 330120
rect 110656 330080 110662 330092
rect 111702 330080 111708 330092
rect 111760 330080 111766 330132
rect 92842 330012 92848 330064
rect 92900 330052 92906 330064
rect 93762 330052 93768 330064
rect 92900 330024 93768 330052
rect 92900 330012 92906 330024
rect 93762 330012 93768 330024
rect 93820 330012 93826 330064
rect 74166 329944 74172 329996
rect 74224 329984 74230 329996
rect 76558 329984 76564 329996
rect 74224 329956 76564 329984
rect 74224 329944 74230 329956
rect 76558 329944 76564 329956
rect 76616 329944 76622 329996
rect 95786 329944 95792 329996
rect 95844 329984 95850 329996
rect 96522 329984 96528 329996
rect 95844 329956 96528 329984
rect 95844 329944 95850 329956
rect 96522 329944 96528 329956
rect 96580 329944 96586 329996
rect 113634 329944 113640 329996
rect 113692 329984 113698 329996
rect 114462 329984 114468 329996
rect 113692 329956 114468 329984
rect 113692 329944 113698 329956
rect 114462 329944 114468 329956
rect 114520 329944 114526 329996
rect 147582 329944 147588 329996
rect 147640 329984 147646 329996
rect 177298 329984 177304 329996
rect 147640 329956 177304 329984
rect 147640 329944 147646 329956
rect 177298 329944 177304 329956
rect 177356 329944 177362 329996
rect 132678 329876 132684 329928
rect 132736 329916 132742 329928
rect 132736 329888 135944 329916
rect 132736 329876 132742 329888
rect 44082 329808 44088 329860
rect 44140 329848 44146 329860
rect 69106 329848 69112 329860
rect 44140 329820 69112 329848
rect 44140 329808 44146 329820
rect 69106 329808 69112 329820
rect 69164 329808 69170 329860
rect 99374 329808 99380 329860
rect 99432 329848 99438 329860
rect 100110 329848 100116 329860
rect 99432 329820 100116 329848
rect 99432 329808 99438 329820
rect 100110 329808 100116 329820
rect 100168 329808 100174 329860
rect 104158 329808 104164 329860
rect 104216 329848 104222 329860
rect 105538 329848 105544 329860
rect 104216 329820 105544 329848
rect 104216 329808 104222 329820
rect 105538 329808 105544 329820
rect 105596 329808 105602 329860
rect 108574 329808 108580 329860
rect 108632 329848 108638 329860
rect 108942 329848 108948 329860
rect 108632 329820 108948 329848
rect 108632 329808 108638 329820
rect 108942 329808 108948 329820
rect 109000 329808 109006 329860
rect 131482 329808 131488 329860
rect 131540 329848 131546 329860
rect 132402 329848 132408 329860
rect 131540 329820 132408 329848
rect 131540 329808 131546 329820
rect 132402 329808 132408 329820
rect 132460 329808 132466 329860
rect 134150 329808 134156 329860
rect 134208 329848 134214 329860
rect 135162 329848 135168 329860
rect 134208 329820 135168 329848
rect 134208 329808 134214 329820
rect 135162 329808 135168 329820
rect 135220 329808 135226 329860
rect 135254 329808 135260 329860
rect 135312 329848 135318 329860
rect 135806 329848 135812 329860
rect 135312 329820 135812 329848
rect 135312 329808 135318 329820
rect 135806 329808 135812 329820
rect 135864 329808 135870 329860
rect 135916 329848 135944 329888
rect 136910 329876 136916 329928
rect 136968 329916 136974 329928
rect 137922 329916 137928 329928
rect 136968 329888 137928 329916
rect 136968 329876 136974 329888
rect 137922 329876 137928 329888
rect 137980 329876 137986 329928
rect 143534 329916 143540 329928
rect 140608 329888 143540 329916
rect 140608 329848 140636 329888
rect 143534 329876 143540 329888
rect 143592 329876 143598 329928
rect 135916 329820 140636 329848
rect 140682 329808 140688 329860
rect 140740 329848 140746 329860
rect 141418 329848 141424 329860
rect 140740 329820 141424 329848
rect 140740 329808 140746 329820
rect 141418 329808 141424 329820
rect 141476 329808 141482 329860
rect 153286 329808 153292 329860
rect 153344 329848 153350 329860
rect 159358 329848 159364 329860
rect 153344 329820 159364 329848
rect 153344 329808 153350 329820
rect 159358 329808 159364 329820
rect 159416 329808 159422 329860
rect 122190 329740 122196 329792
rect 122248 329780 122254 329792
rect 133782 329780 133788 329792
rect 122248 329752 133788 329780
rect 122248 329740 122254 329752
rect 133782 329740 133788 329752
rect 133840 329740 133846 329792
rect 166902 329128 166908 329180
rect 166960 329168 166966 329180
rect 179414 329168 179420 329180
rect 166960 329140 179420 329168
rect 166960 329128 166966 329140
rect 179414 329128 179420 329140
rect 179472 329128 179478 329180
rect 188522 329128 188528 329180
rect 188580 329168 188586 329180
rect 211890 329168 211896 329180
rect 188580 329140 211896 329168
rect 188580 329128 188586 329140
rect 211890 329128 211896 329140
rect 211948 329128 211954 329180
rect 241238 329128 241244 329180
rect 241296 329168 241302 329180
rect 306374 329168 306380 329180
rect 241296 329140 306380 329168
rect 241296 329128 241302 329140
rect 306374 329128 306380 329140
rect 306432 329128 306438 329180
rect 36538 329060 36544 329112
rect 36596 329100 36602 329112
rect 49602 329100 49608 329112
rect 36596 329072 49608 329100
rect 36596 329060 36602 329072
rect 49602 329060 49608 329072
rect 49660 329100 49666 329112
rect 135254 329100 135260 329112
rect 49660 329072 135260 329100
rect 49660 329060 49666 329072
rect 135254 329060 135260 329072
rect 135312 329060 135318 329112
rect 150342 329060 150348 329112
rect 150400 329100 150406 329112
rect 248598 329100 248604 329112
rect 150400 329072 248604 329100
rect 150400 329060 150406 329072
rect 248598 329060 248604 329072
rect 248656 329060 248662 329112
rect 144822 328448 144828 328500
rect 144880 328488 144886 328500
rect 158162 328488 158168 328500
rect 144880 328460 158168 328488
rect 144880 328448 144886 328460
rect 158162 328448 158168 328460
rect 158220 328448 158226 328500
rect 115290 328380 115296 328432
rect 115348 328420 115354 328432
rect 141970 328420 141976 328432
rect 115348 328392 141976 328420
rect 115348 328380 115354 328392
rect 141970 328380 141976 328392
rect 142028 328380 142034 328432
rect 67358 327768 67364 327820
rect 67416 327808 67422 327820
rect 91738 327808 91744 327820
rect 67416 327780 91744 327808
rect 67416 327768 67422 327780
rect 91738 327768 91744 327780
rect 91796 327768 91802 327820
rect 65886 327700 65892 327752
rect 65944 327740 65950 327752
rect 133874 327740 133880 327752
rect 65944 327712 133880 327740
rect 65944 327700 65950 327712
rect 133874 327700 133880 327712
rect 133932 327700 133938 327752
rect 179414 327700 179420 327752
rect 179472 327740 179478 327752
rect 192846 327740 192852 327752
rect 179472 327712 192852 327740
rect 179472 327700 179478 327712
rect 192846 327700 192852 327712
rect 192904 327700 192910 327752
rect 148594 327224 148600 327276
rect 148652 327264 148658 327276
rect 152918 327264 152924 327276
rect 148652 327236 152924 327264
rect 148652 327224 148658 327236
rect 152918 327224 152924 327236
rect 152976 327224 152982 327276
rect 152090 327156 152096 327208
rect 152148 327196 152154 327208
rect 160830 327196 160836 327208
rect 152148 327168 160836 327196
rect 152148 327156 152154 327168
rect 160830 327156 160836 327168
rect 160888 327156 160894 327208
rect 135530 327088 135536 327140
rect 135588 327128 135594 327140
rect 249794 327128 249800 327140
rect 135588 327100 249800 327128
rect 135588 327088 135594 327100
rect 249794 327088 249800 327100
rect 249852 327088 249858 327140
rect 55950 327020 55956 327072
rect 56008 327060 56014 327072
rect 56502 327060 56508 327072
rect 56008 327032 56508 327060
rect 56008 327020 56014 327032
rect 56502 327020 56508 327032
rect 56560 327060 56566 327072
rect 93854 327060 93860 327072
rect 56560 327032 93860 327060
rect 56560 327020 56566 327032
rect 93854 327020 93860 327032
rect 93912 327020 93918 327072
rect 143534 327020 143540 327072
rect 143592 327060 143598 327072
rect 154850 327060 154856 327072
rect 143592 327032 154856 327060
rect 143592 327020 143598 327032
rect 154850 327020 154856 327032
rect 154908 327020 154914 327072
rect 69934 326952 69940 327004
rect 69992 326992 69998 327004
rect 71038 326992 71044 327004
rect 69992 326964 71044 326992
rect 69992 326952 69998 326964
rect 71038 326952 71044 326964
rect 71096 326952 71102 327004
rect 152918 326884 152924 326936
rect 152976 326884 152982 326936
rect 154298 326884 154304 326936
rect 154356 326924 154362 326936
rect 155218 326924 155224 326936
rect 154356 326896 155224 326924
rect 154356 326884 154362 326896
rect 155218 326884 155224 326896
rect 155276 326884 155282 326936
rect 14 326340 20 326392
rect 72 326380 78 326392
rect 55950 326380 55956 326392
rect 72 326352 55956 326380
rect 72 326340 78 326352
rect 55950 326340 55956 326352
rect 56008 326340 56014 326392
rect 152936 326380 152964 326884
rect 159634 326408 159640 326460
rect 159692 326448 159698 326460
rect 199378 326448 199384 326460
rect 159692 326420 199384 326448
rect 159692 326408 159698 326420
rect 199378 326408 199384 326420
rect 199436 326408 199442 326460
rect 196710 326380 196716 326392
rect 152936 326352 196716 326380
rect 196710 326340 196716 326352
rect 196768 326340 196774 326392
rect 203518 326340 203524 326392
rect 203576 326380 203582 326392
rect 228450 326380 228456 326392
rect 203576 326352 228456 326380
rect 203576 326340 203582 326352
rect 228450 326340 228456 326352
rect 228508 326340 228514 326392
rect 156046 326000 156052 326052
rect 156104 326040 156110 326052
rect 159450 326040 159456 326052
rect 156104 326012 159456 326040
rect 156104 326000 156110 326012
rect 159450 326000 159456 326012
rect 159508 326000 159514 326052
rect 156138 324980 156144 325032
rect 156196 325020 156202 325032
rect 255498 325020 255504 325032
rect 156196 324992 255504 325020
rect 156196 324980 156202 324992
rect 255498 324980 255504 324992
rect 255556 324980 255562 325032
rect 181622 324912 181628 324964
rect 181680 324952 181686 324964
rect 313918 324952 313924 324964
rect 181680 324924 313924 324952
rect 181680 324912 181686 324924
rect 313918 324912 313924 324924
rect 313976 324912 313982 324964
rect 59262 324300 59268 324352
rect 59320 324340 59326 324352
rect 66806 324340 66812 324352
rect 59320 324312 66812 324340
rect 59320 324300 59326 324312
rect 66806 324300 66812 324312
rect 66864 324300 66870 324352
rect 159542 323620 159548 323672
rect 159600 323660 159606 323672
rect 220814 323660 220820 323672
rect 159600 323632 220820 323660
rect 159600 323620 159606 323632
rect 220814 323620 220820 323632
rect 220872 323620 220878 323672
rect 160922 323552 160928 323604
rect 160980 323592 160986 323604
rect 349154 323592 349160 323604
rect 160980 323564 349160 323592
rect 160980 323552 160986 323564
rect 349154 323552 349160 323564
rect 349212 323552 349218 323604
rect 61930 322940 61936 322992
rect 61988 322980 61994 322992
rect 66806 322980 66812 322992
rect 61988 322952 66812 322980
rect 61988 322940 61994 322952
rect 66806 322940 66812 322952
rect 66864 322940 66870 322992
rect 156046 322940 156052 322992
rect 156104 322980 156110 322992
rect 161014 322980 161020 322992
rect 156104 322952 161020 322980
rect 156104 322940 156110 322952
rect 161014 322940 161020 322952
rect 161072 322940 161078 322992
rect 230474 322464 230480 322516
rect 230532 322504 230538 322516
rect 236730 322504 236736 322516
rect 230532 322476 236736 322504
rect 230532 322464 230538 322476
rect 236730 322464 236736 322476
rect 236788 322464 236794 322516
rect 185762 322260 185768 322312
rect 185820 322300 185826 322312
rect 202874 322300 202880 322312
rect 185820 322272 202880 322300
rect 185820 322260 185826 322272
rect 202874 322260 202880 322272
rect 202932 322260 202938 322312
rect 166258 322192 166264 322244
rect 166316 322232 166322 322244
rect 232498 322232 232504 322244
rect 166316 322204 232504 322232
rect 166316 322192 166322 322204
rect 232498 322192 232504 322204
rect 232556 322192 232562 322244
rect 156046 321580 156052 321632
rect 156104 321620 156110 321632
rect 166442 321620 166448 321632
rect 156104 321592 166448 321620
rect 156104 321580 156110 321592
rect 166442 321580 166448 321592
rect 166500 321580 166506 321632
rect 193858 320900 193864 320952
rect 193916 320940 193922 320952
rect 235258 320940 235264 320952
rect 193916 320912 235264 320940
rect 193916 320900 193922 320912
rect 235258 320900 235264 320912
rect 235316 320900 235322 320952
rect 156966 320832 156972 320884
rect 157024 320872 157030 320884
rect 233878 320872 233884 320884
rect 157024 320844 233884 320872
rect 157024 320832 157030 320844
rect 233878 320832 233884 320844
rect 233936 320832 233942 320884
rect 157242 319948 157248 320000
rect 157300 319988 157306 320000
rect 161566 319988 161572 320000
rect 157300 319960 161572 319988
rect 157300 319948 157306 319960
rect 161566 319948 161572 319960
rect 161624 319988 161630 320000
rect 162210 319988 162216 320000
rect 161624 319960 162216 319988
rect 161624 319948 161630 319960
rect 162210 319948 162216 319960
rect 162268 319948 162274 320000
rect 4062 319404 4068 319456
rect 4120 319444 4126 319456
rect 15838 319444 15844 319456
rect 4120 319416 15844 319444
rect 4120 319404 4126 319416
rect 15838 319404 15844 319416
rect 15896 319404 15902 319456
rect 171778 319404 171784 319456
rect 171836 319444 171842 319456
rect 248506 319444 248512 319456
rect 171836 319416 248512 319444
rect 171836 319404 171842 319416
rect 248506 319404 248512 319416
rect 248564 319404 248570 319456
rect 56502 318792 56508 318844
rect 56560 318832 56566 318844
rect 66254 318832 66260 318844
rect 56560 318804 66260 318832
rect 56560 318792 56566 318804
rect 66254 318792 66260 318804
rect 66312 318792 66318 318844
rect 157242 318792 157248 318844
rect 157300 318832 157306 318844
rect 178862 318832 178868 318844
rect 157300 318804 178868 318832
rect 157300 318792 157306 318804
rect 178862 318792 178868 318804
rect 178920 318792 178926 318844
rect 215846 318724 215852 318776
rect 215904 318764 215910 318776
rect 216030 318764 216036 318776
rect 215904 318736 216036 318764
rect 215904 318724 215910 318736
rect 216030 318724 216036 318736
rect 216088 318724 216094 318776
rect 166350 318112 166356 318164
rect 166408 318152 166414 318164
rect 202782 318152 202788 318164
rect 166408 318124 202788 318152
rect 166408 318112 166414 318124
rect 202782 318112 202788 318124
rect 202840 318112 202846 318164
rect 11698 318044 11704 318096
rect 11756 318084 11762 318096
rect 46842 318084 46848 318096
rect 11756 318056 46848 318084
rect 11756 318044 11762 318056
rect 46842 318044 46848 318056
rect 46900 318044 46906 318096
rect 184198 318044 184204 318096
rect 184256 318084 184262 318096
rect 227070 318084 227076 318096
rect 184256 318056 227076 318084
rect 184256 318044 184262 318056
rect 227070 318044 227076 318056
rect 227128 318044 227134 318096
rect 60642 317500 60648 317552
rect 60700 317540 60706 317552
rect 66254 317540 66260 317552
rect 60700 317512 66260 317540
rect 60700 317500 60706 317512
rect 66254 317500 66260 317512
rect 66312 317500 66318 317552
rect 46842 317432 46848 317484
rect 46900 317472 46906 317484
rect 66346 317472 66352 317484
rect 46900 317444 66352 317472
rect 46900 317432 46906 317444
rect 66346 317432 66352 317444
rect 66404 317432 66410 317484
rect 215846 317432 215852 317484
rect 215904 317472 215910 317484
rect 300946 317472 300952 317484
rect 215904 317444 300952 317472
rect 215904 317432 215910 317444
rect 300946 317432 300952 317444
rect 301004 317432 301010 317484
rect 157242 316684 157248 316736
rect 157300 316724 157306 316736
rect 189810 316724 189816 316736
rect 157300 316696 189816 316724
rect 157300 316684 157306 316696
rect 189810 316684 189816 316696
rect 189868 316684 189874 316736
rect 156690 316004 156696 316056
rect 156748 316044 156754 316056
rect 254026 316044 254032 316056
rect 156748 316016 254032 316044
rect 156748 316004 156754 316016
rect 254026 316004 254032 316016
rect 254084 316004 254090 316056
rect 61838 315936 61844 315988
rect 61896 315976 61902 315988
rect 66990 315976 66996 315988
rect 61896 315948 66996 315976
rect 61896 315936 61902 315948
rect 66990 315936 66996 315948
rect 67048 315936 67054 315988
rect 157242 315936 157248 315988
rect 157300 315976 157306 315988
rect 166994 315976 167000 315988
rect 157300 315948 167000 315976
rect 157300 315936 157306 315948
rect 166994 315936 167000 315948
rect 167052 315936 167058 315988
rect 236730 315324 236736 315376
rect 236788 315364 236794 315376
rect 242894 315364 242900 315376
rect 236788 315336 242900 315364
rect 236788 315324 236794 315336
rect 242894 315324 242900 315336
rect 242952 315324 242958 315376
rect 166994 315256 167000 315308
rect 167052 315296 167058 315308
rect 178770 315296 178776 315308
rect 167052 315268 178776 315296
rect 167052 315256 167058 315268
rect 178770 315256 178776 315268
rect 178828 315256 178834 315308
rect 178862 315256 178868 315308
rect 178920 315296 178926 315308
rect 245746 315296 245752 315308
rect 178920 315268 245752 315296
rect 178920 315256 178926 315268
rect 245746 315256 245752 315268
rect 245804 315256 245810 315308
rect 35250 314644 35256 314696
rect 35308 314684 35314 314696
rect 66438 314684 66444 314696
rect 35308 314656 66444 314684
rect 35308 314644 35314 314656
rect 66438 314644 66444 314656
rect 66496 314644 66502 314696
rect 61838 314168 61844 314220
rect 61896 314208 61902 314220
rect 66254 314208 66260 314220
rect 61896 314180 66260 314208
rect 61896 314168 61902 314180
rect 66254 314168 66260 314180
rect 66312 314168 66318 314220
rect 195422 313896 195428 313948
rect 195480 313936 195486 313948
rect 225046 313936 225052 313948
rect 195480 313908 225052 313936
rect 195480 313896 195486 313908
rect 225046 313896 225052 313908
rect 225104 313896 225110 313948
rect 60550 313216 60556 313268
rect 60608 313256 60614 313268
rect 66254 313256 66260 313268
rect 60608 313228 66260 313256
rect 60608 313216 60614 313228
rect 66254 313216 66260 313228
rect 66312 313216 66318 313268
rect 52270 312536 52276 312588
rect 52328 312576 52334 312588
rect 61102 312576 61108 312588
rect 52328 312548 61108 312576
rect 52328 312536 52334 312548
rect 61102 312536 61108 312548
rect 61160 312536 61166 312588
rect 157150 312536 157156 312588
rect 157208 312576 157214 312588
rect 244274 312576 244280 312588
rect 157208 312548 244280 312576
rect 157208 312536 157214 312548
rect 244274 312536 244280 312548
rect 244332 312536 244338 312588
rect 157242 311856 157248 311908
rect 157300 311896 157306 311908
rect 193858 311896 193864 311908
rect 157300 311868 193864 311896
rect 157300 311856 157306 311868
rect 193858 311856 193864 311868
rect 193916 311856 193922 311908
rect 207566 311856 207572 311908
rect 207624 311896 207630 311908
rect 282178 311896 282184 311908
rect 207624 311868 282184 311896
rect 207624 311856 207630 311868
rect 282178 311856 282184 311868
rect 282236 311856 282242 311908
rect 62022 311788 62028 311840
rect 62080 311828 62086 311840
rect 66806 311828 66812 311840
rect 62080 311800 66812 311828
rect 62080 311788 62086 311800
rect 66806 311788 66812 311800
rect 66864 311788 66870 311840
rect 181530 311176 181536 311228
rect 181588 311216 181594 311228
rect 230474 311216 230480 311228
rect 181588 311188 230480 311216
rect 181588 311176 181594 311188
rect 230474 311176 230480 311188
rect 230532 311176 230538 311228
rect 161014 311108 161020 311160
rect 161072 311148 161078 311160
rect 210510 311148 210516 311160
rect 161072 311120 210516 311148
rect 161072 311108 161078 311120
rect 210510 311108 210516 311120
rect 210568 311108 210574 311160
rect 218698 311108 218704 311160
rect 218756 311148 218762 311160
rect 309134 311148 309140 311160
rect 218756 311120 309140 311148
rect 218756 311108 218762 311120
rect 309134 311108 309140 311120
rect 309192 311108 309198 311160
rect 157242 310496 157248 310548
rect 157300 310536 157306 310548
rect 166350 310536 166356 310548
rect 157300 310508 166356 310536
rect 157300 310496 157306 310508
rect 166350 310496 166356 310508
rect 166408 310496 166414 310548
rect 201678 310360 201684 310412
rect 201736 310400 201742 310412
rect 202138 310400 202144 310412
rect 201736 310372 202144 310400
rect 201736 310360 201742 310372
rect 202138 310360 202144 310372
rect 202196 310360 202202 310412
rect 160830 309748 160836 309800
rect 160888 309788 160894 309800
rect 244550 309788 244556 309800
rect 160888 309760 244556 309788
rect 160888 309748 160894 309760
rect 244550 309748 244556 309760
rect 244608 309748 244614 309800
rect 67082 309408 67088 309460
rect 67140 309448 67146 309460
rect 67450 309448 67456 309460
rect 67140 309420 67456 309448
rect 67140 309408 67146 309420
rect 67450 309408 67456 309420
rect 67508 309408 67514 309460
rect 53558 309136 53564 309188
rect 53616 309176 53622 309188
rect 66622 309176 66628 309188
rect 53616 309148 66628 309176
rect 53616 309136 53622 309148
rect 66622 309136 66628 309148
rect 66680 309136 66686 309188
rect 157150 309136 157156 309188
rect 157208 309176 157214 309188
rect 177574 309176 177580 309188
rect 157208 309148 177580 309176
rect 157208 309136 157214 309148
rect 177574 309136 177580 309148
rect 177632 309136 177638 309188
rect 201678 309136 201684 309188
rect 201736 309176 201742 309188
rect 580258 309176 580264 309188
rect 201736 309148 580264 309176
rect 201736 309136 201742 309148
rect 580258 309136 580264 309148
rect 580316 309136 580322 309188
rect 157242 309068 157248 309120
rect 157300 309108 157306 309120
rect 172514 309108 172520 309120
rect 157300 309080 172520 309108
rect 157300 309068 157306 309080
rect 172514 309068 172520 309080
rect 172572 309108 172578 309120
rect 173802 309108 173808 309120
rect 172572 309080 173808 309108
rect 172572 309068 172578 309080
rect 173802 309068 173808 309080
rect 173860 309068 173866 309120
rect 214650 309068 214656 309120
rect 214708 309108 214714 309120
rect 215202 309108 215208 309120
rect 214708 309080 215208 309108
rect 214708 309068 214714 309080
rect 215202 309068 215208 309080
rect 215260 309068 215266 309120
rect 231210 309068 231216 309120
rect 231268 309108 231274 309120
rect 236730 309108 236736 309120
rect 231268 309080 236736 309108
rect 231268 309068 231274 309080
rect 236730 309068 236736 309080
rect 236788 309068 236794 309120
rect 49602 308388 49608 308440
rect 49660 308428 49666 308440
rect 67082 308428 67088 308440
rect 49660 308400 67088 308428
rect 49660 308388 49666 308400
rect 67082 308388 67088 308400
rect 67140 308388 67146 308440
rect 173802 308388 173808 308440
rect 173860 308428 173866 308440
rect 187050 308428 187056 308440
rect 173860 308400 187056 308428
rect 173860 308388 173866 308400
rect 187050 308388 187056 308400
rect 187108 308388 187114 308440
rect 18598 307776 18604 307828
rect 18656 307816 18662 307828
rect 49602 307816 49608 307828
rect 18656 307788 49608 307816
rect 18656 307776 18662 307788
rect 49602 307776 49608 307788
rect 49660 307776 49666 307828
rect 215202 307776 215208 307828
rect 215260 307816 215266 307828
rect 273898 307816 273904 307828
rect 215260 307788 273904 307816
rect 215260 307776 215266 307788
rect 273898 307776 273904 307788
rect 273956 307776 273962 307828
rect 65886 307708 65892 307760
rect 65944 307748 65950 307760
rect 67082 307748 67088 307760
rect 65944 307720 67088 307748
rect 65944 307708 65950 307720
rect 67082 307708 67088 307720
rect 67140 307708 67146 307760
rect 39298 307028 39304 307080
rect 39356 307068 39362 307080
rect 67174 307068 67180 307080
rect 39356 307040 67180 307068
rect 39356 307028 39362 307040
rect 67174 307028 67180 307040
rect 67232 307028 67238 307080
rect 164970 306892 164976 306944
rect 165028 306932 165034 306944
rect 171778 306932 171784 306944
rect 165028 306904 171784 306932
rect 165028 306892 165034 306904
rect 171778 306892 171784 306904
rect 171836 306892 171842 306944
rect 232498 306416 232504 306468
rect 232556 306456 232562 306468
rect 271138 306456 271144 306468
rect 232556 306428 271144 306456
rect 232556 306416 232562 306428
rect 271138 306416 271144 306428
rect 271196 306416 271202 306468
rect 173158 306348 173164 306400
rect 173216 306388 173222 306400
rect 247310 306388 247316 306400
rect 173216 306360 247316 306388
rect 173216 306348 173222 306360
rect 247310 306348 247316 306360
rect 247368 306348 247374 306400
rect 3418 306280 3424 306332
rect 3476 306320 3482 306332
rect 36538 306320 36544 306332
rect 3476 306292 36544 306320
rect 3476 306280 3482 306292
rect 36538 306280 36544 306292
rect 36596 306280 36602 306332
rect 157242 306280 157248 306332
rect 157300 306320 157306 306332
rect 160094 306320 160100 306332
rect 157300 306292 160100 306320
rect 157300 306280 157306 306292
rect 160094 306280 160100 306292
rect 160152 306280 160158 306332
rect 233970 305804 233976 305856
rect 234028 305844 234034 305856
rect 234522 305844 234528 305856
rect 234028 305816 234528 305844
rect 234028 305804 234034 305816
rect 234522 305804 234528 305816
rect 234580 305804 234586 305856
rect 170398 305600 170404 305652
rect 170456 305640 170462 305652
rect 192662 305640 192668 305652
rect 170456 305612 192668 305640
rect 170456 305600 170462 305612
rect 192662 305600 192668 305612
rect 192720 305600 192726 305652
rect 191098 305260 191104 305312
rect 191156 305300 191162 305312
rect 191650 305300 191656 305312
rect 191156 305272 191656 305300
rect 191156 305260 191162 305272
rect 191650 305260 191656 305272
rect 191708 305260 191714 305312
rect 157242 305192 157248 305244
rect 157300 305232 157306 305244
rect 162118 305232 162124 305244
rect 157300 305204 162124 305232
rect 157300 305192 157306 305204
rect 162118 305192 162124 305204
rect 162176 305192 162182 305244
rect 234522 305056 234528 305108
rect 234580 305096 234586 305108
rect 287330 305096 287336 305108
rect 234580 305068 287336 305096
rect 234580 305056 234586 305068
rect 287330 305056 287336 305068
rect 287388 305056 287394 305108
rect 191650 304988 191656 305040
rect 191708 305028 191714 305040
rect 261570 305028 261576 305040
rect 191708 305000 261576 305028
rect 191708 304988 191714 305000
rect 261570 304988 261576 305000
rect 261628 304988 261634 305040
rect 160094 304240 160100 304292
rect 160152 304280 160158 304292
rect 181622 304280 181628 304292
rect 160152 304252 181628 304280
rect 160152 304240 160158 304252
rect 181622 304240 181628 304252
rect 181680 304240 181686 304292
rect 222838 304240 222844 304292
rect 222896 304280 222902 304292
rect 232498 304280 232504 304292
rect 222896 304252 232504 304280
rect 222896 304240 222902 304252
rect 232498 304240 232504 304252
rect 232556 304240 232562 304292
rect 238662 304240 238668 304292
rect 238720 304280 238726 304292
rect 299566 304280 299572 304292
rect 238720 304252 299572 304280
rect 238720 304240 238726 304252
rect 299566 304240 299572 304252
rect 299624 304240 299630 304292
rect 156046 303628 156052 303680
rect 156104 303668 156110 303680
rect 204990 303668 204996 303680
rect 156104 303640 204996 303668
rect 156104 303628 156110 303640
rect 204990 303628 204996 303640
rect 205048 303628 205054 303680
rect 206370 303628 206376 303680
rect 206428 303668 206434 303680
rect 207014 303668 207020 303680
rect 206428 303640 207020 303668
rect 206428 303628 206434 303640
rect 207014 303628 207020 303640
rect 207072 303668 207078 303680
rect 256694 303668 256700 303680
rect 207072 303640 256700 303668
rect 207072 303628 207078 303640
rect 256694 303628 256700 303640
rect 256752 303628 256758 303680
rect 163590 302880 163596 302932
rect 163648 302920 163654 302932
rect 176102 302920 176108 302932
rect 163648 302892 176108 302920
rect 163648 302880 163654 302892
rect 176102 302880 176108 302892
rect 176160 302880 176166 302932
rect 222930 302268 222936 302320
rect 222988 302308 222994 302320
rect 223482 302308 223488 302320
rect 222988 302280 223488 302308
rect 222988 302268 222994 302280
rect 223482 302268 223488 302280
rect 223540 302308 223546 302320
rect 261478 302308 261484 302320
rect 223540 302280 261484 302308
rect 223540 302268 223546 302280
rect 261478 302268 261484 302280
rect 261536 302268 261542 302320
rect 157242 302200 157248 302252
rect 157300 302240 157306 302252
rect 165522 302240 165528 302252
rect 157300 302212 165528 302240
rect 157300 302200 157306 302212
rect 165522 302200 165528 302212
rect 165580 302200 165586 302252
rect 167638 302200 167644 302252
rect 167696 302240 167702 302252
rect 255590 302240 255596 302252
rect 167696 302212 255596 302240
rect 167696 302200 167702 302212
rect 255590 302200 255596 302212
rect 255648 302200 255654 302252
rect 64690 302132 64696 302184
rect 64748 302172 64754 302184
rect 66806 302172 66812 302184
rect 64748 302144 66812 302172
rect 64748 302132 64754 302144
rect 66806 302132 66812 302144
rect 66864 302132 66870 302184
rect 199378 302132 199384 302184
rect 199436 302172 199442 302184
rect 200574 302172 200580 302184
rect 199436 302144 200580 302172
rect 199436 302132 199442 302144
rect 200574 302132 200580 302144
rect 200632 302132 200638 302184
rect 170490 300908 170496 300960
rect 170548 300948 170554 300960
rect 241422 300948 241428 300960
rect 170548 300920 241428 300948
rect 170548 300908 170554 300920
rect 241422 300908 241428 300920
rect 241480 300908 241486 300960
rect 200114 300840 200120 300892
rect 200172 300880 200178 300892
rect 200574 300880 200580 300892
rect 200172 300852 200580 300880
rect 200172 300840 200178 300852
rect 200574 300840 200580 300852
rect 200632 300880 200638 300892
rect 269942 300880 269948 300892
rect 200632 300852 269948 300880
rect 200632 300840 200638 300852
rect 269942 300840 269948 300852
rect 270000 300840 270006 300892
rect 64598 300772 64604 300824
rect 64656 300812 64662 300824
rect 66806 300812 66812 300824
rect 64656 300784 66812 300812
rect 64656 300772 64662 300784
rect 66806 300772 66812 300784
rect 66864 300772 66870 300824
rect 162210 300092 162216 300144
rect 162268 300132 162274 300144
rect 225966 300132 225972 300144
rect 162268 300104 225972 300132
rect 162268 300092 162274 300104
rect 225966 300092 225972 300104
rect 226024 300092 226030 300144
rect 184198 299548 184204 299600
rect 184256 299588 184262 299600
rect 253198 299588 253204 299600
rect 184256 299560 253204 299588
rect 184256 299548 184262 299560
rect 253198 299548 253204 299560
rect 253256 299548 253262 299600
rect 58894 299480 58900 299532
rect 58952 299520 58958 299532
rect 66438 299520 66444 299532
rect 58952 299492 66444 299520
rect 58952 299480 58958 299492
rect 66438 299480 66444 299492
rect 66496 299480 66502 299532
rect 227070 299480 227076 299532
rect 227128 299520 227134 299532
rect 228910 299520 228916 299532
rect 227128 299492 228916 299520
rect 227128 299480 227134 299492
rect 228910 299480 228916 299492
rect 228968 299520 228974 299532
rect 303614 299520 303620 299532
rect 228968 299492 303620 299520
rect 228968 299480 228974 299492
rect 303614 299480 303620 299492
rect 303672 299480 303678 299532
rect 157242 299140 157248 299192
rect 157300 299180 157306 299192
rect 164142 299180 164148 299192
rect 157300 299152 164148 299180
rect 157300 299140 157306 299152
rect 164142 299140 164148 299152
rect 164200 299140 164206 299192
rect 155218 298800 155224 298852
rect 155276 298840 155282 298852
rect 173342 298840 173348 298852
rect 155276 298812 173348 298840
rect 155276 298800 155282 298812
rect 173342 298800 173348 298812
rect 173400 298800 173406 298852
rect 165522 298732 165528 298784
rect 165580 298772 165586 298784
rect 246390 298772 246396 298784
rect 165580 298744 246396 298772
rect 165580 298732 165586 298744
rect 246390 298732 246396 298744
rect 246448 298732 246454 298784
rect 200206 298120 200212 298172
rect 200264 298160 200270 298172
rect 202874 298160 202880 298172
rect 200264 298132 202880 298160
rect 200264 298120 200270 298132
rect 202874 298120 202880 298132
rect 202932 298120 202938 298172
rect 209038 298120 209044 298172
rect 209096 298160 209102 298172
rect 209406 298160 209412 298172
rect 209096 298132 209412 298160
rect 209096 298120 209102 298132
rect 209406 298120 209412 298132
rect 209464 298160 209470 298172
rect 265618 298160 265624 298172
rect 209464 298132 265624 298160
rect 209464 298120 209470 298132
rect 265618 298120 265624 298132
rect 265676 298120 265682 298172
rect 246298 297440 246304 297492
rect 246356 297480 246362 297492
rect 254118 297480 254124 297492
rect 246356 297452 254124 297480
rect 246356 297440 246362 297452
rect 254118 297440 254124 297452
rect 254176 297440 254182 297492
rect 202874 297372 202880 297424
rect 202932 297412 202938 297424
rect 295334 297412 295340 297424
rect 202932 297384 295340 297412
rect 202932 297372 202938 297384
rect 295334 297372 295340 297384
rect 295392 297372 295398 297424
rect 164970 297304 164976 297356
rect 165028 297344 165034 297356
rect 165706 297344 165712 297356
rect 165028 297316 165712 297344
rect 165028 297304 165034 297316
rect 165706 297304 165712 297316
rect 165764 297304 165770 297356
rect 64690 296692 64696 296744
rect 64748 296732 64754 296744
rect 66622 296732 66628 296744
rect 64748 296704 66628 296732
rect 64748 296692 64754 296704
rect 66622 296692 66628 296704
rect 66680 296692 66686 296744
rect 191098 296692 191104 296744
rect 191156 296732 191162 296744
rect 245102 296732 245108 296744
rect 191156 296704 245108 296732
rect 191156 296692 191162 296704
rect 245102 296692 245108 296704
rect 245160 296692 245166 296744
rect 53742 296624 53748 296676
rect 53800 296664 53806 296676
rect 66438 296664 66444 296676
rect 53800 296636 66444 296664
rect 53800 296624 53806 296636
rect 66438 296624 66444 296636
rect 66496 296624 66502 296676
rect 155218 296012 155224 296064
rect 155276 296052 155282 296064
rect 175274 296052 175280 296064
rect 155276 296024 175280 296052
rect 155276 296012 155282 296024
rect 175274 296012 175280 296024
rect 175332 296052 175338 296064
rect 240778 296052 240784 296064
rect 175332 296024 240784 296052
rect 175332 296012 175338 296024
rect 240778 296012 240784 296024
rect 240836 296012 240842 296064
rect 156414 295944 156420 295996
rect 156472 295984 156478 295996
rect 244458 295984 244464 295996
rect 156472 295956 244464 295984
rect 156472 295944 156478 295956
rect 244458 295944 244464 295956
rect 244516 295944 244522 295996
rect 245102 295944 245108 295996
rect 245160 295984 245166 295996
rect 259546 295984 259552 295996
rect 245160 295956 259552 295984
rect 245160 295944 245166 295956
rect 259546 295944 259552 295956
rect 259604 295944 259610 295996
rect 156322 295264 156328 295316
rect 156380 295304 156386 295316
rect 172698 295304 172704 295316
rect 156380 295276 172704 295304
rect 156380 295264 156386 295276
rect 172698 295264 172704 295276
rect 172756 295304 172762 295316
rect 173802 295304 173808 295316
rect 172756 295276 173808 295304
rect 172756 295264 172762 295276
rect 173802 295264 173808 295276
rect 173860 295264 173866 295316
rect 173802 294652 173808 294704
rect 173860 294692 173866 294704
rect 197354 294692 197360 294704
rect 173860 294664 197360 294692
rect 173860 294652 173866 294664
rect 197354 294652 197360 294664
rect 197412 294652 197418 294704
rect 193858 294584 193864 294636
rect 193916 294624 193922 294636
rect 245838 294624 245844 294636
rect 193916 294596 245844 294624
rect 193916 294584 193922 294596
rect 245838 294584 245844 294596
rect 245896 294584 245902 294636
rect 61746 294040 61752 294092
rect 61804 294080 61810 294092
rect 66806 294080 66812 294092
rect 61804 294052 66812 294080
rect 61804 294040 61810 294052
rect 66806 294040 66812 294052
rect 66864 294040 66870 294092
rect 15838 293972 15844 294024
rect 15896 294012 15902 294024
rect 67542 294012 67548 294024
rect 15896 293984 67548 294012
rect 15896 293972 15902 293984
rect 67542 293972 67548 293984
rect 67600 293972 67606 294024
rect 200022 293972 200028 294024
rect 200080 294012 200086 294024
rect 222194 294012 222200 294024
rect 200080 293984 222200 294012
rect 200080 293972 200086 293984
rect 222194 293972 222200 293984
rect 222252 293972 222258 294024
rect 227806 293972 227812 294024
rect 227864 294012 227870 294024
rect 228450 294012 228456 294024
rect 227864 293984 228456 294012
rect 227864 293972 227870 293984
rect 228450 293972 228456 293984
rect 228508 294012 228514 294024
rect 278038 294012 278044 294024
rect 228508 293984 278044 294012
rect 228508 293972 228514 293984
rect 278038 293972 278044 293984
rect 278096 293972 278102 294024
rect 59170 293904 59176 293956
rect 59228 293944 59234 293956
rect 66806 293944 66812 293956
rect 59228 293916 66812 293944
rect 59228 293904 59234 293916
rect 66806 293904 66812 293916
rect 66864 293904 66870 293956
rect 238110 293904 238116 293956
rect 238168 293944 238174 293956
rect 240502 293944 240508 293956
rect 238168 293916 240508 293944
rect 238168 293904 238174 293916
rect 240502 293904 240508 293916
rect 240560 293904 240566 293956
rect 204990 293224 204996 293276
rect 205048 293264 205054 293276
rect 235994 293264 236000 293276
rect 205048 293236 236000 293264
rect 205048 293224 205054 293236
rect 235994 293224 236000 293236
rect 236052 293224 236058 293276
rect 2774 292816 2780 292868
rect 2832 292856 2838 292868
rect 4798 292856 4804 292868
rect 2832 292828 4804 292856
rect 2832 292816 2838 292828
rect 4798 292816 4804 292828
rect 4856 292816 4862 292868
rect 156506 292612 156512 292664
rect 156564 292652 156570 292664
rect 166258 292652 166264 292664
rect 156564 292624 166264 292652
rect 156564 292612 156570 292624
rect 166258 292612 166264 292624
rect 166316 292612 166322 292664
rect 157242 292544 157248 292596
rect 157300 292584 157306 292596
rect 220170 292584 220176 292596
rect 157300 292556 220176 292584
rect 157300 292544 157306 292556
rect 220170 292544 220176 292556
rect 220228 292544 220234 292596
rect 231118 292544 231124 292596
rect 231176 292584 231182 292596
rect 233142 292584 233148 292596
rect 231176 292556 233148 292584
rect 231176 292544 231182 292556
rect 233142 292544 233148 292556
rect 233200 292584 233206 292596
rect 583386 292584 583392 292596
rect 233200 292556 583392 292584
rect 233200 292544 233206 292556
rect 583386 292544 583392 292556
rect 583444 292544 583450 292596
rect 14458 292476 14464 292528
rect 14516 292516 14522 292528
rect 60458 292516 60464 292528
rect 14516 292488 60464 292516
rect 14516 292476 14522 292488
rect 60458 292476 60464 292488
rect 60516 292516 60522 292528
rect 66898 292516 66904 292528
rect 60516 292488 66904 292516
rect 60516 292476 60522 292488
rect 66898 292476 66904 292488
rect 66956 292476 66962 292528
rect 197354 291796 197360 291848
rect 197412 291836 197418 291848
rect 209038 291836 209044 291848
rect 197412 291808 209044 291836
rect 197412 291796 197418 291808
rect 209038 291796 209044 291808
rect 209096 291796 209102 291848
rect 222470 291660 222476 291712
rect 222528 291700 222534 291712
rect 223022 291700 223028 291712
rect 222528 291672 223028 291700
rect 222528 291660 222534 291672
rect 223022 291660 223028 291672
rect 223080 291660 223086 291712
rect 223022 291252 223028 291304
rect 223080 291292 223086 291304
rect 253934 291292 253940 291304
rect 223080 291264 253940 291292
rect 223080 291252 223086 291264
rect 253934 291252 253940 291264
rect 253992 291252 253998 291304
rect 156046 291184 156052 291236
rect 156104 291224 156110 291236
rect 193858 291224 193864 291236
rect 156104 291196 193864 291224
rect 156104 291184 156110 291196
rect 193858 291184 193864 291196
rect 193916 291184 193922 291236
rect 204990 291184 204996 291236
rect 205048 291224 205054 291236
rect 218606 291224 218612 291236
rect 205048 291196 218612 291224
rect 205048 291184 205054 291196
rect 218606 291184 218612 291196
rect 218664 291184 218670 291236
rect 236086 291184 236092 291236
rect 236144 291224 236150 291236
rect 236638 291224 236644 291236
rect 236144 291196 236644 291224
rect 236144 291184 236150 291196
rect 236638 291184 236644 291196
rect 236696 291224 236702 291236
rect 306558 291224 306564 291236
rect 236696 291196 306564 291224
rect 236696 291184 236702 291196
rect 306558 291184 306564 291196
rect 306616 291184 306622 291236
rect 63310 289892 63316 289944
rect 63368 289932 63374 289944
rect 66806 289932 66812 289944
rect 63368 289904 66812 289932
rect 63368 289892 63374 289904
rect 66806 289892 66812 289904
rect 66864 289892 66870 289944
rect 199470 289892 199476 289944
rect 199528 289932 199534 289944
rect 256878 289932 256884 289944
rect 199528 289904 256884 289932
rect 199528 289892 199534 289904
rect 256878 289892 256884 289904
rect 256936 289892 256942 289944
rect 157242 289824 157248 289876
rect 157300 289864 157306 289876
rect 247402 289864 247408 289876
rect 157300 289836 247408 289864
rect 157300 289824 157306 289836
rect 247402 289824 247408 289836
rect 247460 289824 247466 289876
rect 238018 289076 238024 289128
rect 238076 289116 238082 289128
rect 242342 289116 242348 289128
rect 238076 289088 242348 289116
rect 238076 289076 238082 289088
rect 242342 289076 242348 289088
rect 242400 289076 242406 289128
rect 157242 288464 157248 288516
rect 157300 288504 157306 288516
rect 224494 288504 224500 288516
rect 157300 288476 224500 288504
rect 157300 288464 157306 288476
rect 224494 288464 224500 288476
rect 224552 288464 224558 288516
rect 242342 288464 242348 288516
rect 242400 288504 242406 288516
rect 280154 288504 280160 288516
rect 242400 288476 280160 288504
rect 242400 288464 242406 288476
rect 280154 288464 280160 288476
rect 280212 288464 280218 288516
rect 171226 288396 171232 288448
rect 171284 288436 171290 288448
rect 244366 288436 244372 288448
rect 171284 288408 244372 288436
rect 171284 288396 171290 288408
rect 244366 288396 244372 288408
rect 244424 288396 244430 288448
rect 180334 287104 180340 287156
rect 180392 287144 180398 287156
rect 223574 287144 223580 287156
rect 180392 287116 223580 287144
rect 180392 287104 180398 287116
rect 223574 287104 223580 287116
rect 223632 287104 223638 287156
rect 230750 287104 230756 287156
rect 230808 287144 230814 287156
rect 230808 287116 231440 287144
rect 230808 287104 230814 287116
rect 52178 287036 52184 287088
rect 52236 287076 52242 287088
rect 66622 287076 66628 287088
rect 52236 287048 66628 287076
rect 52236 287036 52242 287048
rect 66622 287036 66628 287048
rect 66680 287036 66686 287088
rect 157242 287036 157248 287088
rect 157300 287076 157306 287088
rect 231302 287076 231308 287088
rect 157300 287048 231308 287076
rect 157300 287036 157306 287048
rect 231302 287036 231308 287048
rect 231360 287036 231366 287088
rect 231412 287076 231440 287116
rect 233878 287104 233884 287156
rect 233936 287144 233942 287156
rect 244182 287144 244188 287156
rect 233936 287116 244188 287144
rect 233936 287104 233942 287116
rect 244182 287104 244188 287116
rect 244240 287104 244246 287156
rect 255314 287076 255320 287088
rect 231412 287048 255320 287076
rect 255314 287036 255320 287048
rect 255372 287036 255378 287088
rect 224218 286356 224224 286408
rect 224276 286396 224282 286408
rect 229278 286396 229284 286408
rect 224276 286368 229284 286396
rect 224276 286356 224282 286368
rect 229278 286356 229284 286368
rect 229336 286396 229342 286408
rect 230106 286396 230112 286408
rect 229336 286368 230112 286396
rect 229336 286356 229342 286368
rect 230106 286356 230112 286368
rect 230164 286356 230170 286408
rect 163590 286288 163596 286340
rect 163648 286328 163654 286340
rect 191190 286328 191196 286340
rect 163648 286300 191196 286328
rect 163648 286288 163654 286300
rect 191190 286288 191196 286300
rect 191248 286288 191254 286340
rect 210418 286220 210424 286272
rect 210476 286260 210482 286272
rect 211430 286260 211436 286272
rect 210476 286232 211436 286260
rect 210476 286220 210482 286232
rect 211430 286220 211436 286232
rect 211488 286220 211494 286272
rect 220078 285880 220084 285932
rect 220136 285920 220142 285932
rect 220136 285892 229094 285920
rect 220136 285880 220142 285892
rect 198826 285744 198832 285796
rect 198884 285784 198890 285796
rect 205542 285784 205548 285796
rect 198884 285756 205548 285784
rect 198884 285744 198890 285756
rect 205542 285744 205548 285756
rect 205600 285744 205606 285796
rect 55122 285676 55128 285728
rect 55180 285716 55186 285728
rect 66806 285716 66812 285728
rect 55180 285688 66812 285716
rect 55180 285676 55186 285688
rect 66806 285676 66812 285688
rect 66864 285676 66870 285728
rect 199378 285676 199384 285728
rect 199436 285716 199442 285728
rect 204622 285716 204628 285728
rect 199436 285688 204628 285716
rect 199436 285676 199442 285688
rect 204622 285676 204628 285688
rect 204680 285676 204686 285728
rect 204898 285676 204904 285728
rect 204956 285716 204962 285728
rect 208118 285716 208124 285728
rect 204956 285688 208124 285716
rect 204956 285676 204962 285688
rect 208118 285676 208124 285688
rect 208176 285676 208182 285728
rect 211798 285676 211804 285728
rect 211856 285716 211862 285728
rect 213822 285716 213828 285728
rect 211856 285688 213828 285716
rect 211856 285676 211862 285688
rect 213822 285676 213828 285688
rect 213880 285676 213886 285728
rect 220722 285676 220728 285728
rect 220780 285716 220786 285728
rect 222102 285716 222108 285728
rect 220780 285688 222108 285716
rect 220780 285676 220786 285688
rect 222102 285676 222108 285688
rect 222160 285676 222166 285728
rect 229066 285716 229094 285892
rect 237558 285812 237564 285864
rect 237616 285852 237622 285864
rect 238662 285852 238668 285864
rect 237616 285824 238668 285852
rect 237616 285812 237622 285824
rect 238662 285812 238668 285824
rect 238720 285812 238726 285864
rect 230106 285744 230112 285796
rect 230164 285784 230170 285796
rect 246114 285784 246120 285796
rect 230164 285756 246120 285784
rect 230164 285744 230170 285756
rect 246114 285744 246120 285756
rect 246172 285744 246178 285796
rect 269758 285716 269764 285728
rect 229066 285688 269764 285716
rect 269758 285676 269764 285688
rect 269816 285676 269822 285728
rect 200114 285268 200120 285320
rect 200172 285308 200178 285320
rect 200942 285308 200948 285320
rect 200172 285280 200948 285308
rect 200172 285268 200178 285280
rect 200942 285268 200948 285280
rect 201000 285268 201006 285320
rect 222194 285268 222200 285320
rect 222252 285308 222258 285320
rect 222654 285308 222660 285320
rect 222252 285280 222660 285308
rect 222252 285268 222258 285280
rect 222654 285268 222660 285280
rect 222712 285268 222718 285320
rect 57790 284928 57796 284980
rect 57848 284968 57854 284980
rect 65518 284968 65524 284980
rect 57848 284940 65524 284968
rect 57848 284928 57854 284940
rect 65518 284928 65524 284940
rect 65576 284928 65582 284980
rect 159542 284384 159548 284436
rect 159600 284424 159606 284436
rect 216766 284424 216772 284436
rect 159600 284396 216772 284424
rect 159600 284384 159606 284396
rect 216766 284384 216772 284396
rect 216824 284384 216830 284436
rect 230474 284384 230480 284436
rect 230532 284424 230538 284436
rect 231670 284424 231676 284436
rect 230532 284396 231676 284424
rect 230532 284384 230538 284396
rect 231670 284384 231676 284396
rect 231728 284424 231734 284436
rect 281902 284424 281908 284436
rect 231728 284396 281908 284424
rect 231728 284384 231734 284396
rect 281902 284384 281908 284396
rect 281960 284384 281966 284436
rect 156414 284316 156420 284368
rect 156472 284356 156478 284368
rect 243906 284356 243912 284368
rect 156472 284328 243912 284356
rect 156472 284316 156478 284328
rect 243906 284316 243912 284328
rect 243964 284316 243970 284368
rect 191190 283908 191196 283960
rect 191248 283948 191254 283960
rect 201402 283948 201408 283960
rect 191248 283920 201408 283948
rect 191248 283908 191254 283920
rect 201402 283908 201408 283920
rect 201460 283908 201466 283960
rect 244182 283840 244188 283892
rect 244240 283880 244246 283892
rect 282914 283880 282920 283892
rect 244240 283852 282920 283880
rect 244240 283840 244246 283852
rect 282914 283840 282920 283852
rect 282972 283840 282978 283892
rect 162118 283568 162124 283620
rect 162176 283608 162182 283620
rect 188982 283608 188988 283620
rect 162176 283580 188988 283608
rect 162176 283568 162182 283580
rect 188982 283568 188988 283580
rect 189040 283568 189046 283620
rect 157242 283160 157248 283212
rect 157300 283200 157306 283212
rect 162762 283200 162768 283212
rect 157300 283172 162768 283200
rect 157300 283160 157306 283172
rect 162762 283160 162768 283172
rect 162820 283160 162826 283212
rect 246298 283160 246304 283212
rect 246356 283200 246362 283212
rect 247034 283200 247040 283212
rect 246356 283172 247040 283200
rect 246356 283160 246362 283172
rect 247034 283160 247040 283172
rect 247092 283200 247098 283212
rect 250070 283200 250076 283212
rect 247092 283172 250076 283200
rect 247092 283160 247098 283172
rect 250070 283160 250076 283172
rect 250128 283160 250134 283212
rect 245930 282820 245936 282872
rect 245988 282860 245994 282872
rect 254118 282860 254124 282872
rect 245988 282832 254124 282860
rect 245988 282820 245994 282832
rect 254118 282820 254124 282832
rect 254176 282860 254182 282872
rect 582742 282860 582748 282872
rect 254176 282832 582748 282860
rect 254176 282820 254182 282832
rect 582742 282820 582748 282832
rect 582800 282820 582806 282872
rect 162762 282140 162768 282192
rect 162820 282180 162826 282192
rect 184842 282180 184848 282192
rect 162820 282152 184848 282180
rect 162820 282140 162826 282152
rect 184842 282140 184848 282152
rect 184900 282140 184906 282192
rect 185026 282140 185032 282192
rect 185084 282180 185090 282192
rect 197078 282180 197084 282192
rect 185084 282152 197084 282180
rect 185084 282140 185090 282152
rect 197078 282140 197084 282152
rect 197136 282140 197142 282192
rect 60550 281528 60556 281580
rect 60608 281568 60614 281580
rect 66806 281568 66812 281580
rect 60608 281540 66812 281568
rect 60608 281528 60614 281540
rect 66806 281528 66812 281540
rect 66864 281528 66870 281580
rect 184842 281528 184848 281580
rect 184900 281568 184906 281580
rect 197354 281568 197360 281580
rect 184900 281540 197360 281568
rect 184900 281528 184906 281540
rect 197354 281528 197360 281540
rect 197412 281528 197418 281580
rect 157242 281460 157248 281512
rect 157300 281500 157306 281512
rect 184198 281500 184204 281512
rect 157300 281472 184204 281500
rect 157300 281460 157306 281472
rect 184198 281460 184204 281472
rect 184256 281460 184262 281512
rect 181622 281392 181628 281444
rect 181680 281432 181686 281444
rect 197354 281432 197360 281444
rect 181680 281404 197360 281432
rect 181680 281392 181686 281404
rect 197354 281392 197360 281404
rect 197412 281392 197418 281444
rect 156874 280780 156880 280832
rect 156932 280820 156938 280832
rect 171226 280820 171232 280832
rect 156932 280792 171232 280820
rect 156932 280780 156938 280792
rect 171226 280780 171232 280792
rect 171284 280780 171290 280832
rect 245930 280780 245936 280832
rect 245988 280820 245994 280832
rect 248598 280820 248604 280832
rect 245988 280792 248604 280820
rect 245988 280780 245994 280792
rect 248598 280780 248604 280792
rect 248656 280820 248662 280832
rect 311986 280820 311992 280832
rect 248656 280792 311992 280820
rect 248656 280780 248662 280792
rect 311986 280780 311992 280792
rect 312044 280780 312050 280832
rect 63218 280168 63224 280220
rect 63276 280208 63282 280220
rect 66806 280208 66812 280220
rect 63276 280180 66812 280208
rect 63276 280168 63282 280180
rect 66806 280168 66812 280180
rect 66864 280168 66870 280220
rect 245470 280168 245476 280220
rect 245528 280208 245534 280220
rect 273990 280208 273996 280220
rect 245528 280180 273996 280208
rect 245528 280168 245534 280180
rect 273990 280168 273996 280180
rect 274048 280168 274054 280220
rect 195422 279692 195428 279744
rect 195480 279732 195486 279744
rect 198734 279732 198740 279744
rect 195480 279704 198740 279732
rect 195480 279692 195486 279704
rect 198734 279692 198740 279704
rect 198792 279692 198798 279744
rect 158162 279624 158168 279676
rect 158220 279664 158226 279676
rect 162210 279664 162216 279676
rect 158220 279636 162216 279664
rect 158220 279624 158226 279636
rect 162210 279624 162216 279636
rect 162268 279624 162274 279676
rect 157242 279488 157248 279540
rect 157300 279528 157306 279540
rect 158714 279528 158720 279540
rect 157300 279500 158720 279528
rect 157300 279488 157306 279500
rect 158714 279488 158720 279500
rect 158772 279528 158778 279540
rect 158772 279500 161474 279528
rect 158772 279488 158778 279500
rect 161446 279460 161474 279500
rect 171870 279460 171876 279472
rect 161446 279432 171876 279460
rect 171870 279420 171876 279432
rect 171928 279420 171934 279472
rect 245930 279420 245936 279472
rect 245988 279460 245994 279472
rect 251266 279460 251272 279472
rect 245988 279432 251272 279460
rect 245988 279420 245994 279432
rect 251266 279420 251272 279432
rect 251324 279420 251330 279472
rect 245654 278944 245660 278996
rect 245712 278984 245718 278996
rect 247310 278984 247316 278996
rect 245712 278956 247316 278984
rect 245712 278944 245718 278956
rect 247310 278944 247316 278956
rect 247368 278944 247374 278996
rect 192570 278808 192576 278860
rect 192628 278848 192634 278860
rect 197354 278848 197360 278860
rect 192628 278820 197360 278848
rect 192628 278808 192634 278820
rect 197354 278808 197360 278820
rect 197412 278808 197418 278860
rect 11698 278740 11704 278792
rect 11756 278780 11762 278792
rect 59078 278780 59084 278792
rect 11756 278752 59084 278780
rect 11756 278740 11762 278752
rect 59078 278740 59084 278752
rect 59136 278780 59142 278792
rect 67174 278780 67180 278792
rect 59136 278752 67180 278780
rect 59136 278740 59142 278752
rect 67174 278740 67180 278752
rect 67232 278740 67238 278792
rect 251266 278740 251272 278792
rect 251324 278780 251330 278792
rect 583202 278780 583208 278792
rect 251324 278752 583208 278780
rect 251324 278740 251330 278752
rect 583202 278740 583208 278752
rect 583260 278740 583266 278792
rect 191650 278672 191656 278724
rect 191708 278712 191714 278724
rect 197354 278712 197360 278724
rect 191708 278684 197360 278712
rect 191708 278672 191714 278684
rect 197354 278672 197360 278684
rect 197412 278672 197418 278724
rect 157058 278060 157064 278112
rect 157116 278100 157122 278112
rect 170582 278100 170588 278112
rect 157116 278072 170588 278100
rect 157116 278060 157122 278072
rect 170582 278060 170588 278072
rect 170640 278060 170646 278112
rect 180242 278060 180248 278112
rect 180300 278100 180306 278112
rect 198826 278100 198832 278112
rect 180300 278072 198832 278100
rect 180300 278060 180306 278072
rect 198826 278060 198832 278072
rect 198884 278060 198890 278112
rect 245930 278060 245936 278112
rect 245988 278100 245994 278112
rect 249794 278100 249800 278112
rect 245988 278072 249800 278100
rect 245988 278060 245994 278072
rect 249794 278060 249800 278072
rect 249852 278060 249858 278112
rect 158162 277992 158168 278044
rect 158220 278032 158226 278044
rect 185026 278032 185032 278044
rect 158220 278004 185032 278032
rect 158220 277992 158226 278004
rect 185026 277992 185032 278004
rect 185084 277992 185090 278044
rect 246022 277992 246028 278044
rect 246080 278032 246086 278044
rect 249978 278032 249984 278044
rect 246080 278004 249984 278032
rect 246080 277992 246086 278004
rect 249978 277992 249984 278004
rect 250036 278032 250042 278044
rect 583294 278032 583300 278044
rect 250036 278004 583300 278032
rect 250036 277992 250042 278004
rect 583294 277992 583300 278004
rect 583352 277992 583358 278044
rect 57698 277380 57704 277432
rect 57756 277420 57762 277432
rect 66438 277420 66444 277432
rect 57756 277392 66444 277420
rect 57756 277380 57762 277392
rect 66438 277380 66444 277392
rect 66496 277380 66502 277432
rect 157334 276700 157340 276752
rect 157392 276740 157398 276752
rect 197354 276740 197360 276752
rect 157392 276712 197360 276740
rect 157392 276700 157398 276712
rect 197354 276700 197360 276712
rect 197412 276700 197418 276752
rect 199378 276672 199384 276684
rect 155328 276644 199384 276672
rect 155328 276616 155356 276644
rect 199378 276632 199384 276644
rect 199436 276632 199442 276684
rect 245746 276632 245752 276684
rect 245804 276672 245810 276684
rect 278130 276672 278136 276684
rect 245804 276644 278136 276672
rect 245804 276632 245810 276644
rect 278130 276632 278136 276644
rect 278188 276632 278194 276684
rect 155310 276564 155316 276616
rect 155368 276564 155374 276616
rect 53466 276020 53472 276072
rect 53524 276060 53530 276072
rect 66806 276060 66812 276072
rect 53524 276032 66812 276060
rect 53524 276020 53530 276032
rect 66806 276020 66812 276032
rect 66864 276020 66870 276072
rect 245930 275952 245936 276004
rect 245988 275992 245994 276004
rect 254026 275992 254032 276004
rect 245988 275964 254032 275992
rect 245988 275952 245994 275964
rect 254026 275952 254032 275964
rect 254084 275992 254090 276004
rect 582650 275992 582656 276004
rect 254084 275964 582656 275992
rect 254084 275952 254090 275964
rect 582650 275952 582656 275964
rect 582708 275952 582714 276004
rect 157242 275272 157248 275324
rect 157300 275312 157306 275324
rect 173250 275312 173256 275324
rect 157300 275284 173256 275312
rect 157300 275272 157306 275284
rect 173250 275272 173256 275284
rect 173308 275272 173314 275324
rect 160922 274728 160928 274780
rect 160980 274768 160986 274780
rect 197354 274768 197360 274780
rect 160980 274740 197360 274768
rect 160980 274728 160986 274740
rect 197354 274728 197360 274740
rect 197412 274728 197418 274780
rect 56410 274660 56416 274712
rect 56468 274700 56474 274712
rect 66806 274700 66812 274712
rect 56468 274672 66812 274700
rect 56468 274660 56474 274672
rect 66806 274660 66812 274672
rect 66864 274660 66870 274712
rect 157242 274660 157248 274712
rect 157300 274700 157306 274712
rect 161014 274700 161020 274712
rect 157300 274672 161020 274700
rect 157300 274660 157306 274672
rect 161014 274660 161020 274672
rect 161072 274660 161078 274712
rect 156506 274592 156512 274644
rect 156564 274632 156570 274644
rect 191098 274632 191104 274644
rect 156564 274604 191104 274632
rect 156564 274592 156570 274604
rect 191098 274592 191104 274604
rect 191156 274592 191162 274644
rect 196710 274524 196716 274576
rect 196768 274564 196774 274576
rect 200022 274564 200028 274576
rect 196768 274536 200028 274564
rect 196768 274524 196774 274536
rect 200022 274524 200028 274536
rect 200080 274524 200086 274576
rect 182910 273912 182916 273964
rect 182968 273952 182974 273964
rect 195514 273952 195520 273964
rect 182968 273924 195520 273952
rect 182968 273912 182974 273924
rect 195514 273912 195520 273924
rect 195572 273912 195578 273964
rect 62022 273232 62028 273284
rect 62080 273272 62086 273284
rect 66806 273272 66812 273284
rect 62080 273244 66812 273272
rect 62080 273232 62086 273244
rect 66806 273232 66812 273244
rect 66864 273232 66870 273284
rect 245654 273232 245660 273284
rect 245712 273272 245718 273284
rect 254026 273272 254032 273284
rect 245712 273244 254032 273272
rect 245712 273232 245718 273244
rect 254026 273232 254032 273244
rect 254084 273232 254090 273284
rect 176562 273164 176568 273216
rect 176620 273204 176626 273216
rect 197354 273204 197360 273216
rect 176620 273176 197360 273204
rect 176620 273164 176626 273176
rect 197354 273164 197360 273176
rect 197412 273164 197418 273216
rect 185578 273096 185584 273148
rect 185636 273136 185642 273148
rect 197446 273136 197452 273148
rect 185636 273108 197452 273136
rect 185636 273096 185642 273108
rect 197446 273096 197452 273108
rect 197504 273096 197510 273148
rect 260098 272484 260104 272536
rect 260156 272524 260162 272536
rect 302234 272524 302240 272536
rect 260156 272496 302240 272524
rect 260156 272484 260162 272496
rect 302234 272484 302240 272496
rect 302292 272484 302298 272536
rect 63126 271872 63132 271924
rect 63184 271912 63190 271924
rect 66806 271912 66812 271924
rect 63184 271884 66812 271912
rect 63184 271872 63190 271884
rect 66806 271872 66812 271884
rect 66864 271872 66870 271924
rect 245838 271872 245844 271924
rect 245896 271912 245902 271924
rect 251266 271912 251272 271924
rect 245896 271884 251272 271912
rect 245896 271872 245902 271884
rect 251266 271872 251272 271884
rect 251324 271912 251330 271924
rect 259454 271912 259460 271924
rect 251324 271884 259460 271912
rect 251324 271872 251330 271884
rect 259454 271872 259460 271884
rect 259512 271872 259518 271924
rect 156966 271124 156972 271176
rect 157024 271164 157030 271176
rect 191374 271164 191380 271176
rect 157024 271136 191380 271164
rect 157024 271124 157030 271136
rect 191374 271124 191380 271136
rect 191432 271124 191438 271176
rect 48222 270512 48228 270564
rect 48280 270552 48286 270564
rect 66806 270552 66812 270564
rect 48280 270524 66812 270552
rect 48280 270512 48286 270524
rect 66806 270512 66812 270524
rect 66864 270512 66870 270564
rect 166442 270512 166448 270564
rect 166500 270552 166506 270564
rect 197446 270552 197452 270564
rect 166500 270524 197452 270552
rect 166500 270512 166506 270524
rect 197446 270512 197452 270524
rect 197504 270512 197510 270564
rect 245838 270512 245844 270564
rect 245896 270552 245902 270564
rect 252830 270552 252836 270564
rect 245896 270524 252836 270552
rect 245896 270512 245902 270524
rect 252830 270512 252836 270524
rect 252888 270512 252894 270564
rect 164234 270444 164240 270496
rect 164292 270484 164298 270496
rect 197354 270484 197360 270496
rect 164292 270456 197360 270484
rect 164292 270444 164298 270456
rect 197354 270444 197360 270456
rect 197412 270444 197418 270496
rect 256786 270444 256792 270496
rect 256844 270484 256850 270496
rect 583018 270484 583024 270496
rect 256844 270456 583024 270484
rect 256844 270444 256850 270456
rect 583018 270444 583024 270456
rect 583076 270444 583082 270496
rect 163682 270240 163688 270292
rect 163740 270280 163746 270292
rect 164234 270280 164240 270292
rect 163740 270252 164240 270280
rect 163740 270240 163746 270252
rect 164234 270240 164240 270252
rect 164292 270240 164298 270292
rect 246298 269832 246304 269884
rect 246356 269872 246362 269884
rect 247034 269872 247040 269884
rect 246356 269844 247040 269872
rect 246356 269832 246362 269844
rect 247034 269832 247040 269844
rect 247092 269872 247098 269884
rect 252646 269872 252652 269884
rect 247092 269844 252652 269872
rect 247092 269832 247098 269844
rect 252646 269832 252652 269844
rect 252704 269832 252710 269884
rect 4062 269764 4068 269816
rect 4120 269804 4126 269816
rect 21450 269804 21456 269816
rect 4120 269776 21456 269804
rect 4120 269764 4126 269776
rect 21450 269764 21456 269776
rect 21508 269764 21514 269816
rect 245838 269764 245844 269816
rect 245896 269804 245902 269816
rect 256786 269804 256792 269816
rect 245896 269776 256792 269804
rect 245896 269764 245902 269776
rect 256786 269764 256792 269776
rect 256844 269764 256850 269816
rect 181622 269560 181628 269612
rect 181680 269600 181686 269612
rect 186314 269600 186320 269612
rect 181680 269572 186320 269600
rect 181680 269560 181686 269572
rect 186314 269560 186320 269572
rect 186372 269560 186378 269612
rect 64506 269084 64512 269136
rect 64564 269124 64570 269136
rect 66806 269124 66812 269136
rect 64564 269096 66812 269124
rect 64564 269084 64570 269096
rect 66806 269084 66812 269096
rect 66864 269084 66870 269136
rect 157242 269084 157248 269136
rect 157300 269124 157306 269136
rect 178954 269124 178960 269136
rect 157300 269096 178960 269124
rect 157300 269084 157306 269096
rect 178954 269084 178960 269096
rect 179012 269084 179018 269136
rect 21082 269016 21088 269068
rect 21140 269056 21146 269068
rect 22738 269056 22744 269068
rect 21140 269028 22744 269056
rect 21140 269016 21146 269028
rect 22738 269016 22744 269028
rect 22796 269016 22802 269068
rect 67358 269016 67364 269068
rect 67416 269056 67422 269068
rect 67634 269056 67640 269068
rect 67416 269028 67640 269056
rect 67416 269016 67422 269028
rect 67634 269016 67640 269028
rect 67692 269016 67698 269068
rect 156414 269016 156420 269068
rect 156472 269056 156478 269068
rect 180334 269056 180340 269068
rect 156472 269028 180340 269056
rect 156472 269016 156478 269028
rect 180334 269016 180340 269028
rect 180392 269016 180398 269068
rect 245746 269016 245752 269068
rect 245804 269056 245810 269068
rect 255406 269056 255412 269068
rect 245804 269028 255412 269056
rect 245804 269016 245810 269028
rect 255406 269016 255412 269028
rect 255464 269016 255470 269068
rect 178770 268948 178776 269000
rect 178828 268988 178834 269000
rect 197354 268988 197360 269000
rect 178828 268960 197360 268988
rect 178828 268948 178834 268960
rect 197354 268948 197360 268960
rect 197412 268948 197418 269000
rect 55030 268336 55036 268388
rect 55088 268376 55094 268388
rect 66990 268376 66996 268388
rect 55088 268348 66996 268376
rect 55088 268336 55094 268348
rect 66990 268336 66996 268348
rect 67048 268336 67054 268388
rect 180058 268336 180064 268388
rect 180116 268376 180122 268388
rect 197354 268376 197360 268388
rect 180116 268348 197360 268376
rect 180116 268336 180122 268348
rect 197354 268336 197360 268348
rect 197412 268336 197418 268388
rect 255406 268336 255412 268388
rect 255464 268376 255470 268388
rect 582650 268376 582656 268388
rect 255464 268348 582656 268376
rect 255464 268336 255470 268348
rect 582650 268336 582656 268348
rect 582708 268336 582714 268388
rect 195238 267112 195244 267164
rect 195296 267152 195302 267164
rect 197446 267152 197452 267164
rect 195296 267124 197452 267152
rect 195296 267112 195302 267124
rect 197446 267112 197452 267124
rect 197504 267112 197510 267164
rect 3418 266976 3424 267028
rect 3476 267016 3482 267028
rect 21358 267016 21364 267028
rect 3476 266988 21364 267016
rect 3476 266976 3482 266988
rect 21358 266976 21364 266988
rect 21416 266976 21422 267028
rect 245838 266976 245844 267028
rect 245896 267016 245902 267028
rect 288526 267016 288532 267028
rect 245896 266988 288532 267016
rect 245896 266976 245902 266988
rect 288526 266976 288532 266988
rect 288584 266976 288590 267028
rect 64782 266500 64788 266552
rect 64840 266540 64846 266552
rect 66162 266540 66168 266552
rect 64840 266512 66168 266540
rect 64840 266500 64846 266512
rect 66162 266500 66168 266512
rect 66220 266540 66226 266552
rect 66622 266540 66628 266552
rect 66220 266512 66628 266540
rect 66220 266500 66226 266512
rect 66622 266500 66628 266512
rect 66680 266500 66686 266552
rect 173526 266432 173532 266484
rect 173584 266472 173590 266484
rect 197354 266472 197360 266484
rect 173584 266444 197360 266472
rect 173584 266432 173590 266444
rect 197354 266432 197360 266444
rect 197412 266432 197418 266484
rect 157242 266364 157248 266416
rect 157300 266404 157306 266416
rect 184198 266404 184204 266416
rect 157300 266376 184204 266404
rect 157300 266364 157306 266376
rect 184198 266364 184204 266376
rect 184256 266364 184262 266416
rect 245930 266364 245936 266416
rect 245988 266404 245994 266416
rect 263594 266404 263600 266416
rect 245988 266376 263600 266404
rect 245988 266364 245994 266376
rect 263594 266364 263600 266376
rect 263652 266364 263658 266416
rect 245930 265616 245936 265668
rect 245988 265656 245994 265668
rect 251358 265656 251364 265668
rect 245988 265628 251364 265656
rect 245988 265616 245994 265628
rect 251358 265616 251364 265628
rect 251416 265616 251422 265668
rect 263686 265616 263692 265668
rect 263744 265656 263750 265668
rect 583018 265656 583024 265668
rect 263744 265628 583024 265656
rect 263744 265616 263750 265628
rect 583018 265616 583024 265628
rect 583076 265616 583082 265668
rect 41138 264936 41144 264988
rect 41196 264976 41202 264988
rect 66806 264976 66812 264988
rect 41196 264948 66812 264976
rect 41196 264936 41202 264948
rect 66806 264936 66812 264948
rect 66864 264936 66870 264988
rect 157242 264936 157248 264988
rect 157300 264976 157306 264988
rect 171962 264976 171968 264988
rect 157300 264948 171968 264976
rect 157300 264936 157306 264948
rect 171962 264936 171968 264948
rect 172020 264936 172026 264988
rect 186130 264936 186136 264988
rect 186188 264976 186194 264988
rect 197354 264976 197360 264988
rect 186188 264948 197360 264976
rect 186188 264936 186194 264948
rect 197354 264936 197360 264948
rect 197412 264936 197418 264988
rect 188338 264868 188344 264920
rect 188396 264908 188402 264920
rect 197446 264908 197452 264920
rect 188396 264880 197452 264908
rect 188396 264868 188402 264880
rect 197446 264868 197452 264880
rect 197504 264868 197510 264920
rect 41322 264188 41328 264240
rect 41380 264228 41386 264240
rect 58986 264228 58992 264240
rect 41380 264200 58992 264228
rect 41380 264188 41386 264200
rect 58986 264188 58992 264200
rect 59044 264228 59050 264240
rect 66806 264228 66812 264240
rect 59044 264200 66812 264228
rect 59044 264188 59050 264200
rect 66806 264188 66812 264200
rect 66864 264188 66870 264240
rect 166350 264188 166356 264240
rect 166408 264228 166414 264240
rect 187234 264228 187240 264240
rect 166408 264200 187240 264228
rect 166408 264188 166414 264200
rect 187234 264188 187240 264200
rect 187292 264188 187298 264240
rect 246482 264188 246488 264240
rect 246540 264228 246546 264240
rect 299658 264228 299664 264240
rect 246540 264200 299664 264228
rect 246540 264188 246546 264200
rect 299658 264188 299664 264200
rect 299716 264188 299722 264240
rect 245838 263984 245844 264036
rect 245896 264024 245902 264036
rect 248414 264024 248420 264036
rect 245896 263996 248420 264024
rect 245896 263984 245902 263996
rect 248414 263984 248420 263996
rect 248472 263984 248478 264036
rect 60458 263576 60464 263628
rect 60516 263616 60522 263628
rect 66714 263616 66720 263628
rect 60516 263588 66720 263616
rect 60516 263576 60522 263588
rect 66714 263576 66720 263588
rect 66772 263576 66778 263628
rect 195238 263576 195244 263628
rect 195296 263616 195302 263628
rect 197354 263616 197360 263628
rect 195296 263588 197360 263616
rect 195296 263576 195302 263588
rect 197354 263576 197360 263588
rect 197412 263576 197418 263628
rect 52362 262828 52368 262880
rect 52420 262868 52426 262880
rect 66806 262868 66812 262880
rect 52420 262840 66812 262868
rect 52420 262828 52426 262840
rect 66806 262828 66812 262840
rect 66864 262828 66870 262880
rect 251358 262828 251364 262880
rect 251416 262868 251422 262880
rect 259454 262868 259460 262880
rect 251416 262840 259460 262868
rect 251416 262828 251422 262840
rect 259454 262828 259460 262840
rect 259512 262828 259518 262880
rect 156414 262284 156420 262336
rect 156472 262324 156478 262336
rect 170398 262324 170404 262336
rect 156472 262296 170404 262324
rect 156472 262284 156478 262296
rect 170398 262284 170404 262296
rect 170456 262284 170462 262336
rect 159634 262216 159640 262268
rect 159692 262256 159698 262268
rect 195238 262256 195244 262268
rect 159692 262228 195244 262256
rect 159692 262216 159698 262228
rect 195238 262216 195244 262228
rect 195296 262216 195302 262268
rect 164234 262148 164240 262200
rect 164292 262188 164298 262200
rect 169754 262188 169760 262200
rect 164292 262160 169760 262188
rect 164292 262148 164298 262160
rect 169754 262148 169760 262160
rect 169812 262148 169818 262200
rect 161014 261536 161020 261588
rect 161072 261576 161078 261588
rect 177574 261576 177580 261588
rect 161072 261548 177580 261576
rect 161072 261536 161078 261548
rect 177574 261536 177580 261548
rect 177632 261536 177638 261588
rect 186958 261536 186964 261588
rect 187016 261576 187022 261588
rect 197354 261576 197360 261588
rect 187016 261548 197360 261576
rect 187016 261536 187022 261548
rect 197354 261536 197360 261548
rect 197412 261536 197418 261588
rect 246390 261536 246396 261588
rect 246448 261576 246454 261588
rect 247402 261576 247408 261588
rect 246448 261548 247408 261576
rect 246448 261536 246454 261548
rect 247402 261536 247408 261548
rect 247460 261576 247466 261588
rect 248414 261576 248420 261588
rect 247460 261548 248420 261576
rect 247460 261536 247466 261548
rect 248414 261536 248420 261548
rect 248472 261536 248478 261588
rect 21450 261468 21456 261520
rect 21508 261508 21514 261520
rect 63494 261508 63500 261520
rect 21508 261480 63500 261508
rect 21508 261468 21514 261480
rect 63494 261468 63500 261480
rect 63552 261468 63558 261520
rect 173342 261468 173348 261520
rect 173400 261508 173406 261520
rect 199470 261508 199476 261520
rect 173400 261480 199476 261508
rect 173400 261468 173406 261480
rect 199470 261468 199476 261480
rect 199528 261468 199534 261520
rect 265710 261468 265716 261520
rect 265768 261508 265774 261520
rect 580350 261508 580356 261520
rect 265768 261480 580356 261508
rect 265768 261468 265774 261480
rect 580350 261468 580356 261480
rect 580408 261468 580414 261520
rect 63494 260924 63500 260976
rect 63552 260964 63558 260976
rect 64782 260964 64788 260976
rect 63552 260936 64788 260964
rect 63552 260924 63558 260936
rect 64782 260924 64788 260936
rect 64840 260964 64846 260976
rect 66806 260964 66812 260976
rect 64840 260936 66812 260964
rect 64840 260924 64846 260936
rect 66806 260924 66812 260936
rect 66864 260924 66870 260976
rect 157242 260856 157248 260908
rect 157300 260896 157306 260908
rect 164234 260896 164240 260908
rect 157300 260868 164240 260896
rect 157300 260856 157306 260868
rect 164234 260856 164240 260868
rect 164292 260856 164298 260908
rect 156966 260788 156972 260840
rect 157024 260828 157030 260840
rect 177482 260828 177488 260840
rect 157024 260800 177488 260828
rect 157024 260788 157030 260800
rect 177482 260788 177488 260800
rect 177540 260788 177546 260840
rect 245746 260720 245752 260772
rect 245804 260760 245810 260772
rect 251450 260760 251456 260772
rect 245804 260732 251456 260760
rect 245804 260720 245810 260732
rect 251450 260720 251456 260732
rect 251508 260720 251514 260772
rect 156322 260108 156328 260160
rect 156380 260148 156386 260160
rect 179046 260148 179052 260160
rect 156380 260120 179052 260148
rect 156380 260108 156386 260120
rect 179046 260108 179052 260120
rect 179104 260108 179110 260160
rect 253198 259496 253204 259548
rect 253256 259536 253262 259548
rect 276658 259536 276664 259548
rect 253256 259508 276664 259536
rect 253256 259496 253262 259508
rect 276658 259496 276664 259508
rect 276716 259496 276722 259548
rect 178954 259428 178960 259480
rect 179012 259468 179018 259480
rect 182174 259468 182180 259480
rect 179012 259440 182180 259468
rect 179012 259428 179018 259440
rect 182174 259428 182180 259440
rect 182232 259428 182238 259480
rect 193950 259428 193956 259480
rect 194008 259468 194014 259480
rect 197354 259468 197360 259480
rect 194008 259440 197360 259468
rect 194008 259428 194014 259440
rect 197354 259428 197360 259440
rect 197412 259428 197418 259480
rect 244458 259428 244464 259480
rect 244516 259468 244522 259480
rect 291194 259468 291200 259480
rect 244516 259440 291200 259468
rect 244516 259428 244522 259440
rect 291194 259428 291200 259440
rect 291252 259428 291258 259480
rect 169110 259360 169116 259412
rect 169168 259400 169174 259412
rect 197446 259400 197452 259412
rect 169168 259372 197452 259400
rect 169168 259360 169174 259372
rect 197446 259360 197452 259372
rect 197504 259360 197510 259412
rect 245930 259360 245936 259412
rect 245988 259400 245994 259412
rect 253198 259400 253204 259412
rect 245988 259372 253204 259400
rect 245988 259360 245994 259372
rect 253198 259360 253204 259372
rect 253256 259360 253262 259412
rect 264238 259360 264244 259412
rect 264296 259400 264302 259412
rect 579798 259400 579804 259412
rect 264296 259372 579804 259400
rect 264296 259360 264302 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 184290 259292 184296 259344
rect 184348 259332 184354 259344
rect 184750 259332 184756 259344
rect 184348 259304 184756 259332
rect 184348 259292 184354 259304
rect 184750 259292 184756 259304
rect 184808 259292 184814 259344
rect 184750 258680 184756 258732
rect 184808 258720 184814 258732
rect 197354 258720 197360 258732
rect 184808 258692 197360 258720
rect 184808 258680 184814 258692
rect 197354 258680 197360 258692
rect 197412 258680 197418 258732
rect 53742 258068 53748 258120
rect 53800 258108 53806 258120
rect 66254 258108 66260 258120
rect 53800 258080 66260 258108
rect 53800 258068 53806 258080
rect 66254 258068 66260 258080
rect 66312 258068 66318 258120
rect 245838 258068 245844 258120
rect 245896 258108 245902 258120
rect 279418 258108 279424 258120
rect 245896 258080 279424 258108
rect 245896 258068 245902 258080
rect 279418 258068 279424 258080
rect 279476 258068 279482 258120
rect 245654 258000 245660 258052
rect 245712 258040 245718 258052
rect 255590 258040 255596 258052
rect 245712 258012 255596 258040
rect 245712 258000 245718 258012
rect 255590 258000 255596 258012
rect 255648 258000 255654 258052
rect 156874 257932 156880 257984
rect 156932 257972 156938 257984
rect 159542 257972 159548 257984
rect 156932 257944 159548 257972
rect 156932 257932 156938 257944
rect 159542 257932 159548 257944
rect 159600 257932 159606 257984
rect 157242 257320 157248 257372
rect 157300 257360 157306 257372
rect 192570 257360 192576 257372
rect 157300 257332 192576 257360
rect 157300 257320 157306 257332
rect 192570 257320 192576 257332
rect 192628 257320 192634 257372
rect 255590 257320 255596 257372
rect 255648 257360 255654 257372
rect 271230 257360 271236 257372
rect 255648 257332 271236 257360
rect 255648 257320 255654 257332
rect 271230 257320 271236 257332
rect 271288 257320 271294 257372
rect 162762 256708 162768 256760
rect 162820 256748 162826 256760
rect 177942 256748 177948 256760
rect 162820 256720 177948 256748
rect 162820 256708 162826 256720
rect 177942 256708 177948 256720
rect 178000 256748 178006 256760
rect 197446 256748 197452 256760
rect 178000 256720 197452 256748
rect 178000 256708 178006 256720
rect 197446 256708 197452 256720
rect 197504 256708 197510 256760
rect 189810 256640 189816 256692
rect 189868 256680 189874 256692
rect 197354 256680 197360 256692
rect 189868 256652 197360 256680
rect 189868 256640 189874 256652
rect 197354 256640 197360 256652
rect 197412 256640 197418 256692
rect 245930 256572 245936 256624
rect 245988 256612 245994 256624
rect 259546 256612 259552 256624
rect 245988 256584 259552 256612
rect 245988 256572 245994 256584
rect 259546 256572 259552 256584
rect 259604 256612 259610 256624
rect 260742 256612 260748 256624
rect 259604 256584 260748 256612
rect 259604 256572 259610 256584
rect 260742 256572 260748 256584
rect 260800 256572 260806 256624
rect 178678 256164 178684 256216
rect 178736 256204 178742 256216
rect 182910 256204 182916 256216
rect 178736 256176 182916 256204
rect 178736 256164 178742 256176
rect 182910 256164 182916 256176
rect 182968 256164 182974 256216
rect 155218 255960 155224 256012
rect 155276 256000 155282 256012
rect 186958 256000 186964 256012
rect 155276 255972 186964 256000
rect 155276 255960 155282 255972
rect 186958 255960 186964 255972
rect 187016 255960 187022 256012
rect 260742 255960 260748 256012
rect 260800 256000 260806 256012
rect 296714 256000 296720 256012
rect 260800 255972 296720 256000
rect 260800 255960 260806 255972
rect 296714 255960 296720 255972
rect 296772 255960 296778 256012
rect 64598 255280 64604 255332
rect 64656 255320 64662 255332
rect 66806 255320 66812 255332
rect 64656 255292 66812 255320
rect 64656 255280 64662 255292
rect 66806 255280 66812 255292
rect 66864 255280 66870 255332
rect 191098 255280 191104 255332
rect 191156 255320 191162 255332
rect 195422 255320 195428 255332
rect 191156 255292 195428 255320
rect 191156 255280 191162 255292
rect 195422 255280 195428 255292
rect 195480 255280 195486 255332
rect 3418 255212 3424 255264
rect 3476 255252 3482 255264
rect 18598 255252 18604 255264
rect 3476 255224 18604 255252
rect 3476 255212 3482 255224
rect 18598 255212 18604 255224
rect 18656 255212 18662 255264
rect 245838 255212 245844 255264
rect 245896 255252 245902 255264
rect 255498 255252 255504 255264
rect 245896 255224 255504 255252
rect 245896 255212 245902 255224
rect 255498 255212 255504 255224
rect 255556 255212 255562 255264
rect 245930 255144 245936 255196
rect 245988 255184 245994 255196
rect 249794 255184 249800 255196
rect 245988 255156 249800 255184
rect 245988 255144 245994 255156
rect 249794 255144 249800 255156
rect 249852 255144 249858 255196
rect 157242 254600 157248 254652
rect 157300 254640 157306 254652
rect 161658 254640 161664 254652
rect 157300 254612 161664 254640
rect 157300 254600 157306 254612
rect 161658 254600 161664 254612
rect 161716 254640 161722 254652
rect 162670 254640 162676 254652
rect 161716 254612 162676 254640
rect 161716 254600 161722 254612
rect 162670 254600 162676 254612
rect 162728 254600 162734 254652
rect 156506 254532 156512 254584
rect 156564 254572 156570 254584
rect 173802 254572 173808 254584
rect 156564 254544 173808 254572
rect 156564 254532 156570 254544
rect 173802 254532 173808 254544
rect 173860 254532 173866 254584
rect 187694 254532 187700 254584
rect 187752 254572 187758 254584
rect 188798 254572 188804 254584
rect 187752 254544 188804 254572
rect 187752 254532 187758 254544
rect 188798 254532 188804 254544
rect 188856 254572 188862 254584
rect 197998 254572 198004 254584
rect 188856 254544 198004 254572
rect 188856 254532 188862 254544
rect 197998 254532 198004 254544
rect 198056 254532 198062 254584
rect 56318 253920 56324 253972
rect 56376 253960 56382 253972
rect 66806 253960 66812 253972
rect 56376 253932 66812 253960
rect 56376 253920 56382 253932
rect 66806 253920 66812 253932
rect 66864 253920 66870 253972
rect 162118 253920 162124 253972
rect 162176 253960 162182 253972
rect 163682 253960 163688 253972
rect 162176 253932 163688 253960
rect 162176 253920 162182 253932
rect 163682 253920 163688 253932
rect 163740 253920 163746 253972
rect 165062 253920 165068 253972
rect 165120 253960 165126 253972
rect 187694 253960 187700 253972
rect 165120 253932 187700 253960
rect 165120 253920 165126 253932
rect 187694 253920 187700 253932
rect 187752 253920 187758 253972
rect 193030 253920 193036 253972
rect 193088 253960 193094 253972
rect 197354 253960 197360 253972
rect 193088 253932 197360 253960
rect 193088 253920 193094 253932
rect 197354 253920 197360 253932
rect 197412 253920 197418 253972
rect 54938 253852 54944 253904
rect 54996 253892 55002 253904
rect 57146 253892 57152 253904
rect 54996 253864 57152 253892
rect 54996 253852 55002 253864
rect 57146 253852 57152 253864
rect 57204 253852 57210 253904
rect 245930 253852 245936 253904
rect 245988 253892 245994 253904
rect 256878 253892 256884 253904
rect 245988 253864 256884 253892
rect 245988 253852 245994 253864
rect 256878 253852 256884 253864
rect 256936 253852 256942 253904
rect 157242 253580 157248 253632
rect 157300 253620 157306 253632
rect 162762 253620 162768 253632
rect 157300 253592 162768 253620
rect 157300 253580 157306 253592
rect 162762 253580 162768 253592
rect 162820 253580 162826 253632
rect 54938 253172 54944 253224
rect 54996 253212 55002 253224
rect 66898 253212 66904 253224
rect 54996 253184 66904 253212
rect 54996 253172 55002 253184
rect 66898 253172 66904 253184
rect 66956 253172 66962 253224
rect 160738 253172 160744 253224
rect 160796 253212 160802 253224
rect 168374 253212 168380 253224
rect 160796 253184 168380 253212
rect 160796 253172 160802 253184
rect 168374 253172 168380 253184
rect 168432 253172 168438 253224
rect 256878 253172 256884 253224
rect 256936 253212 256942 253224
rect 294046 253212 294052 253224
rect 256936 253184 294052 253212
rect 256936 253172 256942 253184
rect 294046 253172 294052 253184
rect 294104 253172 294110 253224
rect 187602 252628 187608 252680
rect 187660 252668 187666 252680
rect 197354 252668 197360 252680
rect 187660 252640 197360 252668
rect 187660 252628 187666 252640
rect 197354 252628 197360 252640
rect 197412 252628 197418 252680
rect 57146 252560 57152 252612
rect 57204 252600 57210 252612
rect 57606 252600 57612 252612
rect 57204 252572 57612 252600
rect 57204 252560 57210 252572
rect 57606 252560 57612 252572
rect 57664 252600 57670 252612
rect 66806 252600 66812 252612
rect 57664 252572 66812 252600
rect 57664 252560 57670 252572
rect 66806 252560 66812 252572
rect 66864 252560 66870 252612
rect 168374 252560 168380 252612
rect 168432 252600 168438 252612
rect 169570 252600 169576 252612
rect 168432 252572 169576 252600
rect 168432 252560 168438 252572
rect 169570 252560 169576 252572
rect 169628 252600 169634 252612
rect 197446 252600 197452 252612
rect 169628 252572 197452 252600
rect 169628 252560 169634 252572
rect 197446 252560 197452 252572
rect 197504 252560 197510 252612
rect 245838 252492 245844 252544
rect 245896 252532 245902 252544
rect 262214 252532 262220 252544
rect 245896 252504 262220 252532
rect 245896 252492 245902 252504
rect 262214 252492 262220 252504
rect 262272 252532 262278 252544
rect 262674 252532 262680 252544
rect 262272 252504 262680 252532
rect 262272 252492 262278 252504
rect 262674 252492 262680 252504
rect 262732 252492 262738 252544
rect 245930 252288 245936 252340
rect 245988 252328 245994 252340
rect 248690 252328 248696 252340
rect 245988 252300 248696 252328
rect 245988 252288 245994 252300
rect 248690 252288 248696 252300
rect 248748 252288 248754 252340
rect 173802 251812 173808 251864
rect 173860 251852 173866 251864
rect 187694 251852 187700 251864
rect 173860 251824 187700 251852
rect 173860 251812 173866 251824
rect 187694 251812 187700 251824
rect 187752 251812 187758 251864
rect 262674 251812 262680 251864
rect 262732 251852 262738 251864
rect 583570 251852 583576 251864
rect 262732 251824 583576 251852
rect 262732 251812 262738 251824
rect 583570 251812 583576 251824
rect 583628 251812 583634 251864
rect 157242 251268 157248 251320
rect 157300 251308 157306 251320
rect 169754 251308 169760 251320
rect 157300 251280 169760 251308
rect 157300 251268 157306 251280
rect 169754 251268 169760 251280
rect 169812 251268 169818 251320
rect 157150 251200 157156 251252
rect 157208 251240 157214 251252
rect 180058 251240 180064 251252
rect 157208 251212 180064 251240
rect 157208 251200 157214 251212
rect 180058 251200 180064 251212
rect 180116 251200 180122 251252
rect 187694 251200 187700 251252
rect 187752 251240 187758 251252
rect 188890 251240 188896 251252
rect 187752 251212 188896 251240
rect 187752 251200 187758 251212
rect 188890 251200 188896 251212
rect 188948 251240 188954 251252
rect 197354 251240 197360 251252
rect 188948 251212 197360 251240
rect 188948 251200 188954 251212
rect 197354 251200 197360 251212
rect 197412 251200 197418 251252
rect 245654 250520 245660 250572
rect 245712 250560 245718 250572
rect 269850 250560 269856 250572
rect 245712 250532 269856 250560
rect 245712 250520 245718 250532
rect 269850 250520 269856 250532
rect 269908 250520 269914 250572
rect 170582 250452 170588 250504
rect 170640 250492 170646 250504
rect 180334 250492 180340 250504
rect 170640 250464 180340 250492
rect 170640 250452 170646 250464
rect 180334 250452 180340 250464
rect 180392 250452 180398 250504
rect 185670 250452 185676 250504
rect 185728 250492 185734 250504
rect 197078 250492 197084 250504
rect 185728 250464 197084 250492
rect 185728 250452 185734 250464
rect 197078 250452 197084 250464
rect 197136 250452 197142 250504
rect 265618 250452 265624 250504
rect 265676 250492 265682 250504
rect 289814 250492 289820 250504
rect 265676 250464 289820 250492
rect 265676 250452 265682 250464
rect 289814 250452 289820 250464
rect 289872 250452 289878 250504
rect 60366 249772 60372 249824
rect 60424 249812 60430 249824
rect 66438 249812 66444 249824
rect 60424 249784 66444 249812
rect 60424 249772 60430 249784
rect 66438 249772 66444 249784
rect 66496 249772 66502 249824
rect 157242 249772 157248 249824
rect 157300 249812 157306 249824
rect 186958 249812 186964 249824
rect 157300 249784 186964 249812
rect 157300 249772 157306 249784
rect 186958 249772 186964 249784
rect 187016 249772 187022 249824
rect 191190 249772 191196 249824
rect 191248 249812 191254 249824
rect 197354 249812 197360 249824
rect 191248 249784 197360 249812
rect 191248 249772 191254 249784
rect 197354 249772 197360 249784
rect 197412 249772 197418 249824
rect 192662 249704 192668 249756
rect 192720 249744 192726 249756
rect 195882 249744 195888 249756
rect 192720 249716 195888 249744
rect 192720 249704 192726 249716
rect 195882 249704 195888 249716
rect 195940 249704 195946 249756
rect 191374 249636 191380 249688
rect 191432 249676 191438 249688
rect 193122 249676 193128 249688
rect 191432 249648 193128 249676
rect 191432 249636 191438 249648
rect 193122 249636 193128 249648
rect 193180 249676 193186 249688
rect 197354 249676 197360 249688
rect 193180 249648 197360 249676
rect 193180 249636 193186 249648
rect 197354 249636 197360 249648
rect 197412 249636 197418 249688
rect 245930 249636 245936 249688
rect 245988 249676 245994 249688
rect 249886 249676 249892 249688
rect 245988 249648 249892 249676
rect 245988 249636 245994 249648
rect 249886 249636 249892 249648
rect 249944 249636 249950 249688
rect 156966 249364 156972 249416
rect 157024 249404 157030 249416
rect 159634 249404 159640 249416
rect 157024 249376 159640 249404
rect 157024 249364 157030 249376
rect 159634 249364 159640 249376
rect 159692 249364 159698 249416
rect 169018 249024 169024 249076
rect 169076 249064 169082 249076
rect 191282 249064 191288 249076
rect 169076 249036 191288 249064
rect 169076 249024 169082 249036
rect 191282 249024 191288 249036
rect 191340 249024 191346 249076
rect 195882 248684 195888 248736
rect 195940 248724 195946 248736
rect 197354 248724 197360 248736
rect 195940 248696 197360 248724
rect 195940 248684 195946 248696
rect 197354 248684 197360 248696
rect 197412 248684 197418 248736
rect 156506 248412 156512 248464
rect 156564 248452 156570 248464
rect 172514 248452 172520 248464
rect 156564 248424 172520 248452
rect 156564 248412 156570 248424
rect 172514 248412 172520 248424
rect 172572 248412 172578 248464
rect 156230 247664 156236 247716
rect 156288 247704 156294 247716
rect 164970 247704 164976 247716
rect 156288 247676 164976 247704
rect 156288 247664 156294 247676
rect 164970 247664 164976 247676
rect 165028 247664 165034 247716
rect 185854 247664 185860 247716
rect 185912 247704 185918 247716
rect 199562 247704 199568 247716
rect 185912 247676 199568 247704
rect 185912 247664 185918 247676
rect 199562 247664 199568 247676
rect 199620 247664 199626 247716
rect 245930 247664 245936 247716
rect 245988 247704 245994 247716
rect 582834 247704 582840 247716
rect 245988 247676 582840 247704
rect 245988 247664 245994 247676
rect 582834 247664 582840 247676
rect 582892 247664 582898 247716
rect 50982 247052 50988 247104
rect 51040 247092 51046 247104
rect 66806 247092 66812 247104
rect 51040 247064 66812 247092
rect 51040 247052 51046 247064
rect 66806 247052 66812 247064
rect 66864 247052 66870 247104
rect 164142 247052 164148 247104
rect 164200 247092 164206 247104
rect 185854 247092 185860 247104
rect 164200 247064 185860 247092
rect 164200 247052 164206 247064
rect 185854 247052 185860 247064
rect 185912 247092 185918 247104
rect 186222 247092 186228 247104
rect 185912 247064 186228 247092
rect 185912 247052 185918 247064
rect 186222 247052 186228 247064
rect 186280 247052 186286 247104
rect 187142 247052 187148 247104
rect 187200 247092 187206 247104
rect 197354 247092 197360 247104
rect 187200 247064 197360 247092
rect 187200 247052 187206 247064
rect 197354 247052 197360 247064
rect 197412 247052 197418 247104
rect 171962 246304 171968 246356
rect 172020 246344 172026 246356
rect 189810 246344 189816 246356
rect 172020 246316 189816 246344
rect 172020 246304 172026 246316
rect 189810 246304 189816 246316
rect 189868 246304 189874 246356
rect 157242 246032 157248 246084
rect 157300 246072 157306 246084
rect 160830 246072 160836 246084
rect 157300 246044 160836 246072
rect 157300 246032 157306 246044
rect 160830 246032 160836 246044
rect 160888 246032 160894 246084
rect 246390 245692 246396 245744
rect 246448 245732 246454 245744
rect 247218 245732 247224 245744
rect 246448 245704 247224 245732
rect 246448 245692 246454 245704
rect 247218 245692 247224 245704
rect 247276 245732 247282 245744
rect 247276 245704 258074 245732
rect 247276 245692 247282 245704
rect 158254 245624 158260 245676
rect 158312 245664 158318 245676
rect 191742 245664 191748 245676
rect 158312 245636 191748 245664
rect 158312 245624 158318 245636
rect 191742 245624 191748 245636
rect 191800 245664 191806 245676
rect 197354 245664 197360 245676
rect 191800 245636 197360 245664
rect 191800 245624 191806 245636
rect 197354 245624 197360 245636
rect 197412 245624 197418 245676
rect 245838 245624 245844 245676
rect 245896 245664 245902 245676
rect 248598 245664 248604 245676
rect 245896 245636 248604 245664
rect 245896 245624 245902 245636
rect 248598 245624 248604 245636
rect 248656 245624 248662 245676
rect 258046 245664 258074 245704
rect 298186 245664 298192 245676
rect 258046 245636 298192 245664
rect 298186 245624 298192 245636
rect 298244 245624 298250 245676
rect 53650 244876 53656 244928
rect 53708 244916 53714 244928
rect 66070 244916 66076 244928
rect 53708 244888 66076 244916
rect 53708 244876 53714 244888
rect 66070 244876 66076 244888
rect 66128 244916 66134 244928
rect 66622 244916 66628 244928
rect 66128 244888 66628 244916
rect 66128 244876 66134 244888
rect 66622 244876 66628 244888
rect 66680 244876 66686 244928
rect 245930 244400 245936 244452
rect 245988 244440 245994 244452
rect 248690 244440 248696 244452
rect 245988 244412 248696 244440
rect 245988 244400 245994 244412
rect 248690 244400 248696 244412
rect 248748 244400 248754 244452
rect 157978 244332 157984 244384
rect 158036 244372 158042 244384
rect 193398 244372 193404 244384
rect 158036 244344 193404 244372
rect 158036 244332 158042 244344
rect 193398 244332 193404 244344
rect 193456 244332 193462 244384
rect 155678 244264 155684 244316
rect 155736 244304 155742 244316
rect 198826 244304 198832 244316
rect 155736 244276 198832 244304
rect 155736 244264 155742 244276
rect 198826 244264 198832 244276
rect 198884 244264 198890 244316
rect 192478 244128 192484 244180
rect 192536 244168 192542 244180
rect 197170 244168 197176 244180
rect 192536 244140 197176 244168
rect 192536 244128 192542 244140
rect 197170 244128 197176 244140
rect 197228 244168 197234 244180
rect 197446 244168 197452 244180
rect 197228 244140 197452 244168
rect 197228 244128 197234 244140
rect 197446 244128 197452 244140
rect 197504 244128 197510 244180
rect 193398 243584 193404 243636
rect 193456 243624 193462 243636
rect 197354 243624 197360 243636
rect 193456 243596 197360 243624
rect 193456 243584 193462 243596
rect 197354 243584 197360 243596
rect 197412 243584 197418 243636
rect 154942 243516 154948 243568
rect 155000 243556 155006 243568
rect 164234 243556 164240 243568
rect 155000 243528 164240 243556
rect 155000 243516 155006 243528
rect 164234 243516 164240 243528
rect 164292 243556 164298 243568
rect 164970 243556 164976 243568
rect 164292 243528 164976 243556
rect 164292 243516 164298 243528
rect 164970 243516 164976 243528
rect 165028 243516 165034 243568
rect 172514 243516 172520 243568
rect 172572 243556 172578 243568
rect 194042 243556 194048 243568
rect 172572 243528 194048 243556
rect 172572 243516 172578 243528
rect 194042 243516 194048 243528
rect 194100 243516 194106 243568
rect 63402 242904 63408 242956
rect 63460 242944 63466 242956
rect 66806 242944 66812 242956
rect 63460 242916 66812 242944
rect 63460 242904 63466 242916
rect 66806 242904 66812 242916
rect 66864 242904 66870 242956
rect 156046 242904 156052 242956
rect 156104 242944 156110 242956
rect 192662 242944 192668 242956
rect 156104 242916 192668 242944
rect 156104 242904 156110 242916
rect 192662 242904 192668 242916
rect 192720 242904 192726 242956
rect 244458 242904 244464 242956
rect 244516 242944 244522 242956
rect 244642 242944 244648 242956
rect 244516 242916 244648 242944
rect 244516 242904 244522 242916
rect 244642 242904 244648 242916
rect 244700 242944 244706 242956
rect 265618 242944 265624 242956
rect 244700 242916 265624 242944
rect 244700 242904 244706 242916
rect 265618 242904 265624 242916
rect 265676 242904 265682 242956
rect 164142 242264 164148 242276
rect 152568 242236 164148 242264
rect 64506 242156 64512 242208
rect 64564 242196 64570 242208
rect 64564 242168 64874 242196
rect 64564 242156 64570 242168
rect 64846 242060 64874 242168
rect 82814 242060 82820 242072
rect 64846 242032 82820 242060
rect 82814 242020 82820 242032
rect 82872 242020 82878 242072
rect 152458 242020 152464 242072
rect 152516 242060 152522 242072
rect 152568 242060 152596 242236
rect 164142 242224 164148 242236
rect 164200 242224 164206 242276
rect 269942 242224 269948 242276
rect 270000 242264 270006 242276
rect 285674 242264 285680 242276
rect 270000 242236 285680 242264
rect 270000 242224 270006 242236
rect 285674 242224 285680 242236
rect 285732 242224 285738 242276
rect 168374 242156 168380 242208
rect 168432 242196 168438 242208
rect 169662 242196 169668 242208
rect 168432 242168 169668 242196
rect 168432 242156 168438 242168
rect 169662 242156 169668 242168
rect 169720 242196 169726 242208
rect 197354 242196 197360 242208
rect 169720 242168 197360 242196
rect 169720 242156 169726 242168
rect 197354 242156 197360 242168
rect 197412 242156 197418 242208
rect 245102 242156 245108 242208
rect 245160 242196 245166 242208
rect 252738 242196 252744 242208
rect 245160 242168 252744 242196
rect 245160 242156 245166 242168
rect 252738 242156 252744 242168
rect 252796 242156 252802 242208
rect 261570 242156 261576 242208
rect 261628 242196 261634 242208
rect 278222 242196 278228 242208
rect 261628 242168 278228 242196
rect 261628 242156 261634 242168
rect 278222 242156 278228 242168
rect 278280 242156 278286 242208
rect 152516 242032 152596 242060
rect 152516 242020 152522 242032
rect 154114 242020 154120 242072
rect 154172 242060 154178 242072
rect 165062 242060 165068 242072
rect 154172 242032 165068 242060
rect 154172 242020 154178 242032
rect 165062 242020 165068 242032
rect 165120 242020 165126 242072
rect 70394 241816 70400 241868
rect 70452 241856 70458 241868
rect 71038 241856 71044 241868
rect 70452 241828 71044 241856
rect 70452 241816 70458 241828
rect 71038 241816 71044 241828
rect 71096 241816 71102 241868
rect 149146 241544 149152 241596
rect 149204 241584 149210 241596
rect 154022 241584 154028 241596
rect 149204 241556 154028 241584
rect 149204 241544 149210 241556
rect 154022 241544 154028 241556
rect 154080 241544 154086 241596
rect 163682 241476 163688 241528
rect 163740 241516 163746 241528
rect 191650 241516 191656 241528
rect 163740 241488 191656 241516
rect 163740 241476 163746 241488
rect 191650 241476 191656 241488
rect 191708 241476 191714 241528
rect 195330 241476 195336 241528
rect 195388 241516 195394 241528
rect 197538 241516 197544 241528
rect 195388 241488 197544 241516
rect 195388 241476 195394 241488
rect 197538 241476 197544 241488
rect 197596 241476 197602 241528
rect 245930 241476 245936 241528
rect 245988 241516 245994 241528
rect 255498 241516 255504 241528
rect 245988 241488 255504 241516
rect 245988 241476 245994 241488
rect 255498 241476 255504 241488
rect 255556 241476 255562 241528
rect 141464 241408 141470 241460
rect 141522 241448 141528 241460
rect 149054 241448 149060 241460
rect 141522 241420 149060 241448
rect 141522 241408 141528 241420
rect 149054 241408 149060 241420
rect 149112 241408 149118 241460
rect 193858 241408 193864 241460
rect 193916 241448 193922 241460
rect 197354 241448 197360 241460
rect 193916 241420 197360 241448
rect 193916 241408 193922 241420
rect 197354 241408 197360 241420
rect 197412 241408 197418 241460
rect 3418 241068 3424 241120
rect 3476 241108 3482 241120
rect 7558 241108 7564 241120
rect 3476 241080 7564 241108
rect 3476 241068 3482 241080
rect 7558 241068 7564 241080
rect 7616 241068 7622 241120
rect 115842 240796 115848 240848
rect 115900 240836 115906 240848
rect 155678 240836 155684 240848
rect 115900 240808 155684 240836
rect 115900 240796 115906 240808
rect 155678 240796 155684 240808
rect 155736 240796 155742 240848
rect 65978 240728 65984 240780
rect 66036 240768 66042 240780
rect 76650 240768 76656 240780
rect 66036 240740 76656 240768
rect 66036 240728 66042 240740
rect 76650 240728 76656 240740
rect 76708 240728 76714 240780
rect 82814 240728 82820 240780
rect 82872 240768 82878 240780
rect 128814 240768 128820 240780
rect 82872 240740 128820 240768
rect 82872 240728 82878 240740
rect 128814 240728 128820 240740
rect 128872 240728 128878 240780
rect 149514 240728 149520 240780
rect 149572 240768 149578 240780
rect 199562 240768 199568 240780
rect 149572 240740 199568 240768
rect 149572 240728 149578 240740
rect 199562 240728 199568 240740
rect 199620 240728 199626 240780
rect 198734 240320 198740 240372
rect 198792 240360 198798 240372
rect 198792 240332 202184 240360
rect 198792 240320 198798 240332
rect 200114 240252 200120 240304
rect 200172 240292 200178 240304
rect 200172 240264 200344 240292
rect 200172 240252 200178 240264
rect 200316 240168 200344 240264
rect 202156 240168 202184 240332
rect 67818 240116 67824 240168
rect 67876 240156 67882 240168
rect 76558 240156 76564 240168
rect 67876 240128 76564 240156
rect 67876 240116 67882 240128
rect 76558 240116 76564 240128
rect 76616 240116 76622 240168
rect 104894 240116 104900 240168
rect 104952 240156 104958 240168
rect 105446 240156 105452 240168
rect 104952 240128 105452 240156
rect 104952 240116 104958 240128
rect 105446 240116 105452 240128
rect 105504 240116 105510 240168
rect 198642 240116 198648 240168
rect 198700 240156 198706 240168
rect 200114 240156 200120 240168
rect 198700 240128 200120 240156
rect 198700 240116 198706 240128
rect 200114 240116 200120 240128
rect 200172 240116 200178 240168
rect 200298 240116 200304 240168
rect 200356 240116 200362 240168
rect 202138 240116 202144 240168
rect 202196 240116 202202 240168
rect 242250 240116 242256 240168
rect 242308 240156 242314 240168
rect 244090 240156 244096 240168
rect 242308 240128 244096 240156
rect 242308 240116 242314 240128
rect 244090 240116 244096 240128
rect 244148 240116 244154 240168
rect 67542 240048 67548 240100
rect 67600 240088 67606 240100
rect 69750 240088 69756 240100
rect 67600 240060 69756 240088
rect 67600 240048 67606 240060
rect 69750 240048 69756 240060
rect 69808 240048 69814 240100
rect 70302 240048 70308 240100
rect 70360 240088 70366 240100
rect 115842 240088 115848 240100
rect 70360 240060 115848 240088
rect 70360 240048 70366 240060
rect 115842 240048 115848 240060
rect 115900 240048 115906 240100
rect 117222 240048 117228 240100
rect 117280 240088 117286 240100
rect 224310 240088 224316 240100
rect 117280 240060 224316 240088
rect 117280 240048 117286 240060
rect 224310 240048 224316 240060
rect 224368 240048 224374 240100
rect 240870 240048 240876 240100
rect 240928 240088 240934 240100
rect 243906 240088 243912 240100
rect 240928 240060 243912 240088
rect 240928 240048 240934 240060
rect 243906 240048 243912 240060
rect 243964 240048 243970 240100
rect 252830 240088 252836 240100
rect 248386 240060 252836 240088
rect 79042 239980 79048 240032
rect 79100 240020 79106 240032
rect 79870 240020 79876 240032
rect 79100 239992 79876 240020
rect 79100 239980 79106 239992
rect 79870 239980 79876 239992
rect 79928 239980 79934 240032
rect 80514 239980 80520 240032
rect 80572 240020 80578 240032
rect 81342 240020 81348 240032
rect 80572 239992 81348 240020
rect 80572 239980 80578 239992
rect 81342 239980 81348 239992
rect 81400 239980 81406 240032
rect 81526 239980 81532 240032
rect 81584 240020 81590 240032
rect 82722 240020 82728 240032
rect 81584 239992 82728 240020
rect 81584 239980 81590 239992
rect 82722 239980 82728 239992
rect 82780 239980 82786 240032
rect 86034 239980 86040 240032
rect 86092 240020 86098 240032
rect 86862 240020 86868 240032
rect 86092 239992 86868 240020
rect 86092 239980 86098 239992
rect 86862 239980 86868 239992
rect 86920 239980 86926 240032
rect 90450 239980 90456 240032
rect 90508 240020 90514 240032
rect 90910 240020 90916 240032
rect 90508 239992 90916 240020
rect 90508 239980 90514 239992
rect 90910 239980 90916 239992
rect 90968 239980 90974 240032
rect 121730 239980 121736 240032
rect 121788 240020 121794 240032
rect 122742 240020 122748 240032
rect 121788 239992 122748 240020
rect 121788 239980 121794 239992
rect 122742 239980 122748 239992
rect 122800 239980 122806 240032
rect 127434 239980 127440 240032
rect 127492 240020 127498 240032
rect 128262 240020 128268 240032
rect 127492 239992 128268 240020
rect 127492 239980 127498 239992
rect 128262 239980 128268 239992
rect 128320 239980 128326 240032
rect 131850 239980 131856 240032
rect 131908 240020 131914 240032
rect 132310 240020 132316 240032
rect 131908 239992 132316 240020
rect 131908 239980 131914 239992
rect 132310 239980 132316 239992
rect 132368 239980 132374 240032
rect 228726 240020 228732 240032
rect 132466 239992 228732 240020
rect 128906 239912 128912 239964
rect 128964 239952 128970 239964
rect 129642 239952 129648 239964
rect 128964 239924 129648 239952
rect 128964 239912 128970 239924
rect 129642 239912 129648 239924
rect 129700 239912 129706 239964
rect 126146 239844 126152 239896
rect 126204 239884 126210 239896
rect 132466 239884 132494 239992
rect 228726 239980 228732 239992
rect 228784 239980 228790 240032
rect 240042 239980 240048 240032
rect 240100 240020 240106 240032
rect 248386 240020 248414 240060
rect 252830 240048 252836 240060
rect 252888 240048 252894 240100
rect 240100 239992 248414 240020
rect 240100 239980 240106 239992
rect 138106 239912 138112 239964
rect 138164 239952 138170 239964
rect 138934 239952 138940 239964
rect 138164 239924 138940 239952
rect 138164 239912 138170 239924
rect 138934 239912 138940 239924
rect 138992 239912 138998 239964
rect 142246 239912 142252 239964
rect 142304 239952 142310 239964
rect 143350 239952 143356 239964
rect 142304 239924 143356 239952
rect 142304 239912 142310 239924
rect 143350 239912 143356 239924
rect 143408 239912 143414 239964
rect 145282 239912 145288 239964
rect 145340 239952 145346 239964
rect 146018 239952 146024 239964
rect 145340 239924 146024 239952
rect 145340 239912 145346 239924
rect 146018 239912 146024 239924
rect 146076 239912 146082 239964
rect 126204 239856 132494 239884
rect 126204 239844 126210 239856
rect 106826 239776 106832 239828
rect 106884 239816 106890 239828
rect 107562 239816 107568 239828
rect 106884 239788 107568 239816
rect 106884 239776 106890 239788
rect 107562 239776 107568 239788
rect 107620 239776 107626 239828
rect 148226 239776 148232 239828
rect 148284 239816 148290 239828
rect 148962 239816 148968 239828
rect 148284 239788 148968 239816
rect 148284 239776 148290 239788
rect 148962 239776 148968 239788
rect 149020 239776 149026 239828
rect 101122 239640 101128 239692
rect 101180 239680 101186 239692
rect 102042 239680 102048 239692
rect 101180 239652 102048 239680
rect 101180 239640 101186 239652
rect 102042 239640 102048 239652
rect 102100 239640 102106 239692
rect 120166 239640 120172 239692
rect 120224 239680 120230 239692
rect 121362 239680 121368 239692
rect 120224 239652 121368 239680
rect 120224 239640 120230 239652
rect 121362 239640 121368 239652
rect 121420 239640 121426 239692
rect 88978 239504 88984 239556
rect 89036 239544 89042 239556
rect 89530 239544 89536 239556
rect 89036 239516 89536 239544
rect 89036 239504 89042 239516
rect 89530 239504 89536 239516
rect 89588 239504 89594 239556
rect 99374 239504 99380 239556
rect 99432 239544 99438 239556
rect 100662 239544 100668 239556
rect 99432 239516 100668 239544
rect 99432 239504 99438 239516
rect 100662 239504 100668 239516
rect 100720 239504 100726 239556
rect 107746 239504 107752 239556
rect 107804 239544 107810 239556
rect 108390 239544 108396 239556
rect 107804 239516 108396 239544
rect 107804 239504 107810 239516
rect 108390 239504 108396 239516
rect 108448 239504 108454 239556
rect 109586 239504 109592 239556
rect 109644 239544 109650 239556
rect 110230 239544 110236 239556
rect 109644 239516 110236 239544
rect 109644 239504 109650 239516
rect 110230 239504 110236 239516
rect 110288 239504 110294 239556
rect 111058 239504 111064 239556
rect 111116 239544 111122 239556
rect 111610 239544 111616 239556
rect 111116 239516 111616 239544
rect 111116 239504 111122 239516
rect 111610 239504 111616 239516
rect 111668 239504 111674 239556
rect 71682 239368 71688 239420
rect 71740 239408 71746 239420
rect 79318 239408 79324 239420
rect 71740 239380 79324 239408
rect 71740 239368 71746 239380
rect 79318 239368 79324 239380
rect 79376 239368 79382 239420
rect 124674 239368 124680 239420
rect 124732 239408 124738 239420
rect 125410 239408 125416 239420
rect 124732 239380 125416 239408
rect 124732 239368 124738 239380
rect 125410 239368 125416 239380
rect 125468 239368 125474 239420
rect 97626 239300 97632 239352
rect 97684 239340 97690 239352
rect 104158 239340 104164 239352
rect 97684 239312 104164 239340
rect 97684 239300 97690 239312
rect 104158 239300 104164 239312
rect 104216 239300 104222 239352
rect 115290 239232 115296 239284
rect 115348 239272 115354 239284
rect 115842 239272 115848 239284
rect 115348 239244 115848 239272
rect 115348 239232 115354 239244
rect 115842 239232 115848 239244
rect 115900 239232 115906 239284
rect 130378 239232 130384 239284
rect 130436 239272 130442 239284
rect 130930 239272 130936 239284
rect 130436 239244 130936 239272
rect 130436 239232 130442 239244
rect 130930 239232 130936 239244
rect 130988 239232 130994 239284
rect 133138 239164 133144 239216
rect 133196 239204 133202 239216
rect 133690 239204 133696 239216
rect 133196 239176 133696 239204
rect 133196 239164 133202 239176
rect 133690 239164 133696 239176
rect 133748 239164 133754 239216
rect 134610 239164 134616 239216
rect 134668 239204 134674 239216
rect 135162 239204 135168 239216
rect 134668 239176 135168 239204
rect 134668 239164 134674 239176
rect 135162 239164 135168 239176
rect 135220 239164 135226 239216
rect 141050 239096 141056 239148
rect 141108 239136 141114 239148
rect 142062 239136 142068 239148
rect 141108 239108 142068 239136
rect 141108 239096 141114 239108
rect 142062 239096 142068 239108
rect 142120 239096 142126 239148
rect 143994 239096 144000 239148
rect 144052 239136 144058 239148
rect 144730 239136 144736 239148
rect 144052 239108 144736 239136
rect 144052 239096 144058 239108
rect 144730 239096 144736 239108
rect 144788 239096 144794 239148
rect 149054 239096 149060 239148
rect 149112 239136 149118 239148
rect 149606 239136 149612 239148
rect 149112 239108 149612 239136
rect 149112 239096 149118 239108
rect 149606 239096 149612 239108
rect 149664 239096 149670 239148
rect 153930 239096 153936 239148
rect 153988 239136 153994 239148
rect 154482 239136 154488 239148
rect 153988 239108 154488 239136
rect 153988 239096 153994 239108
rect 154482 239096 154488 239108
rect 154540 239096 154546 239148
rect 226886 238756 226892 238808
rect 226944 238796 226950 238808
rect 238938 238796 238944 238808
rect 226944 238768 238944 238796
rect 226944 238756 226950 238768
rect 238938 238756 238944 238768
rect 238996 238796 239002 238808
rect 240042 238796 240048 238808
rect 238996 238768 240048 238796
rect 238996 238756 239002 238768
rect 240042 238756 240048 238768
rect 240100 238756 240106 238808
rect 219434 238688 219440 238740
rect 219492 238728 219498 238740
rect 222838 238728 222844 238740
rect 219492 238700 222844 238728
rect 219492 238688 219498 238700
rect 222838 238688 222844 238700
rect 222896 238688 222902 238740
rect 242158 238688 242164 238740
rect 242216 238728 242222 238740
rect 248506 238728 248512 238740
rect 242216 238700 248512 238728
rect 242216 238688 242222 238700
rect 248506 238688 248512 238700
rect 248564 238688 248570 238740
rect 107654 238620 107660 238672
rect 107712 238660 107718 238672
rect 219894 238660 219900 238672
rect 107712 238632 219900 238660
rect 107712 238620 107718 238632
rect 219894 238620 219900 238632
rect 219952 238620 219958 238672
rect 60366 238076 60372 238128
rect 60424 238116 60430 238128
rect 73798 238116 73804 238128
rect 60424 238088 73804 238116
rect 60424 238076 60430 238088
rect 73798 238076 73804 238088
rect 73856 238076 73862 238128
rect 224310 238076 224316 238128
rect 224368 238116 224374 238128
rect 236638 238116 236644 238128
rect 224368 238088 236644 238116
rect 224368 238076 224374 238088
rect 236638 238076 236644 238088
rect 236696 238076 236702 238128
rect 67910 238008 67916 238060
rect 67968 238048 67974 238060
rect 108298 238048 108304 238060
rect 67968 238020 108304 238048
rect 67968 238008 67974 238020
rect 108298 238008 108304 238020
rect 108356 238008 108362 238060
rect 215294 238008 215300 238060
rect 215352 238048 215358 238060
rect 244458 238048 244464 238060
rect 215352 238020 244464 238048
rect 215352 238008 215358 238020
rect 244458 238008 244464 238020
rect 244516 238008 244522 238060
rect 199470 237804 199476 237856
rect 199528 237844 199534 237856
rect 199930 237844 199936 237856
rect 199528 237816 199936 237844
rect 199528 237804 199534 237816
rect 199930 237804 199936 237816
rect 199988 237844 199994 237856
rect 201034 237844 201040 237856
rect 199988 237816 201040 237844
rect 199988 237804 199994 237816
rect 201034 237804 201040 237816
rect 201092 237804 201098 237856
rect 230566 237804 230572 237856
rect 230624 237844 230630 237856
rect 231762 237844 231768 237856
rect 230624 237816 231768 237844
rect 230624 237804 230630 237816
rect 231762 237804 231768 237816
rect 231820 237804 231826 237856
rect 84194 237668 84200 237720
rect 84252 237708 84258 237720
rect 93118 237708 93124 237720
rect 84252 237680 93124 237708
rect 84252 237668 84258 237680
rect 93118 237668 93124 237680
rect 93176 237668 93182 237720
rect 200114 237396 200120 237448
rect 200172 237436 200178 237448
rect 201586 237436 201592 237448
rect 200172 237408 201592 237436
rect 200172 237396 200178 237408
rect 201586 237396 201592 237408
rect 201644 237396 201650 237448
rect 206830 237396 206836 237448
rect 206888 237436 206894 237448
rect 207658 237436 207664 237448
rect 206888 237408 207664 237436
rect 206888 237396 206894 237408
rect 207658 237396 207664 237408
rect 207716 237396 207722 237448
rect 207934 237396 207940 237448
rect 207992 237436 207998 237448
rect 209038 237436 209044 237448
rect 207992 237408 209044 237436
rect 207992 237396 207998 237408
rect 209038 237396 209044 237408
rect 209096 237396 209102 237448
rect 211246 237396 211252 237448
rect 211304 237436 211310 237448
rect 211798 237436 211804 237448
rect 211304 237408 211804 237436
rect 211304 237396 211310 237408
rect 211798 237396 211804 237408
rect 211856 237396 211862 237448
rect 223022 237396 223028 237448
rect 223080 237436 223086 237448
rect 223758 237436 223764 237448
rect 223080 237408 223764 237436
rect 223080 237396 223086 237408
rect 223758 237396 223764 237408
rect 223816 237396 223822 237448
rect 4798 237328 4804 237380
rect 4856 237368 4862 237380
rect 53834 237368 53840 237380
rect 4856 237340 53840 237368
rect 4856 237328 4862 237340
rect 53834 237328 53840 237340
rect 53892 237328 53898 237380
rect 103514 237328 103520 237380
rect 103572 237368 103578 237380
rect 137094 237368 137100 237380
rect 103572 237340 137100 237368
rect 103572 237328 103578 237340
rect 137094 237328 137100 237340
rect 137152 237328 137158 237380
rect 138014 237328 138020 237380
rect 138072 237368 138078 237380
rect 164878 237368 164884 237380
rect 138072 237340 164884 237368
rect 138072 237328 138078 237340
rect 164878 237328 164884 237340
rect 164936 237328 164942 237380
rect 216030 237328 216036 237380
rect 216088 237368 216094 237380
rect 265710 237368 265716 237380
rect 216088 237340 265716 237368
rect 216088 237328 216094 237340
rect 265710 237328 265716 237340
rect 265768 237328 265774 237380
rect 118694 237260 118700 237312
rect 118752 237300 118758 237312
rect 152458 237300 152464 237312
rect 118752 237272 152464 237300
rect 118752 237260 118758 237272
rect 152458 237260 152464 237272
rect 152516 237260 152522 237312
rect 196894 237260 196900 237312
rect 196952 237300 196958 237312
rect 208854 237300 208860 237312
rect 196952 237272 208860 237300
rect 196952 237260 196958 237272
rect 208854 237260 208860 237272
rect 208912 237260 208918 237312
rect 186958 237192 186964 237244
rect 187016 237232 187022 237244
rect 215294 237232 215300 237244
rect 187016 237204 215300 237232
rect 187016 237192 187022 237204
rect 215294 237192 215300 237204
rect 215352 237192 215358 237244
rect 53834 236648 53840 236700
rect 53892 236688 53898 236700
rect 54846 236688 54852 236700
rect 53892 236660 54852 236688
rect 53892 236648 53898 236660
rect 54846 236648 54852 236660
rect 54904 236688 54910 236700
rect 86218 236688 86224 236700
rect 54904 236660 86224 236688
rect 54904 236648 54910 236660
rect 86218 236648 86224 236660
rect 86276 236648 86282 236700
rect 91094 236648 91100 236700
rect 91152 236688 91158 236700
rect 104250 236688 104256 236700
rect 91152 236660 104256 236688
rect 91152 236648 91158 236660
rect 104250 236648 104256 236660
rect 104308 236648 104314 236700
rect 152458 236648 152464 236700
rect 152516 236688 152522 236700
rect 161474 236688 161480 236700
rect 152516 236660 161480 236688
rect 152516 236648 152522 236660
rect 161474 236648 161480 236660
rect 161532 236688 161538 236700
rect 162762 236688 162768 236700
rect 161532 236660 162768 236688
rect 161532 236648 161538 236660
rect 162762 236648 162768 236660
rect 162820 236648 162826 236700
rect 176010 236648 176016 236700
rect 176068 236688 176074 236700
rect 185578 236688 185584 236700
rect 176068 236660 185584 236688
rect 176068 236648 176074 236660
rect 185578 236648 185584 236660
rect 185636 236648 185642 236700
rect 195882 236444 195888 236496
rect 195940 236484 195946 236496
rect 196802 236484 196808 236496
rect 195940 236456 196808 236484
rect 195940 236444 195946 236456
rect 196802 236444 196808 236456
rect 196860 236444 196866 236496
rect 214650 236104 214656 236156
rect 214708 236144 214714 236156
rect 216030 236144 216036 236156
rect 214708 236116 216036 236144
rect 214708 236104 214714 236116
rect 216030 236104 216036 236116
rect 216088 236104 216094 236156
rect 226978 236036 226984 236088
rect 227036 236076 227042 236088
rect 229646 236076 229652 236088
rect 227036 236048 229652 236076
rect 227036 236036 227042 236048
rect 229646 236036 229652 236048
rect 229704 236036 229710 236088
rect 128814 235900 128820 235952
rect 128872 235940 128878 235952
rect 181622 235940 181628 235952
rect 128872 235912 181628 235940
rect 128872 235900 128878 235912
rect 181622 235900 181628 235912
rect 181680 235900 181686 235952
rect 189902 235900 189908 235952
rect 189960 235940 189966 235952
rect 204438 235940 204444 235952
rect 189960 235912 204444 235940
rect 189960 235900 189966 235912
rect 204438 235900 204444 235912
rect 204496 235900 204502 235952
rect 235350 235900 235356 235952
rect 235408 235940 235414 235952
rect 252922 235940 252928 235952
rect 235408 235912 252928 235940
rect 235408 235900 235414 235912
rect 252922 235900 252928 235912
rect 252980 235900 252986 235952
rect 103698 235288 103704 235340
rect 103756 235328 103762 235340
rect 119430 235328 119436 235340
rect 103756 235300 119436 235328
rect 103756 235288 103762 235300
rect 119430 235288 119436 235300
rect 119488 235288 119494 235340
rect 115934 235220 115940 235272
rect 115992 235260 115998 235272
rect 137278 235260 137284 235272
rect 115992 235232 137284 235260
rect 115992 235220 115998 235232
rect 137278 235220 137284 235232
rect 137336 235220 137342 235272
rect 243630 235220 243636 235272
rect 243688 235260 243694 235272
rect 284294 235260 284300 235272
rect 243688 235232 284300 235260
rect 243688 235220 243694 235232
rect 284294 235220 284300 235232
rect 284352 235220 284358 235272
rect 194686 234676 194692 234728
rect 194744 234716 194750 234728
rect 211062 234716 211068 234728
rect 194744 234688 211068 234716
rect 194744 234676 194750 234688
rect 211062 234676 211068 234688
rect 211120 234676 211126 234728
rect 231118 234676 231124 234728
rect 231176 234716 231182 234728
rect 232038 234716 232044 234728
rect 231176 234688 232044 234716
rect 231176 234676 231182 234688
rect 232038 234676 232044 234688
rect 232096 234676 232102 234728
rect 208394 234608 208400 234660
rect 208452 234648 208458 234660
rect 240318 234648 240324 234660
rect 208452 234620 240324 234648
rect 208452 234608 208458 234620
rect 240318 234608 240324 234620
rect 240376 234648 240382 234660
rect 240778 234648 240784 234660
rect 240376 234620 240784 234648
rect 240376 234608 240382 234620
rect 240778 234608 240784 234620
rect 240836 234608 240842 234660
rect 252922 234608 252928 234660
rect 252980 234648 252986 234660
rect 582834 234648 582840 234660
rect 252980 234620 582840 234648
rect 252980 234608 252986 234620
rect 582834 234608 582840 234620
rect 582892 234608 582898 234660
rect 21358 234540 21364 234592
rect 21416 234580 21422 234592
rect 92474 234580 92480 234592
rect 21416 234552 92480 234580
rect 21416 234540 21422 234552
rect 92474 234540 92480 234552
rect 92532 234540 92538 234592
rect 122926 234540 122932 234592
rect 122984 234580 122990 234592
rect 145926 234580 145932 234592
rect 122984 234552 145932 234580
rect 122984 234540 122990 234552
rect 145926 234540 145932 234552
rect 145984 234540 145990 234592
rect 146018 234540 146024 234592
rect 146076 234580 146082 234592
rect 161014 234580 161020 234592
rect 146076 234552 161020 234580
rect 146076 234540 146082 234552
rect 161014 234540 161020 234552
rect 161072 234540 161078 234592
rect 177574 234540 177580 234592
rect 177632 234580 177638 234592
rect 249886 234580 249892 234592
rect 177632 234552 249892 234580
rect 177632 234540 177638 234552
rect 249886 234540 249892 234552
rect 249944 234540 249950 234592
rect 133598 234472 133604 234524
rect 133656 234512 133662 234524
rect 184382 234512 184388 234524
rect 133656 234484 184388 234512
rect 133656 234472 133662 234484
rect 184382 234472 184388 234484
rect 184440 234472 184446 234524
rect 188798 234472 188804 234524
rect 188856 234512 188862 234524
rect 192478 234512 192484 234524
rect 188856 234484 192484 234512
rect 188856 234472 188862 234484
rect 192478 234472 192484 234484
rect 192536 234472 192542 234524
rect 192662 234472 192668 234524
rect 192720 234512 192726 234524
rect 240962 234512 240968 234524
rect 192720 234484 240968 234512
rect 192720 234472 192726 234484
rect 240962 234472 240968 234484
rect 241020 234512 241026 234524
rect 241238 234512 241244 234524
rect 241020 234484 241244 234512
rect 241020 234472 241026 234484
rect 241238 234472 241244 234484
rect 241296 234472 241302 234524
rect 63218 233860 63224 233912
rect 63276 233900 63282 233912
rect 75178 233900 75184 233912
rect 63276 233872 75184 233900
rect 63276 233860 63282 233872
rect 75178 233860 75184 233872
rect 75236 233860 75242 233912
rect 92474 233860 92480 233912
rect 92532 233900 92538 233912
rect 111058 233900 111064 233912
rect 92532 233872 111064 233900
rect 92532 233860 92538 233872
rect 111058 233860 111064 233872
rect 111116 233860 111122 233912
rect 57698 233180 57704 233232
rect 57756 233220 57762 233232
rect 124306 233220 124312 233232
rect 57756 233192 124312 233220
rect 57756 233180 57762 233192
rect 124306 233180 124312 233192
rect 124364 233180 124370 233232
rect 126698 233180 126704 233232
rect 126756 233220 126762 233232
rect 173342 233220 173348 233232
rect 126756 233192 173348 233220
rect 126756 233180 126762 233192
rect 173342 233180 173348 233192
rect 173400 233220 173406 233232
rect 173526 233220 173532 233232
rect 173400 233192 173532 233220
rect 173400 233180 173406 233192
rect 173526 233180 173532 233192
rect 173584 233180 173590 233232
rect 182910 233180 182916 233232
rect 182968 233220 182974 233232
rect 225230 233220 225236 233232
rect 182968 233192 225236 233220
rect 182968 233180 182974 233192
rect 225230 233180 225236 233192
rect 225288 233180 225294 233232
rect 155494 233112 155500 233164
rect 155552 233152 155558 233164
rect 158254 233152 158260 233164
rect 155552 233124 158260 233152
rect 155552 233112 155558 233124
rect 158254 233112 158260 233124
rect 158312 233112 158318 233164
rect 194042 233112 194048 233164
rect 194100 233152 194106 233164
rect 219526 233152 219532 233164
rect 194100 233124 219532 233152
rect 194100 233112 194106 233124
rect 219526 233112 219532 233124
rect 219584 233112 219590 233164
rect 107746 232500 107752 232552
rect 107804 232540 107810 232552
rect 128998 232540 129004 232552
rect 107804 232512 129004 232540
rect 107804 232500 107810 232512
rect 128998 232500 129004 232512
rect 129056 232500 129062 232552
rect 138106 232500 138112 232552
rect 138164 232540 138170 232552
rect 153102 232540 153108 232552
rect 138164 232512 153108 232540
rect 138164 232500 138170 232512
rect 153102 232500 153108 232512
rect 153160 232540 153166 232552
rect 155310 232540 155316 232552
rect 153160 232512 155316 232540
rect 153160 232500 153166 232512
rect 155310 232500 155316 232512
rect 155368 232500 155374 232552
rect 157334 232500 157340 232552
rect 157392 232540 157398 232552
rect 173802 232540 173808 232552
rect 157392 232512 173808 232540
rect 157392 232500 157398 232512
rect 173802 232500 173808 232512
rect 173860 232500 173866 232552
rect 225598 231820 225604 231872
rect 225656 231860 225662 231872
rect 226150 231860 226156 231872
rect 225656 231832 226156 231860
rect 225656 231820 225662 231832
rect 226150 231820 226156 231832
rect 226208 231860 226214 231872
rect 292574 231860 292580 231872
rect 226208 231832 292580 231860
rect 226208 231820 226214 231832
rect 292574 231820 292580 231832
rect 292632 231820 292638 231872
rect 54938 231752 54944 231804
rect 54996 231792 55002 231804
rect 126238 231792 126244 231804
rect 54996 231764 126244 231792
rect 54996 231752 55002 231764
rect 126238 231752 126244 231764
rect 126296 231752 126302 231804
rect 148870 231752 148876 231804
rect 148928 231792 148934 231804
rect 166442 231792 166448 231804
rect 148928 231764 166448 231792
rect 148928 231752 148934 231764
rect 166442 231752 166448 231764
rect 166500 231752 166506 231804
rect 180334 231752 180340 231804
rect 180392 231792 180398 231804
rect 223022 231792 223028 231804
rect 180392 231764 223028 231792
rect 180392 231752 180398 231764
rect 223022 231752 223028 231764
rect 223080 231752 223086 231804
rect 147582 231684 147588 231736
rect 147640 231724 147646 231736
rect 158162 231724 158168 231736
rect 147640 231696 158168 231724
rect 147640 231684 147646 231696
rect 158162 231684 158168 231696
rect 158220 231684 158226 231736
rect 199562 231684 199568 231736
rect 199620 231724 199626 231736
rect 208394 231724 208400 231736
rect 199620 231696 208400 231724
rect 199620 231684 199626 231696
rect 208394 231684 208400 231696
rect 208452 231684 208458 231736
rect 226702 231140 226708 231192
rect 226760 231180 226766 231192
rect 295426 231180 295432 231192
rect 226760 231152 295432 231180
rect 226760 231140 226766 231152
rect 295426 231140 295432 231152
rect 295484 231140 295490 231192
rect 77386 231072 77392 231124
rect 77444 231112 77450 231124
rect 148502 231112 148508 231124
rect 77444 231084 148508 231112
rect 77444 231072 77450 231084
rect 148502 231072 148508 231084
rect 148560 231072 148566 231124
rect 158254 231072 158260 231124
rect 158312 231112 158318 231124
rect 167638 231112 167644 231124
rect 158312 231084 167644 231112
rect 158312 231072 158318 231084
rect 167638 231072 167644 231084
rect 167696 231072 167702 231124
rect 228726 231072 228732 231124
rect 228784 231112 228790 231124
rect 305178 231112 305184 231124
rect 228784 231084 305184 231112
rect 228784 231072 228790 231084
rect 305178 231072 305184 231084
rect 305236 231072 305242 231124
rect 187694 230500 187700 230512
rect 167012 230472 187700 230500
rect 63126 230392 63132 230444
rect 63184 230432 63190 230444
rect 167012 230432 167040 230472
rect 187694 230460 187700 230472
rect 187752 230460 187758 230512
rect 63184 230404 167040 230432
rect 63184 230392 63190 230404
rect 187234 230392 187240 230444
rect 187292 230432 187298 230444
rect 207658 230432 207664 230444
rect 187292 230404 207664 230432
rect 187292 230392 187298 230404
rect 207658 230392 207664 230404
rect 207716 230392 207722 230444
rect 142062 230324 142068 230376
rect 142120 230364 142126 230376
rect 234062 230364 234068 230376
rect 142120 230336 234068 230364
rect 142120 230324 142126 230336
rect 234062 230324 234068 230336
rect 234120 230324 234126 230376
rect 213178 229712 213184 229764
rect 213236 229752 213242 229764
rect 231946 229752 231952 229764
rect 213236 229724 231952 229752
rect 213236 229712 213242 229724
rect 231946 229712 231952 229724
rect 232004 229752 232010 229764
rect 287146 229752 287152 229764
rect 232004 229724 287152 229752
rect 232004 229712 232010 229724
rect 287146 229712 287152 229724
rect 287204 229712 287210 229764
rect 64782 229032 64788 229084
rect 64840 229072 64846 229084
rect 170490 229072 170496 229084
rect 64840 229044 170496 229072
rect 64840 229032 64846 229044
rect 170490 229032 170496 229044
rect 170548 229032 170554 229084
rect 202138 229032 202144 229084
rect 202196 229072 202202 229084
rect 252738 229072 252744 229084
rect 202196 229044 252744 229072
rect 202196 229032 202202 229044
rect 252738 229032 252744 229044
rect 252796 229032 252802 229084
rect 123018 228964 123024 229016
rect 123076 229004 123082 229016
rect 199378 229004 199384 229016
rect 123076 228976 199384 229004
rect 123076 228964 123082 228976
rect 199378 228964 199384 228976
rect 199436 228964 199442 229016
rect 173250 228896 173256 228948
rect 173308 228936 173314 228948
rect 220446 228936 220452 228948
rect 173308 228908 220452 228936
rect 173308 228896 173314 228908
rect 220446 228896 220452 228908
rect 220504 228896 220510 228948
rect 252738 228352 252744 228404
rect 252796 228392 252802 228404
rect 313366 228392 313372 228404
rect 252796 228364 313372 228392
rect 252796 228352 252802 228364
rect 313366 228352 313372 228364
rect 313424 228352 313430 228404
rect 220078 227740 220084 227792
rect 220136 227780 220142 227792
rect 220446 227780 220452 227792
rect 220136 227752 220452 227780
rect 220136 227740 220142 227752
rect 220446 227740 220452 227752
rect 220504 227740 220510 227792
rect 224218 227740 224224 227792
rect 224276 227780 224282 227792
rect 224276 227752 226380 227780
rect 224276 227740 224282 227752
rect 115750 227672 115756 227724
rect 115808 227712 115814 227724
rect 130378 227712 130384 227724
rect 115808 227684 130384 227712
rect 115808 227672 115814 227684
rect 130378 227672 130384 227684
rect 130436 227672 130442 227724
rect 226352 227712 226380 227752
rect 227254 227740 227260 227792
rect 227312 227780 227318 227792
rect 227806 227780 227812 227792
rect 227312 227752 227812 227780
rect 227312 227740 227318 227752
rect 227806 227740 227812 227752
rect 227864 227780 227870 227792
rect 284386 227780 284392 227792
rect 227864 227752 284392 227780
rect 227864 227740 227870 227752
rect 284386 227740 284392 227752
rect 284444 227740 284450 227792
rect 229738 227712 229744 227724
rect 226352 227684 229744 227712
rect 229738 227672 229744 227684
rect 229796 227672 229802 227724
rect 135162 227060 135168 227112
rect 135220 227100 135226 227112
rect 146754 227100 146760 227112
rect 135220 227072 146760 227100
rect 135220 227060 135226 227072
rect 146754 227060 146760 227072
rect 146812 227060 146818 227112
rect 148502 227060 148508 227112
rect 148560 227100 148566 227112
rect 215938 227100 215944 227112
rect 148560 227072 215944 227100
rect 148560 227060 148566 227072
rect 215938 227060 215944 227072
rect 215996 227060 216002 227112
rect 217134 227060 217140 227112
rect 217192 227100 217198 227112
rect 226334 227100 226340 227112
rect 217192 227072 226340 227100
rect 217192 227060 217198 227072
rect 226334 227060 226340 227072
rect 226392 227060 226398 227112
rect 56318 226992 56324 227044
rect 56376 227032 56382 227044
rect 115198 227032 115204 227044
rect 56376 227004 115204 227032
rect 56376 226992 56382 227004
rect 115198 226992 115204 227004
rect 115256 226992 115262 227044
rect 119430 226992 119436 227044
rect 119488 227032 119494 227044
rect 194962 227032 194968 227044
rect 119488 227004 194968 227032
rect 119488 226992 119494 227004
rect 194962 226992 194968 227004
rect 195020 226992 195026 227044
rect 214098 226992 214104 227044
rect 214156 227032 214162 227044
rect 225598 227032 225604 227044
rect 214156 227004 225604 227032
rect 214156 226992 214162 227004
rect 225598 226992 225604 227004
rect 225656 226992 225662 227044
rect 282178 226992 282184 227044
rect 282236 227032 282242 227044
rect 292666 227032 292672 227044
rect 282236 227004 292672 227032
rect 282236 226992 282242 227004
rect 292666 226992 292672 227004
rect 292724 226992 292730 227044
rect 236822 226352 236828 226364
rect 236012 226324 236828 226352
rect 86218 226244 86224 226296
rect 86276 226284 86282 226296
rect 137370 226284 137376 226296
rect 86276 226256 137376 226284
rect 86276 226244 86282 226256
rect 137370 226244 137376 226256
rect 137428 226244 137434 226296
rect 144730 226244 144736 226296
rect 144788 226284 144794 226296
rect 236012 226284 236040 226324
rect 236822 226312 236828 226324
rect 236880 226352 236886 226364
rect 313274 226352 313280 226364
rect 236880 226324 313280 226352
rect 236880 226312 236886 226324
rect 313274 226312 313280 226324
rect 313332 226312 313338 226364
rect 144788 226256 236040 226284
rect 144788 226244 144794 226256
rect 57790 225564 57796 225616
rect 57848 225604 57854 225616
rect 142890 225604 142896 225616
rect 57848 225576 142896 225604
rect 57848 225564 57854 225576
rect 142890 225564 142896 225576
rect 142948 225564 142954 225616
rect 143350 225564 143356 225616
rect 143408 225604 143414 225616
rect 230382 225604 230388 225616
rect 143408 225576 230388 225604
rect 143408 225564 143414 225576
rect 230382 225564 230388 225576
rect 230440 225604 230446 225616
rect 231118 225604 231124 225616
rect 230440 225576 231124 225604
rect 230440 225564 230446 225576
rect 231118 225564 231124 225576
rect 231176 225564 231182 225616
rect 238294 225564 238300 225616
rect 238352 225604 238358 225616
rect 245838 225604 245844 225616
rect 238352 225576 245844 225604
rect 238352 225564 238358 225576
rect 245838 225564 245844 225576
rect 245896 225564 245902 225616
rect 76650 224884 76656 224936
rect 76708 224924 76714 224936
rect 244274 224924 244280 224936
rect 76708 224896 244280 224924
rect 76708 224884 76714 224896
rect 244274 224884 244280 224896
rect 244332 224884 244338 224936
rect 132310 224204 132316 224256
rect 132368 224244 132374 224256
rect 164878 224244 164884 224256
rect 132368 224216 164884 224244
rect 132368 224204 132374 224216
rect 164878 224204 164884 224216
rect 164936 224204 164942 224256
rect 193030 223592 193036 223644
rect 193088 223632 193094 223644
rect 582466 223632 582472 223644
rect 193088 223604 582472 223632
rect 193088 223592 193094 223604
rect 582466 223592 582472 223604
rect 582524 223592 582530 223644
rect 160002 223524 160008 223576
rect 160060 223564 160066 223576
rect 160922 223564 160928 223576
rect 160060 223536 160928 223564
rect 160060 223524 160066 223536
rect 160922 223524 160928 223536
rect 160980 223524 160986 223576
rect 188062 223524 188068 223576
rect 188120 223564 188126 223576
rect 188798 223564 188804 223576
rect 188120 223536 188804 223564
rect 188120 223524 188126 223536
rect 188798 223524 188804 223536
rect 188856 223564 188862 223576
rect 191098 223564 191104 223576
rect 188856 223536 191104 223564
rect 188856 223524 188862 223536
rect 191098 223524 191104 223536
rect 191156 223524 191162 223576
rect 194962 223524 194968 223576
rect 195020 223564 195026 223576
rect 217502 223564 217508 223576
rect 195020 223536 217508 223564
rect 195020 223524 195026 223536
rect 217502 223524 217508 223536
rect 217560 223524 217566 223576
rect 136542 222912 136548 222964
rect 136600 222952 136606 222964
rect 160002 222952 160008 222964
rect 136600 222924 160008 222952
rect 136600 222912 136606 222924
rect 160002 222912 160008 222924
rect 160060 222912 160066 222964
rect 162210 222912 162216 222964
rect 162268 222952 162274 222964
rect 199470 222952 199476 222964
rect 162268 222924 199476 222952
rect 162268 222912 162274 222924
rect 199470 222912 199476 222924
rect 199528 222912 199534 222964
rect 86954 222844 86960 222896
rect 87012 222884 87018 222896
rect 188062 222884 188068 222896
rect 87012 222856 188068 222884
rect 87012 222844 87018 222856
rect 188062 222844 188068 222856
rect 188120 222844 188126 222896
rect 204990 222844 204996 222896
rect 205048 222884 205054 222896
rect 582742 222884 582748 222896
rect 205048 222856 582748 222884
rect 205048 222844 205054 222856
rect 582742 222844 582748 222856
rect 582800 222844 582806 222896
rect 187694 222096 187700 222148
rect 187752 222136 187758 222148
rect 193030 222136 193036 222148
rect 187752 222108 193036 222136
rect 187752 222096 187758 222108
rect 193030 222096 193036 222108
rect 193088 222096 193094 222148
rect 50522 222028 50528 222080
rect 50580 222068 50586 222080
rect 50798 222068 50804 222080
rect 50580 222040 50804 222068
rect 50580 222028 50586 222040
rect 50798 222028 50804 222040
rect 50856 222068 50862 222080
rect 93854 222068 93860 222080
rect 50856 222040 93860 222068
rect 50856 222028 50862 222040
rect 93854 222028 93860 222040
rect 93912 222028 93918 222080
rect 99466 222028 99472 222080
rect 99524 222068 99530 222080
rect 211246 222068 211252 222080
rect 99524 222040 211252 222068
rect 99524 222028 99530 222040
rect 211246 222028 211252 222040
rect 211304 222068 211310 222080
rect 211798 222068 211804 222080
rect 211304 222040 211804 222068
rect 211304 222028 211310 222040
rect 211798 222028 211804 222040
rect 211856 222028 211862 222080
rect 57606 221960 57612 222012
rect 57664 222000 57670 222012
rect 188430 222000 188436 222012
rect 57664 221972 188436 222000
rect 57664 221960 57670 221972
rect 188430 221960 188436 221972
rect 188488 221960 188494 222012
rect 215938 221484 215944 221536
rect 215996 221524 216002 221536
rect 246298 221524 246304 221536
rect 215996 221496 246304 221524
rect 215996 221484 216002 221496
rect 246298 221484 246304 221496
rect 246356 221484 246362 221536
rect 4798 221416 4804 221468
rect 4856 221456 4862 221468
rect 50522 221456 50528 221468
rect 4856 221428 50528 221456
rect 4856 221416 4862 221428
rect 50522 221416 50528 221428
rect 50580 221416 50586 221468
rect 197078 221416 197084 221468
rect 197136 221456 197142 221468
rect 255406 221456 255412 221468
rect 197136 221428 255412 221456
rect 197136 221416 197142 221428
rect 255406 221416 255412 221428
rect 255464 221416 255470 221468
rect 580902 220940 580908 220992
rect 580960 220980 580966 220992
rect 583202 220980 583208 220992
rect 580960 220952 583208 220980
rect 580960 220940 580966 220952
rect 583202 220940 583208 220952
rect 583260 220940 583266 220992
rect 144822 220736 144828 220788
rect 144880 220776 144886 220788
rect 235258 220776 235264 220788
rect 144880 220748 235264 220776
rect 144880 220736 144886 220748
rect 235258 220736 235264 220748
rect 235316 220736 235322 220788
rect 193030 220668 193036 220720
rect 193088 220708 193094 220720
rect 193950 220708 193956 220720
rect 193088 220680 193956 220708
rect 193088 220668 193094 220680
rect 193950 220668 193956 220680
rect 194008 220668 194014 220720
rect 104986 220056 104992 220108
rect 105044 220096 105050 220108
rect 193030 220096 193036 220108
rect 105044 220068 193036 220096
rect 105044 220056 105050 220068
rect 193030 220056 193036 220068
rect 193088 220056 193094 220108
rect 201494 220056 201500 220108
rect 201552 220096 201558 220108
rect 301038 220096 301044 220108
rect 201552 220068 301044 220096
rect 201552 220056 201558 220068
rect 301038 220056 301044 220068
rect 301096 220056 301102 220108
rect 155402 219376 155408 219428
rect 155460 219416 155466 219428
rect 242894 219416 242900 219428
rect 155460 219388 242900 219416
rect 155460 219376 155466 219388
rect 242894 219376 242900 219388
rect 242952 219376 242958 219428
rect 304258 219376 304264 219428
rect 304316 219416 304322 219428
rect 580166 219416 580172 219428
rect 304316 219388 580172 219416
rect 304316 219376 304322 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 137922 219308 137928 219360
rect 137980 219348 137986 219360
rect 213178 219348 213184 219360
rect 137980 219320 213184 219348
rect 137980 219308 137986 219320
rect 213178 219308 213184 219320
rect 213236 219308 213242 219360
rect 242894 218764 242900 218816
rect 242952 218804 242958 218816
rect 243906 218804 243912 218816
rect 242952 218776 243912 218804
rect 242952 218764 242958 218776
rect 243906 218764 243912 218776
rect 243964 218764 243970 218816
rect 52178 218696 52184 218748
rect 52236 218736 52242 218748
rect 143350 218736 143356 218748
rect 52236 218708 143356 218736
rect 52236 218696 52242 218708
rect 143350 218696 143356 218708
rect 143408 218696 143414 218748
rect 67726 217948 67732 218000
rect 67784 217988 67790 218000
rect 137462 217988 137468 218000
rect 67784 217960 137468 217988
rect 67784 217948 67790 217960
rect 137462 217948 137468 217960
rect 137520 217948 137526 218000
rect 130930 217880 130936 217932
rect 130988 217920 130994 217932
rect 181530 217920 181536 217932
rect 130988 217892 181536 217920
rect 130988 217880 130994 217892
rect 181530 217880 181536 217892
rect 181588 217880 181594 217932
rect 189074 217336 189080 217388
rect 189132 217376 189138 217388
rect 231854 217376 231860 217388
rect 189132 217348 231860 217376
rect 189132 217336 189138 217348
rect 231854 217336 231860 217348
rect 231912 217336 231918 217388
rect 142890 217268 142896 217320
rect 142948 217308 142954 217320
rect 218054 217308 218060 217320
rect 142948 217280 218060 217308
rect 142948 217268 142954 217280
rect 218054 217268 218060 217280
rect 218112 217268 218118 217320
rect 218974 217268 218980 217320
rect 219032 217308 219038 217320
rect 219434 217308 219440 217320
rect 219032 217280 219440 217308
rect 219032 217268 219038 217280
rect 219434 217268 219440 217280
rect 219492 217268 219498 217320
rect 220262 217268 220268 217320
rect 220320 217308 220326 217320
rect 291378 217308 291384 217320
rect 220320 217280 291384 217308
rect 220320 217268 220326 217280
rect 291378 217268 291384 217280
rect 291436 217268 291442 217320
rect 81618 216588 81624 216640
rect 81676 216628 81682 216640
rect 191282 216628 191288 216640
rect 81676 216600 191288 216628
rect 81676 216588 81682 216600
rect 191282 216588 191288 216600
rect 191340 216588 191346 216640
rect 180058 216520 180064 216572
rect 180116 216560 180122 216572
rect 255498 216560 255504 216572
rect 180116 216532 255504 216560
rect 180116 216520 180122 216532
rect 255498 216520 255504 216532
rect 255556 216520 255562 216572
rect 100662 215908 100668 215960
rect 100720 215948 100726 215960
rect 173158 215948 173164 215960
rect 100720 215920 173164 215948
rect 100720 215908 100726 215920
rect 173158 215908 173164 215920
rect 173216 215908 173222 215960
rect 193950 215908 193956 215960
rect 194008 215948 194014 215960
rect 207382 215948 207388 215960
rect 194008 215920 207388 215948
rect 194008 215908 194014 215920
rect 207382 215908 207388 215920
rect 207440 215908 207446 215960
rect 298738 215908 298744 215960
rect 298796 215948 298802 215960
rect 309318 215948 309324 215960
rect 298796 215920 309324 215948
rect 298796 215908 298802 215920
rect 309318 215908 309324 215920
rect 309376 215908 309382 215960
rect 255498 215296 255504 215348
rect 255556 215336 255562 215348
rect 255958 215336 255964 215348
rect 255556 215308 255964 215336
rect 255556 215296 255562 215308
rect 255958 215296 255964 215308
rect 256016 215296 256022 215348
rect 3326 215228 3332 215280
rect 3384 215268 3390 215280
rect 40678 215268 40684 215280
rect 3384 215240 40684 215268
rect 3384 215228 3390 215240
rect 40678 215228 40684 215240
rect 40736 215228 40742 215280
rect 199378 214616 199384 214668
rect 199436 214656 199442 214668
rect 230566 214656 230572 214668
rect 199436 214628 230572 214656
rect 199436 214616 199442 214628
rect 230566 214616 230572 214628
rect 230624 214616 230630 214668
rect 61746 214548 61752 214600
rect 61804 214588 61810 214600
rect 115290 214588 115296 214600
rect 61804 214560 115296 214588
rect 61804 214548 61810 214560
rect 115290 214548 115296 214560
rect 115348 214548 115354 214600
rect 126882 214548 126888 214600
rect 126940 214588 126946 214600
rect 197354 214588 197360 214600
rect 126940 214560 197360 214588
rect 126940 214548 126946 214560
rect 197354 214548 197360 214560
rect 197412 214548 197418 214600
rect 203334 214548 203340 214600
rect 203392 214588 203398 214600
rect 211154 214588 211160 214600
rect 203392 214560 211160 214588
rect 203392 214548 203398 214560
rect 211154 214548 211160 214560
rect 211212 214588 211218 214600
rect 307938 214588 307944 214600
rect 211212 214560 307944 214588
rect 211212 214548 211218 214560
rect 307938 214548 307944 214560
rect 307996 214548 308002 214600
rect 167638 213936 167644 213988
rect 167696 213976 167702 213988
rect 202966 213976 202972 213988
rect 167696 213948 202972 213976
rect 167696 213936 167702 213948
rect 202966 213936 202972 213948
rect 203024 213976 203030 213988
rect 203610 213976 203616 213988
rect 203024 213948 203616 213976
rect 203024 213936 203030 213948
rect 203610 213936 203616 213948
rect 203668 213936 203674 213988
rect 75178 213868 75184 213920
rect 75236 213908 75242 213920
rect 195330 213908 195336 213920
rect 75236 213880 195336 213908
rect 75236 213868 75242 213880
rect 195330 213868 195336 213880
rect 195388 213868 195394 213920
rect 197354 213868 197360 213920
rect 197412 213908 197418 213920
rect 227806 213908 227812 213920
rect 197412 213880 227812 213908
rect 197412 213868 197418 213880
rect 227806 213868 227812 213880
rect 227864 213868 227870 213920
rect 133874 213800 133880 213852
rect 133932 213840 133938 213852
rect 244366 213840 244372 213852
rect 133932 213812 244372 213840
rect 133932 213800 133938 213812
rect 244366 213800 244372 213812
rect 244424 213800 244430 213852
rect 240962 213188 240968 213240
rect 241020 213228 241026 213240
rect 285766 213228 285772 213240
rect 241020 213200 285772 213228
rect 241020 213188 241026 213200
rect 285766 213188 285772 213200
rect 285824 213188 285830 213240
rect 71038 212440 71044 212492
rect 71096 212480 71102 212492
rect 233510 212480 233516 212492
rect 71096 212452 233516 212480
rect 71096 212440 71102 212452
rect 233510 212440 233516 212452
rect 233568 212480 233574 212492
rect 234430 212480 234436 212492
rect 233568 212452 234436 212480
rect 233568 212440 233574 212452
rect 234430 212440 234436 212452
rect 234488 212440 234494 212492
rect 146202 212372 146208 212424
rect 146260 212412 146266 212424
rect 244550 212412 244556 212424
rect 146260 212384 244556 212412
rect 146260 212372 146266 212384
rect 244550 212372 244556 212384
rect 244608 212372 244614 212424
rect 69014 211080 69020 211132
rect 69072 211120 69078 211132
rect 189074 211120 189080 211132
rect 69072 211092 189080 211120
rect 69072 211080 69078 211092
rect 189074 211080 189080 211092
rect 189132 211080 189138 211132
rect 162302 211012 162308 211064
rect 162360 211052 162366 211064
rect 256786 211052 256792 211064
rect 162360 211024 256792 211052
rect 162360 211012 162366 211024
rect 256786 211012 256792 211024
rect 256844 211012 256850 211064
rect 197906 209788 197912 209840
rect 197964 209828 197970 209840
rect 214466 209828 214472 209840
rect 197964 209800 214472 209828
rect 197964 209788 197970 209800
rect 214466 209788 214472 209800
rect 214524 209828 214530 209840
rect 239398 209828 239404 209840
rect 214524 209800 239404 209828
rect 214524 209788 214530 209800
rect 239398 209788 239404 209800
rect 239456 209788 239462 209840
rect 103422 209108 103428 209160
rect 103480 209148 103486 209160
rect 133138 209148 133144 209160
rect 103480 209120 133144 209148
rect 103480 209108 103486 209120
rect 133138 209108 133144 209120
rect 133196 209108 133202 209160
rect 133690 209108 133696 209160
rect 133748 209148 133754 209160
rect 193858 209148 193864 209160
rect 133748 209120 193864 209148
rect 133748 209108 133754 209120
rect 193858 209108 193864 209120
rect 193916 209108 193922 209160
rect 204898 209108 204904 209160
rect 204956 209148 204962 209160
rect 302510 209148 302516 209160
rect 204956 209120 302516 209148
rect 204956 209108 204962 209120
rect 302510 209108 302516 209120
rect 302568 209108 302574 209160
rect 67634 209040 67640 209092
rect 67692 209080 67698 209092
rect 205542 209080 205548 209092
rect 67692 209052 205548 209080
rect 67692 209040 67698 209052
rect 205542 209040 205548 209052
rect 205600 209040 205606 209092
rect 236638 209040 236644 209092
rect 236696 209080 236702 209092
rect 298738 209080 298744 209092
rect 236696 209052 298744 209080
rect 236696 209040 236702 209052
rect 298738 209040 298744 209052
rect 298796 209040 298802 209092
rect 205542 208836 205548 208888
rect 205600 208876 205606 208888
rect 206462 208876 206468 208888
rect 205600 208848 206468 208876
rect 205600 208836 205606 208848
rect 206462 208836 206468 208848
rect 206520 208836 206526 208888
rect 85574 208292 85580 208344
rect 85632 208332 85638 208344
rect 197906 208332 197912 208344
rect 85632 208304 197912 208332
rect 85632 208292 85638 208304
rect 197906 208292 197912 208304
rect 197964 208292 197970 208344
rect 200022 207680 200028 207732
rect 200080 207720 200086 207732
rect 230474 207720 230480 207732
rect 200080 207692 230480 207720
rect 200080 207680 200086 207692
rect 230474 207680 230480 207692
rect 230532 207680 230538 207732
rect 235258 207680 235264 207732
rect 235316 207720 235322 207732
rect 294138 207720 294144 207732
rect 235316 207692 294144 207720
rect 235316 207680 235322 207692
rect 294138 207680 294144 207692
rect 294196 207680 294202 207732
rect 113082 207612 113088 207664
rect 113140 207652 113146 207664
rect 236270 207652 236276 207664
rect 113140 207624 236276 207652
rect 113140 207612 113146 207624
rect 236270 207612 236276 207624
rect 236328 207652 236334 207664
rect 248690 207652 248696 207664
rect 236328 207624 248696 207652
rect 236328 207612 236334 207624
rect 248690 207612 248696 207624
rect 248748 207612 248754 207664
rect 93118 206932 93124 206984
rect 93176 206972 93182 206984
rect 208302 206972 208308 206984
rect 93176 206944 208308 206972
rect 93176 206932 93182 206944
rect 208302 206932 208308 206944
rect 208360 206932 208366 206984
rect 110230 206864 110236 206916
rect 110288 206904 110294 206916
rect 219434 206904 219440 206916
rect 110288 206876 219440 206904
rect 110288 206864 110294 206876
rect 219434 206864 219440 206876
rect 219492 206904 219498 206916
rect 220722 206904 220728 206916
rect 219492 206876 220728 206904
rect 219492 206864 219498 206876
rect 220722 206864 220728 206876
rect 220780 206864 220786 206916
rect 220722 206252 220728 206304
rect 220780 206292 220786 206304
rect 280246 206292 280252 206304
rect 220780 206264 280252 206292
rect 220780 206252 220786 206264
rect 280246 206252 280252 206264
rect 280304 206252 280310 206304
rect 207842 206116 207848 206168
rect 207900 206156 207906 206168
rect 208302 206156 208308 206168
rect 207900 206128 208308 206156
rect 207900 206116 207906 206128
rect 208302 206116 208308 206128
rect 208360 206116 208366 206168
rect 81342 205572 81348 205624
rect 81400 205612 81406 205624
rect 157334 205612 157340 205624
rect 81400 205584 157340 205612
rect 81400 205572 81406 205584
rect 157334 205572 157340 205584
rect 157392 205572 157398 205624
rect 164878 205572 164884 205624
rect 164936 205612 164942 205624
rect 240134 205612 240140 205624
rect 164936 205584 240140 205612
rect 164936 205572 164942 205584
rect 240134 205572 240140 205584
rect 240192 205612 240198 205624
rect 240870 205612 240876 205624
rect 240192 205584 240876 205612
rect 240192 205572 240198 205584
rect 240870 205572 240876 205584
rect 240928 205572 240934 205624
rect 95234 204892 95240 204944
rect 95292 204932 95298 204944
rect 242986 204932 242992 204944
rect 95292 204904 242992 204932
rect 95292 204892 95298 204904
rect 242986 204892 242992 204904
rect 243044 204892 243050 204944
rect 70394 204212 70400 204264
rect 70452 204252 70458 204264
rect 215478 204252 215484 204264
rect 70452 204224 215484 204252
rect 70452 204212 70458 204224
rect 215478 204212 215484 204224
rect 215536 204212 215542 204264
rect 74534 204144 74540 204196
rect 74592 204184 74598 204196
rect 167638 204184 167644 204196
rect 74592 204156 167644 204184
rect 74592 204144 74598 204156
rect 167638 204144 167644 204156
rect 167696 204144 167702 204196
rect 215478 203600 215484 203652
rect 215536 203640 215542 203652
rect 228542 203640 228548 203652
rect 215536 203612 228548 203640
rect 215536 203600 215542 203612
rect 228542 203600 228548 203612
rect 228600 203600 228606 203652
rect 262858 203600 262864 203652
rect 262916 203640 262922 203652
rect 306650 203640 306656 203652
rect 262916 203612 306656 203640
rect 262916 203600 262922 203612
rect 306650 203600 306656 203612
rect 306708 203600 306714 203652
rect 173158 203532 173164 203584
rect 173216 203572 173222 203584
rect 195422 203572 195428 203584
rect 173216 203544 195428 203572
rect 173216 203532 173222 203544
rect 195422 203532 195428 203544
rect 195480 203532 195486 203584
rect 225598 203532 225604 203584
rect 225656 203572 225662 203584
rect 291286 203572 291292 203584
rect 225656 203544 291292 203572
rect 225656 203532 225662 203544
rect 291286 203532 291292 203544
rect 291344 203532 291350 203584
rect 3418 202784 3424 202836
rect 3476 202824 3482 202836
rect 119430 202824 119436 202836
rect 3476 202796 119436 202824
rect 3476 202784 3482 202796
rect 119430 202784 119436 202796
rect 119488 202784 119494 202836
rect 121362 202784 121368 202836
rect 121420 202824 121426 202836
rect 155218 202824 155224 202836
rect 121420 202796 155224 202824
rect 121420 202784 121426 202796
rect 155218 202784 155224 202796
rect 155276 202784 155282 202836
rect 171778 202172 171784 202224
rect 171836 202212 171842 202224
rect 186958 202212 186964 202224
rect 171836 202184 186964 202212
rect 171836 202172 171842 202184
rect 186958 202172 186964 202184
rect 187016 202172 187022 202224
rect 193122 202172 193128 202224
rect 193180 202212 193186 202224
rect 252646 202212 252652 202224
rect 193180 202184 252652 202212
rect 193180 202172 193186 202184
rect 252646 202172 252652 202184
rect 252704 202172 252710 202224
rect 125502 202104 125508 202156
rect 125560 202144 125566 202156
rect 237374 202144 237380 202156
rect 125560 202116 237380 202144
rect 125560 202104 125566 202116
rect 237374 202104 237380 202116
rect 237432 202144 237438 202156
rect 247126 202144 247132 202156
rect 237432 202116 247132 202144
rect 237432 202104 237438 202116
rect 247126 202104 247132 202116
rect 247184 202104 247190 202156
rect 264238 202104 264244 202156
rect 264296 202144 264302 202156
rect 310606 202144 310612 202156
rect 264296 202116 310612 202144
rect 264296 202104 264302 202116
rect 310606 202104 310612 202116
rect 310664 202104 310670 202156
rect 63310 201424 63316 201476
rect 63368 201464 63374 201476
rect 214650 201464 214656 201476
rect 63368 201436 214656 201464
rect 63368 201424 63374 201436
rect 214650 201424 214656 201436
rect 214708 201424 214714 201476
rect 223022 200812 223028 200864
rect 223080 200852 223086 200864
rect 229094 200852 229100 200864
rect 223080 200824 229100 200852
rect 223080 200812 223086 200824
rect 229094 200812 229100 200824
rect 229152 200812 229158 200864
rect 214926 200200 214932 200252
rect 214984 200240 214990 200252
rect 225690 200240 225696 200252
rect 214984 200212 225696 200240
rect 214984 200200 214990 200212
rect 225690 200200 225696 200212
rect 225748 200200 225754 200252
rect 186130 200132 186136 200184
rect 186188 200172 186194 200184
rect 247678 200172 247684 200184
rect 186188 200144 247684 200172
rect 186188 200132 186194 200144
rect 247678 200132 247684 200144
rect 247736 200132 247742 200184
rect 46842 200064 46848 200116
rect 46900 200104 46906 200116
rect 217410 200104 217416 200116
rect 46900 200076 217416 200104
rect 46900 200064 46906 200076
rect 217410 200064 217416 200076
rect 217468 200064 217474 200116
rect 131022 199996 131028 200048
rect 131080 200036 131086 200048
rect 187050 200036 187056 200048
rect 131080 200008 187056 200036
rect 131080 199996 131086 200008
rect 187050 199996 187056 200008
rect 187108 199996 187114 200048
rect 222102 198772 222108 198824
rect 222160 198812 222166 198824
rect 238110 198812 238116 198824
rect 222160 198784 238116 198812
rect 222160 198772 222166 198784
rect 238110 198772 238116 198784
rect 238168 198772 238174 198824
rect 296898 198744 296904 198756
rect 187620 198716 296904 198744
rect 187620 198688 187648 198716
rect 296898 198704 296904 198716
rect 296956 198704 296962 198756
rect 110322 198636 110328 198688
rect 110380 198676 110386 198688
rect 187602 198676 187608 198688
rect 110380 198648 187608 198676
rect 110380 198636 110386 198648
rect 187602 198636 187608 198648
rect 187660 198636 187666 198688
rect 192570 198636 192576 198688
rect 192628 198676 192634 198688
rect 222102 198676 222108 198688
rect 192628 198648 222108 198676
rect 192628 198636 192634 198648
rect 222102 198636 222108 198648
rect 222160 198636 222166 198688
rect 58894 197956 58900 198008
rect 58952 197996 58958 198008
rect 133782 197996 133788 198008
rect 58952 197968 133788 197996
rect 58952 197956 58958 197968
rect 133782 197956 133788 197968
rect 133840 197956 133846 198008
rect 202230 197956 202236 198008
rect 202288 197996 202294 198008
rect 286318 197996 286324 198008
rect 202288 197968 286324 197996
rect 202288 197956 202294 197968
rect 286318 197956 286324 197968
rect 286376 197956 286382 198008
rect 133782 197276 133788 197328
rect 133840 197316 133846 197328
rect 186130 197316 186136 197328
rect 133840 197288 186136 197316
rect 133840 197276 133846 197288
rect 186130 197276 186136 197288
rect 186188 197276 186194 197328
rect 207842 197276 207848 197328
rect 207900 197316 207906 197328
rect 214926 197316 214932 197328
rect 207900 197288 214932 197316
rect 207900 197276 207906 197288
rect 214926 197276 214932 197288
rect 214984 197276 214990 197328
rect 195238 196664 195244 196716
rect 195296 196704 195302 196716
rect 227070 196704 227076 196716
rect 195296 196676 227076 196704
rect 195296 196664 195302 196676
rect 227070 196664 227076 196676
rect 227128 196664 227134 196716
rect 228358 196664 228364 196716
rect 228416 196704 228422 196716
rect 303798 196704 303804 196716
rect 228416 196676 303804 196704
rect 228416 196664 228422 196676
rect 303798 196664 303804 196676
rect 303856 196664 303862 196716
rect 89530 196596 89536 196648
rect 89588 196636 89594 196648
rect 196894 196636 196900 196648
rect 89588 196608 196900 196636
rect 89588 196596 89594 196608
rect 196894 196596 196900 196608
rect 196952 196596 196958 196648
rect 214558 196596 214564 196648
rect 214616 196636 214622 196648
rect 295610 196636 295616 196648
rect 214616 196608 295616 196636
rect 214616 196596 214622 196608
rect 295610 196596 295616 196608
rect 295668 196596 295674 196648
rect 56410 195916 56416 195968
rect 56468 195956 56474 195968
rect 174630 195956 174636 195968
rect 56468 195928 174636 195956
rect 56468 195916 56474 195928
rect 174630 195916 174636 195928
rect 174688 195916 174694 195968
rect 79962 195848 79968 195900
rect 80020 195888 80026 195900
rect 189258 195888 189264 195900
rect 80020 195860 189264 195888
rect 80020 195848 80026 195860
rect 189258 195848 189264 195860
rect 189316 195848 189322 195900
rect 189258 195304 189264 195356
rect 189316 195344 189322 195356
rect 190362 195344 190368 195356
rect 189316 195316 190368 195344
rect 189316 195304 189322 195316
rect 190362 195304 190368 195316
rect 190420 195344 190426 195356
rect 228358 195344 228364 195356
rect 190420 195316 228364 195344
rect 190420 195304 190426 195316
rect 228358 195304 228364 195316
rect 228416 195304 228422 195356
rect 203610 195236 203616 195288
rect 203668 195276 203674 195288
rect 279050 195276 279056 195288
rect 203668 195248 279056 195276
rect 203668 195236 203674 195248
rect 279050 195236 279056 195248
rect 279108 195236 279114 195288
rect 316678 195236 316684 195288
rect 316736 195276 316742 195288
rect 325694 195276 325700 195288
rect 316736 195248 325700 195276
rect 316736 195236 316742 195248
rect 325694 195236 325700 195248
rect 325752 195236 325758 195288
rect 86862 194488 86868 194540
rect 86920 194528 86926 194540
rect 168374 194528 168380 194540
rect 86920 194500 168380 194528
rect 86920 194488 86926 194500
rect 168374 194488 168380 194500
rect 168432 194488 168438 194540
rect 188890 193876 188896 193928
rect 188948 193916 188954 193928
rect 251818 193916 251824 193928
rect 188948 193888 251824 193916
rect 188948 193876 188954 193888
rect 251818 193876 251824 193888
rect 251876 193876 251882 193928
rect 255958 193876 255964 193928
rect 256016 193916 256022 193928
rect 268470 193916 268476 193928
rect 256016 193888 268476 193916
rect 256016 193876 256022 193888
rect 268470 193876 268476 193888
rect 268528 193876 268534 193928
rect 177942 193808 177948 193860
rect 178000 193848 178006 193860
rect 302326 193848 302332 193860
rect 178000 193820 302332 193848
rect 178000 193808 178006 193820
rect 302326 193808 302332 193820
rect 302384 193808 302390 193860
rect 115198 193128 115204 193180
rect 115256 193168 115262 193180
rect 197998 193168 198004 193180
rect 115256 193140 198004 193168
rect 115256 193128 115262 193140
rect 197998 193128 198004 193140
rect 198056 193128 198062 193180
rect 197262 192516 197268 192568
rect 197320 192556 197326 192568
rect 228450 192556 228456 192568
rect 197320 192528 228456 192556
rect 197320 192516 197326 192528
rect 228450 192516 228456 192528
rect 228508 192516 228514 192568
rect 228634 192516 228640 192568
rect 228692 192556 228698 192568
rect 235350 192556 235356 192568
rect 228692 192528 235356 192556
rect 228692 192516 228698 192528
rect 235350 192516 235356 192528
rect 235408 192516 235414 192568
rect 268378 192516 268384 192568
rect 268436 192556 268442 192568
rect 296806 192556 296812 192568
rect 268436 192528 296812 192556
rect 268436 192516 268442 192528
rect 296806 192516 296812 192528
rect 296864 192516 296870 192568
rect 202782 192448 202788 192500
rect 202840 192488 202846 192500
rect 305270 192488 305276 192500
rect 202840 192460 305276 192488
rect 202840 192448 202846 192460
rect 305270 192448 305276 192460
rect 305328 192448 305334 192500
rect 143442 191768 143448 191820
rect 143500 191808 143506 191820
rect 209222 191808 209228 191820
rect 143500 191780 209228 191808
rect 143500 191768 143506 191780
rect 209222 191768 209228 191780
rect 209280 191768 209286 191820
rect 179322 191700 179328 191752
rect 179380 191740 179386 191752
rect 180242 191740 180248 191752
rect 179380 191712 180248 191740
rect 179380 191700 179386 191712
rect 180242 191700 180248 191712
rect 180300 191700 180306 191752
rect 191282 191156 191288 191208
rect 191340 191196 191346 191208
rect 233970 191196 233976 191208
rect 191340 191168 233976 191196
rect 191340 191156 191346 191168
rect 233970 191156 233976 191168
rect 234028 191156 234034 191208
rect 104894 191088 104900 191140
rect 104952 191128 104958 191140
rect 179322 191128 179328 191140
rect 104952 191100 179328 191128
rect 104952 191088 104958 191100
rect 179322 191088 179328 191100
rect 179380 191088 179386 191140
rect 209038 191088 209044 191140
rect 209096 191128 209102 191140
rect 281810 191128 281816 191140
rect 209096 191100 281816 191128
rect 209096 191088 209102 191100
rect 281810 191088 281816 191100
rect 281868 191088 281874 191140
rect 69658 190408 69664 190460
rect 69716 190448 69722 190460
rect 193950 190448 193956 190460
rect 69716 190420 193956 190448
rect 69716 190408 69722 190420
rect 193950 190408 193956 190420
rect 194008 190408 194014 190460
rect 228542 189796 228548 189848
rect 228600 189836 228606 189848
rect 244458 189836 244464 189848
rect 228600 189808 244464 189836
rect 228600 189796 228606 189808
rect 244458 189796 244464 189808
rect 244516 189796 244522 189848
rect 188982 189728 188988 189780
rect 189040 189768 189046 189780
rect 231946 189768 231952 189780
rect 189040 189740 231952 189768
rect 189040 189728 189046 189740
rect 231946 189728 231952 189740
rect 232004 189728 232010 189780
rect 129642 189048 129648 189100
rect 129700 189088 129706 189100
rect 166258 189088 166264 189100
rect 129700 189060 166264 189088
rect 129700 189048 129706 189060
rect 166258 189048 166264 189060
rect 166316 189048 166322 189100
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 35250 189020 35256 189032
rect 3568 188992 35256 189020
rect 3568 188980 3574 188992
rect 35250 188980 35256 188992
rect 35308 188980 35314 189032
rect 187050 188368 187056 188420
rect 187108 188408 187114 188420
rect 221366 188408 221372 188420
rect 187108 188380 221372 188408
rect 187108 188368 187114 188380
rect 221366 188368 221372 188380
rect 221424 188368 221430 188420
rect 35158 188300 35164 188352
rect 35216 188340 35222 188352
rect 162118 188340 162124 188352
rect 35216 188312 162124 188340
rect 35216 188300 35222 188312
rect 162118 188300 162124 188312
rect 162176 188300 162182 188352
rect 174630 188300 174636 188352
rect 174688 188340 174694 188352
rect 288618 188340 288624 188352
rect 174688 188312 288624 188340
rect 174688 188300 174694 188312
rect 288618 188300 288624 188312
rect 288676 188300 288682 188352
rect 135162 187688 135168 187740
rect 135220 187728 135226 187740
rect 163498 187728 163504 187740
rect 135220 187700 163504 187728
rect 135220 187688 135226 187700
rect 163498 187688 163504 187700
rect 163556 187688 163562 187740
rect 221366 187008 221372 187060
rect 221424 187048 221430 187060
rect 232130 187048 232136 187060
rect 221424 187020 232136 187048
rect 221424 187008 221430 187020
rect 232130 187008 232136 187020
rect 232188 187008 232194 187060
rect 184842 186940 184848 186992
rect 184900 186980 184906 186992
rect 247218 186980 247224 186992
rect 184900 186952 247224 186980
rect 184900 186940 184906 186952
rect 247218 186940 247224 186952
rect 247276 186940 247282 186992
rect 122742 186396 122748 186448
rect 122800 186436 122806 186448
rect 174630 186436 174636 186448
rect 122800 186408 174636 186436
rect 122800 186396 122806 186408
rect 174630 186396 174636 186408
rect 174688 186396 174694 186448
rect 108942 186328 108948 186380
rect 109000 186368 109006 186380
rect 193950 186368 193956 186380
rect 109000 186340 193956 186368
rect 109000 186328 109006 186340
rect 193950 186328 193956 186340
rect 194008 186328 194014 186380
rect 230382 185852 230388 185904
rect 230440 185892 230446 185904
rect 231854 185892 231860 185904
rect 230440 185864 231860 185892
rect 230440 185852 230446 185864
rect 231854 185852 231860 185864
rect 231912 185852 231918 185904
rect 217962 185648 217968 185700
rect 218020 185688 218026 185700
rect 229186 185688 229192 185700
rect 218020 185660 229192 185688
rect 218020 185648 218026 185660
rect 229186 185648 229192 185660
rect 229244 185648 229250 185700
rect 181530 185580 181536 185632
rect 181588 185620 181594 185632
rect 240226 185620 240232 185632
rect 181588 185592 240232 185620
rect 181588 185580 181594 185592
rect 240226 185580 240232 185592
rect 240284 185580 240290 185632
rect 240778 185580 240784 185632
rect 240836 185620 240842 185632
rect 296990 185620 296996 185632
rect 240836 185592 296996 185620
rect 240836 185580 240842 185592
rect 296990 185580 296996 185592
rect 297048 185580 297054 185632
rect 124122 184968 124128 185020
rect 124180 185008 124186 185020
rect 164878 185008 164884 185020
rect 124180 184980 164884 185008
rect 124180 184968 124186 184980
rect 164878 184968 164884 184980
rect 164936 184968 164942 185020
rect 106182 184900 106188 184952
rect 106240 184940 106246 184952
rect 182910 184940 182916 184952
rect 106240 184912 182916 184940
rect 106240 184900 106246 184912
rect 182910 184900 182916 184912
rect 182968 184900 182974 184952
rect 207658 184220 207664 184272
rect 207716 184260 207722 184272
rect 238754 184260 238760 184272
rect 207716 184232 238760 184260
rect 207716 184220 207722 184232
rect 238754 184220 238760 184232
rect 238812 184220 238818 184272
rect 276658 184220 276664 184272
rect 276716 184260 276722 184272
rect 292850 184260 292856 184272
rect 276716 184232 292856 184260
rect 276716 184220 276722 184232
rect 292850 184220 292856 184232
rect 292908 184220 292914 184272
rect 180150 184152 180156 184204
rect 180208 184192 180214 184204
rect 192478 184192 192484 184204
rect 180208 184164 192484 184192
rect 180208 184152 180214 184164
rect 192478 184152 192484 184164
rect 192536 184152 192542 184204
rect 217318 184152 217324 184204
rect 217376 184192 217382 184204
rect 284478 184192 284484 184204
rect 217376 184164 284484 184192
rect 217376 184152 217382 184164
rect 284478 184152 284484 184164
rect 284536 184152 284542 184204
rect 103422 183608 103428 183660
rect 103480 183648 103486 183660
rect 169018 183648 169024 183660
rect 103480 183620 169024 183648
rect 103480 183608 103486 183620
rect 169018 183608 169024 183620
rect 169076 183608 169082 183660
rect 128262 183540 128268 183592
rect 128320 183580 128326 183592
rect 214650 183580 214656 183592
rect 128320 183552 214656 183580
rect 128320 183540 128326 183552
rect 214650 183540 214656 183552
rect 214708 183540 214714 183592
rect 215202 182860 215208 182912
rect 215260 182900 215266 182912
rect 234706 182900 234712 182912
rect 215260 182872 234712 182900
rect 215260 182860 215266 182872
rect 234706 182860 234712 182872
rect 234764 182860 234770 182912
rect 282270 182860 282276 182912
rect 282328 182900 282334 182912
rect 294230 182900 294236 182912
rect 282328 182872 294236 182900
rect 282328 182860 282334 182872
rect 294230 182860 294236 182872
rect 294288 182860 294294 182912
rect 179322 182792 179328 182844
rect 179380 182832 179386 182844
rect 226334 182832 226340 182844
rect 179380 182804 226340 182832
rect 179380 182792 179386 182804
rect 226334 182792 226340 182804
rect 226392 182792 226398 182844
rect 242250 182792 242256 182844
rect 242308 182832 242314 182844
rect 253934 182832 253940 182844
rect 242308 182804 253940 182832
rect 242308 182792 242314 182804
rect 253934 182792 253940 182804
rect 253992 182792 253998 182844
rect 265618 182792 265624 182844
rect 265676 182832 265682 182844
rect 281626 182832 281632 182844
rect 265676 182804 281632 182832
rect 265676 182792 265682 182804
rect 281626 182792 281632 182804
rect 281684 182792 281690 182844
rect 282178 182792 282184 182844
rect 282236 182832 282242 182844
rect 309410 182832 309416 182844
rect 282236 182804 309416 182832
rect 282236 182792 282242 182804
rect 309410 182792 309416 182804
rect 309468 182792 309474 182844
rect 133138 182248 133144 182300
rect 133196 182288 133202 182300
rect 164510 182288 164516 182300
rect 133196 182260 164516 182288
rect 133196 182248 133202 182260
rect 164510 182248 164516 182260
rect 164568 182248 164574 182300
rect 148226 182180 148232 182232
rect 148284 182220 148290 182232
rect 214558 182220 214564 182232
rect 148284 182192 214564 182220
rect 148284 182180 148290 182192
rect 214558 182180 214564 182192
rect 214616 182180 214622 182232
rect 229738 182112 229744 182164
rect 229796 182152 229802 182164
rect 230750 182152 230756 182164
rect 229796 182124 230756 182152
rect 229796 182112 229802 182124
rect 230750 182112 230756 182124
rect 230808 182112 230814 182164
rect 233970 181568 233976 181620
rect 234028 181608 234034 181620
rect 245746 181608 245752 181620
rect 234028 181580 245752 181608
rect 234028 181568 234034 181580
rect 245746 181568 245752 181580
rect 245804 181568 245810 181620
rect 220078 181500 220084 181552
rect 220136 181540 220142 181552
rect 234890 181540 234896 181552
rect 220136 181512 234896 181540
rect 220136 181500 220142 181512
rect 234890 181500 234896 181512
rect 234948 181500 234954 181552
rect 273898 181500 273904 181552
rect 273956 181540 273962 181552
rect 295518 181540 295524 181552
rect 273956 181512 295524 181540
rect 273956 181500 273962 181512
rect 295518 181500 295524 181512
rect 295576 181500 295582 181552
rect 211798 181432 211804 181484
rect 211856 181472 211862 181484
rect 226886 181472 226892 181484
rect 211856 181444 226892 181472
rect 211856 181432 211862 181444
rect 226886 181432 226892 181444
rect 226944 181432 226950 181484
rect 235442 181432 235448 181484
rect 235500 181472 235506 181484
rect 248598 181472 248604 181484
rect 235500 181444 248604 181472
rect 235500 181432 235506 181444
rect 248598 181432 248604 181444
rect 248656 181432 248662 181484
rect 251818 181432 251824 181484
rect 251876 181472 251882 181484
rect 298278 181472 298284 181484
rect 251876 181444 298284 181472
rect 251876 181432 251882 181444
rect 298278 181432 298284 181444
rect 298336 181432 298342 181484
rect 125962 180888 125968 180940
rect 126020 180928 126026 180940
rect 170490 180928 170496 180940
rect 126020 180900 170496 180928
rect 126020 180888 126026 180900
rect 170490 180888 170496 180900
rect 170548 180888 170554 180940
rect 132402 180820 132408 180872
rect 132460 180860 132466 180872
rect 203610 180860 203616 180872
rect 132460 180832 203616 180860
rect 132460 180820 132466 180832
rect 203610 180820 203616 180832
rect 203668 180820 203674 180872
rect 222930 180208 222936 180260
rect 222988 180248 222994 180260
rect 240318 180248 240324 180260
rect 222988 180220 240324 180248
rect 222988 180208 222994 180220
rect 240318 180208 240324 180220
rect 240376 180208 240382 180260
rect 279418 180208 279424 180260
rect 279476 180248 279482 180260
rect 290090 180248 290096 180260
rect 279476 180220 290096 180248
rect 279476 180208 279482 180220
rect 290090 180208 290096 180220
rect 290148 180208 290154 180260
rect 186222 180140 186228 180192
rect 186280 180180 186286 180192
rect 223390 180180 223396 180192
rect 186280 180152 223396 180180
rect 186280 180140 186286 180152
rect 223390 180140 223396 180152
rect 223448 180140 223454 180192
rect 269850 180140 269856 180192
rect 269908 180180 269914 180192
rect 291470 180180 291476 180192
rect 269908 180152 291476 180180
rect 269908 180140 269914 180152
rect 291470 180140 291476 180152
rect 291528 180140 291534 180192
rect 169570 180072 169576 180124
rect 169628 180112 169634 180124
rect 226334 180112 226340 180124
rect 169628 180084 226340 180112
rect 169628 180072 169634 180084
rect 226334 180072 226340 180084
rect 226392 180072 226398 180124
rect 238110 180072 238116 180124
rect 238168 180112 238174 180124
rect 278774 180112 278780 180124
rect 238168 180084 278780 180112
rect 238168 180072 238174 180084
rect 278774 180072 278780 180084
rect 278832 180072 278838 180124
rect 229278 179936 229284 179988
rect 229336 179976 229342 179988
rect 237466 179976 237472 179988
rect 229336 179948 237472 179976
rect 229336 179936 229342 179948
rect 237466 179936 237472 179948
rect 237524 179936 237530 179988
rect 120994 179460 121000 179512
rect 121052 179500 121058 179512
rect 167822 179500 167828 179512
rect 121052 179472 167828 179500
rect 121052 179460 121058 179472
rect 167822 179460 167828 179472
rect 167880 179460 167886 179512
rect 112254 179392 112260 179444
rect 112312 179432 112318 179444
rect 171778 179432 171784 179444
rect 112312 179404 171784 179432
rect 112312 179392 112318 179404
rect 171778 179392 171784 179404
rect 171836 179392 171842 179444
rect 246298 179392 246304 179444
rect 246356 179432 246362 179444
rect 247126 179432 247132 179444
rect 246356 179404 247132 179432
rect 246356 179392 246362 179404
rect 247126 179392 247132 179404
rect 247184 179392 247190 179444
rect 574738 179324 574744 179376
rect 574796 179364 574802 179376
rect 580166 179364 580172 179376
rect 574796 179336 580172 179364
rect 574796 179324 574802 179336
rect 580166 179324 580172 179336
rect 580224 179324 580230 179376
rect 278774 179052 278780 179104
rect 278832 179092 278838 179104
rect 280338 179092 280344 179104
rect 278832 179064 280344 179092
rect 278832 179052 278838 179064
rect 280338 179052 280344 179064
rect 280396 179052 280402 179104
rect 278222 178916 278228 178968
rect 278280 178956 278286 178968
rect 278774 178956 278780 178968
rect 278280 178928 278780 178956
rect 278280 178916 278286 178928
rect 278774 178916 278780 178928
rect 278832 178916 278838 178968
rect 227070 178712 227076 178764
rect 227128 178752 227134 178764
rect 234798 178752 234804 178764
rect 227128 178724 234804 178752
rect 227128 178712 227134 178724
rect 234798 178712 234804 178724
rect 234856 178712 234862 178764
rect 199930 178644 199936 178696
rect 199988 178684 199994 178696
rect 245838 178684 245844 178696
rect 199988 178656 245844 178684
rect 199988 178644 199994 178656
rect 245838 178644 245844 178656
rect 245896 178644 245902 178696
rect 271230 178644 271236 178696
rect 271288 178684 271294 178696
rect 285858 178684 285864 178696
rect 271288 178656 285864 178684
rect 271288 178644 271294 178656
rect 285858 178644 285864 178656
rect 285916 178644 285922 178696
rect 124490 178100 124496 178152
rect 124548 178140 124554 178152
rect 187050 178140 187056 178152
rect 124548 178112 187056 178140
rect 124548 178100 124554 178112
rect 187050 178100 187056 178112
rect 187108 178100 187114 178152
rect 116946 178032 116952 178084
rect 117004 178072 117010 178084
rect 196802 178072 196808 178084
rect 117004 178044 196808 178072
rect 117004 178032 117010 178044
rect 196802 178032 196808 178044
rect 196860 178032 196866 178084
rect 298738 178032 298744 178084
rect 298796 178072 298802 178084
rect 299750 178072 299756 178084
rect 298796 178044 299756 178072
rect 298796 178032 298802 178044
rect 299750 178032 299756 178044
rect 299808 178032 299814 178084
rect 201126 177964 201132 178016
rect 201184 178004 201190 178016
rect 227806 178004 227812 178016
rect 201184 177976 227812 178004
rect 201184 177964 201190 177976
rect 227806 177964 227812 177976
rect 227864 177964 227870 178016
rect 286318 177964 286324 178016
rect 286376 178004 286382 178016
rect 287054 178004 287060 178016
rect 286376 177976 287060 178004
rect 286376 177964 286382 177976
rect 287054 177964 287060 177976
rect 287112 177964 287118 178016
rect 205542 177896 205548 177948
rect 205600 177936 205606 177948
rect 223482 177936 223488 177948
rect 205600 177908 223488 177936
rect 205600 177896 205606 177908
rect 223482 177896 223488 177908
rect 223540 177896 223546 177948
rect 226886 177352 226892 177404
rect 226944 177392 226950 177404
rect 238938 177392 238944 177404
rect 226944 177364 238944 177392
rect 226944 177352 226950 177364
rect 238938 177352 238944 177364
rect 238996 177352 239002 177404
rect 273990 177352 273996 177404
rect 274048 177392 274054 177404
rect 284570 177392 284576 177404
rect 274048 177364 284576 177392
rect 274048 177352 274054 177364
rect 284570 177352 284576 177364
rect 284628 177352 284634 177404
rect 228450 177284 228456 177336
rect 228508 177324 228514 177336
rect 233234 177324 233240 177336
rect 228508 177296 233240 177324
rect 228508 177284 228514 177296
rect 233234 177284 233240 177296
rect 233292 177284 233298 177336
rect 233878 177284 233884 177336
rect 233936 177324 233942 177336
rect 251174 177324 251180 177336
rect 233936 177296 251180 177324
rect 233936 177284 233942 177296
rect 251174 177284 251180 177296
rect 251232 177284 251238 177336
rect 268470 177284 268476 177336
rect 268528 177324 268534 177336
rect 283190 177324 283196 177336
rect 268528 177296 283196 177324
rect 268528 177284 268534 177296
rect 283190 177284 283196 177296
rect 283248 177284 283254 177336
rect 128170 176740 128176 176792
rect 128228 176780 128234 176792
rect 166442 176780 166448 176792
rect 128228 176752 166448 176780
rect 128228 176740 128234 176752
rect 166442 176740 166448 176752
rect 166500 176740 166506 176792
rect 136082 176672 136088 176724
rect 136140 176712 136146 176724
rect 136140 176684 142154 176712
rect 136140 176672 136146 176684
rect 142126 176644 142154 176684
rect 158990 176672 158996 176724
rect 159048 176712 159054 176724
rect 203518 176712 203524 176724
rect 159048 176684 203524 176712
rect 159048 176672 159054 176684
rect 203518 176672 203524 176684
rect 203576 176672 203582 176724
rect 213914 176644 213920 176656
rect 142126 176616 213920 176644
rect 213914 176604 213920 176616
rect 213972 176604 213978 176656
rect 188798 176536 188804 176588
rect 188856 176576 188862 176588
rect 228358 176576 228364 176588
rect 188856 176548 228364 176576
rect 188856 176536 188862 176548
rect 228358 176536 228364 176548
rect 228416 176536 228422 176588
rect 278130 176196 278136 176248
rect 278188 176236 278194 176248
rect 285950 176236 285956 176248
rect 278188 176208 285956 176236
rect 278188 176196 278194 176208
rect 285950 176196 285956 176208
rect 286008 176196 286014 176248
rect 226334 175992 226340 176044
rect 226392 176032 226398 176044
rect 233878 176032 233884 176044
rect 226392 176004 233884 176032
rect 226392 175992 226398 176004
rect 233878 175992 233884 176004
rect 233936 175992 233942 176044
rect 130746 175924 130752 175976
rect 130804 175964 130810 175976
rect 165522 175964 165528 175976
rect 130804 175936 165528 175964
rect 130804 175924 130810 175936
rect 165522 175924 165528 175936
rect 165580 175924 165586 175976
rect 231762 175924 231768 175976
rect 231820 175964 231826 175976
rect 245930 175964 245936 175976
rect 231820 175936 245936 175964
rect 231820 175924 231826 175936
rect 245930 175924 245936 175936
rect 245988 175924 245994 175976
rect 246390 175924 246396 175976
rect 246448 175964 246454 175976
rect 253934 175964 253940 175976
rect 246448 175936 253940 175964
rect 246448 175924 246454 175936
rect 253934 175924 253940 175936
rect 253992 175924 253998 175976
rect 223666 175788 223672 175840
rect 223724 175788 223730 175840
rect 163498 175176 163504 175228
rect 163556 175216 163562 175228
rect 213914 175216 213920 175228
rect 163556 175188 213920 175216
rect 163556 175176 163562 175188
rect 213914 175176 213920 175188
rect 213972 175176 213978 175228
rect 223684 175216 223712 175788
rect 279326 175420 279332 175432
rect 267706 175392 279332 175420
rect 243538 175312 243544 175364
rect 243596 175352 243602 175364
rect 264974 175352 264980 175364
rect 243596 175324 264980 175352
rect 243596 175312 243602 175324
rect 264974 175312 264980 175324
rect 265032 175312 265038 175364
rect 253934 175244 253940 175296
rect 253992 175284 253998 175296
rect 267706 175284 267734 175392
rect 279326 175380 279332 175392
rect 279384 175380 279390 175432
rect 253992 175256 267734 175284
rect 253992 175244 253998 175256
rect 223684 175188 229094 175216
rect 164510 175108 164516 175160
rect 164568 175148 164574 175160
rect 214006 175148 214012 175160
rect 164568 175120 214012 175148
rect 164568 175108 164574 175120
rect 214006 175108 214012 175120
rect 214064 175108 214070 175160
rect 229066 175148 229094 175188
rect 231762 175176 231768 175228
rect 231820 175216 231826 175228
rect 240134 175216 240140 175228
rect 231820 175188 240140 175216
rect 231820 175176 231826 175188
rect 240134 175176 240140 175188
rect 240192 175176 240198 175228
rect 230934 175148 230940 175160
rect 229066 175120 230940 175148
rect 230934 175108 230940 175120
rect 230992 175108 230998 175160
rect 229738 174768 229744 174820
rect 229796 174808 229802 174820
rect 232038 174808 232044 174820
rect 229796 174780 232044 174808
rect 229796 174768 229802 174780
rect 232038 174768 232044 174780
rect 232096 174768 232102 174820
rect 214098 174496 214104 174548
rect 214156 174536 214162 174548
rect 229278 174536 229284 174548
rect 214156 174508 229284 174536
rect 214156 174496 214162 174508
rect 229278 174496 229284 174508
rect 229336 174496 229342 174548
rect 255958 173952 255964 174004
rect 256016 173992 256022 174004
rect 264974 173992 264980 174004
rect 256016 173964 264980 173992
rect 256016 173952 256022 173964
rect 264974 173952 264980 173964
rect 265032 173952 265038 174004
rect 247770 173884 247776 173936
rect 247828 173924 247834 173936
rect 265066 173924 265072 173936
rect 247828 173896 265072 173924
rect 247828 173884 247834 173896
rect 265066 173884 265072 173896
rect 265124 173884 265130 173936
rect 165522 173816 165528 173868
rect 165580 173856 165586 173868
rect 214006 173856 214012 173868
rect 165580 173828 214012 173856
rect 165580 173816 165586 173828
rect 214006 173816 214012 173828
rect 214064 173816 214070 173868
rect 231578 173816 231584 173868
rect 231636 173856 231642 173868
rect 247034 173856 247040 173868
rect 231636 173828 247040 173856
rect 231636 173816 231642 173828
rect 247034 173816 247040 173828
rect 247092 173816 247098 173868
rect 203610 173748 203616 173800
rect 203668 173788 203674 173800
rect 213914 173788 213920 173800
rect 203668 173760 213920 173788
rect 203668 173748 203674 173760
rect 213914 173748 213920 173760
rect 213972 173748 213978 173800
rect 250530 172592 250536 172644
rect 250588 172632 250594 172644
rect 264974 172632 264980 172644
rect 250588 172604 264980 172632
rect 250588 172592 250594 172604
rect 264974 172592 264980 172604
rect 265032 172592 265038 172644
rect 247678 172524 247684 172576
rect 247736 172564 247742 172576
rect 265066 172564 265072 172576
rect 247736 172536 265072 172564
rect 247736 172524 247742 172536
rect 265066 172524 265072 172536
rect 265124 172524 265130 172576
rect 166258 172456 166264 172508
rect 166316 172496 166322 172508
rect 213914 172496 213920 172508
rect 166316 172468 213920 172496
rect 166316 172456 166322 172468
rect 213914 172456 213920 172468
rect 213972 172456 213978 172508
rect 236362 172456 236368 172508
rect 236420 172496 236426 172508
rect 238018 172496 238024 172508
rect 236420 172468 238024 172496
rect 236420 172456 236426 172468
rect 238018 172456 238024 172468
rect 238076 172456 238082 172508
rect 281534 172456 281540 172508
rect 281592 172496 281598 172508
rect 291378 172496 291384 172508
rect 281592 172468 291384 172496
rect 281592 172456 281598 172468
rect 291378 172456 291384 172468
rect 291436 172456 291442 172508
rect 167638 172388 167644 172440
rect 167696 172428 167702 172440
rect 215294 172428 215300 172440
rect 167696 172400 215300 172428
rect 167696 172388 167702 172400
rect 215294 172388 215300 172400
rect 215352 172388 215358 172440
rect 231118 172184 231124 172236
rect 231176 172224 231182 172236
rect 233326 172224 233332 172236
rect 231176 172196 233332 172224
rect 231176 172184 231182 172196
rect 233326 172184 233332 172196
rect 233384 172184 233390 172236
rect 231762 171844 231768 171896
rect 231820 171884 231826 171896
rect 237374 171884 237380 171896
rect 231820 171856 237380 171884
rect 231820 171844 231826 171856
rect 237374 171844 237380 171856
rect 237432 171844 237438 171896
rect 240870 171164 240876 171216
rect 240928 171204 240934 171216
rect 264974 171204 264980 171216
rect 240928 171176 264980 171204
rect 240928 171164 240934 171176
rect 264974 171164 264980 171176
rect 265032 171164 265038 171216
rect 238110 171096 238116 171148
rect 238168 171136 238174 171148
rect 265066 171136 265072 171148
rect 238168 171108 265072 171136
rect 238168 171096 238174 171108
rect 265066 171096 265072 171108
rect 265124 171096 265130 171148
rect 166442 171028 166448 171080
rect 166500 171068 166506 171080
rect 214006 171068 214012 171080
rect 166500 171040 214012 171068
rect 166500 171028 166506 171040
rect 214006 171028 214012 171040
rect 214064 171028 214070 171080
rect 170490 170960 170496 171012
rect 170548 171000 170554 171012
rect 213914 171000 213920 171012
rect 170548 170972 213920 171000
rect 170548 170960 170554 170972
rect 213914 170960 213920 170972
rect 213972 170960 213978 171012
rect 230658 170756 230664 170808
rect 230716 170796 230722 170808
rect 232130 170796 232136 170808
rect 230716 170768 232136 170796
rect 230716 170756 230722 170768
rect 232130 170756 232136 170768
rect 232188 170756 232194 170808
rect 231210 170008 231216 170060
rect 231268 170048 231274 170060
rect 233234 170048 233240 170060
rect 231268 170020 233240 170048
rect 231268 170008 231274 170020
rect 233234 170008 233240 170020
rect 233292 170008 233298 170060
rect 249242 169804 249248 169856
rect 249300 169844 249306 169856
rect 264974 169844 264980 169856
rect 249300 169816 264980 169844
rect 249300 169804 249306 169816
rect 264974 169804 264980 169816
rect 265032 169804 265038 169856
rect 232130 169736 232136 169788
rect 232188 169776 232194 169788
rect 236178 169776 236184 169788
rect 232188 169748 236184 169776
rect 232188 169736 232194 169748
rect 236178 169736 236184 169748
rect 236236 169736 236242 169788
rect 240962 169736 240968 169788
rect 241020 169776 241026 169788
rect 265066 169776 265072 169788
rect 241020 169748 265072 169776
rect 241020 169736 241026 169748
rect 265066 169736 265072 169748
rect 265124 169736 265130 169788
rect 169294 169668 169300 169720
rect 169352 169708 169358 169720
rect 214006 169708 214012 169720
rect 169352 169680 214012 169708
rect 169352 169668 169358 169680
rect 214006 169668 214012 169680
rect 214064 169668 214070 169720
rect 187050 169600 187056 169652
rect 187108 169640 187114 169652
rect 213914 169640 213920 169652
rect 187108 169612 213920 169640
rect 187108 169600 187114 169612
rect 213914 169600 213920 169612
rect 213972 169600 213978 169652
rect 281534 169600 281540 169652
rect 281592 169640 281598 169652
rect 287054 169640 287060 169652
rect 281592 169612 287060 169640
rect 281592 169600 281598 169612
rect 287054 169600 287060 169612
rect 287112 169600 287118 169652
rect 231670 169396 231676 169448
rect 231728 169436 231734 169448
rect 234890 169436 234896 169448
rect 231728 169408 234896 169436
rect 231728 169396 231734 169408
rect 234890 169396 234896 169408
rect 234948 169396 234954 169448
rect 238386 168512 238392 168564
rect 238444 168552 238450 168564
rect 238846 168552 238852 168564
rect 238444 168524 238852 168552
rect 238444 168512 238450 168524
rect 238846 168512 238852 168524
rect 238904 168512 238910 168564
rect 233970 168376 233976 168428
rect 234028 168416 234034 168428
rect 264974 168416 264980 168428
rect 234028 168388 264980 168416
rect 234028 168376 234034 168388
rect 264974 168376 264980 168388
rect 265032 168376 265038 168428
rect 167822 168308 167828 168360
rect 167880 168348 167886 168360
rect 214006 168348 214012 168360
rect 167880 168320 214012 168348
rect 167880 168308 167886 168320
rect 214006 168308 214012 168320
rect 214064 168308 214070 168360
rect 174630 168240 174636 168292
rect 174688 168280 174694 168292
rect 213914 168280 213920 168292
rect 174688 168252 213920 168280
rect 174688 168240 174694 168252
rect 213914 168240 213920 168252
rect 213972 168240 213978 168292
rect 230934 168240 230940 168292
rect 230992 168280 230998 168292
rect 233418 168280 233424 168292
rect 230992 168252 233424 168280
rect 230992 168240 230998 168252
rect 233418 168240 233424 168252
rect 233476 168240 233482 168292
rect 231670 167424 231676 167476
rect 231728 167464 231734 167476
rect 236270 167464 236276 167476
rect 231728 167436 236276 167464
rect 231728 167424 231734 167436
rect 236270 167424 236276 167436
rect 236328 167424 236334 167476
rect 242158 167084 242164 167136
rect 242216 167124 242222 167136
rect 264974 167124 264980 167136
rect 242216 167096 264980 167124
rect 242216 167084 242222 167096
rect 264974 167084 264980 167096
rect 265032 167084 265038 167136
rect 235258 167016 235264 167068
rect 235316 167056 235322 167068
rect 265066 167056 265072 167068
rect 235316 167028 265072 167056
rect 235316 167016 235322 167028
rect 265066 167016 265072 167028
rect 265124 167016 265130 167068
rect 169110 166948 169116 167000
rect 169168 166988 169174 167000
rect 213914 166988 213920 167000
rect 169168 166960 213920 166988
rect 169168 166948 169174 166960
rect 213914 166948 213920 166960
rect 213972 166948 213978 167000
rect 231302 166948 231308 167000
rect 231360 166988 231366 167000
rect 234798 166988 234804 167000
rect 231360 166960 234804 166988
rect 231360 166948 231366 166960
rect 234798 166948 234804 166960
rect 234856 166948 234862 167000
rect 196802 166880 196808 166932
rect 196860 166920 196866 166932
rect 214006 166920 214012 166932
rect 196860 166892 214012 166920
rect 196860 166880 196866 166892
rect 214006 166880 214012 166892
rect 214064 166880 214070 166932
rect 282822 166404 282828 166456
rect 282880 166444 282886 166456
rect 288710 166444 288716 166456
rect 282880 166416 288716 166444
rect 282880 166404 282886 166416
rect 288710 166404 288716 166416
rect 288768 166404 288774 166456
rect 230566 166268 230572 166320
rect 230624 166308 230630 166320
rect 230934 166308 230940 166320
rect 230624 166280 230940 166308
rect 230624 166268 230630 166280
rect 230934 166268 230940 166280
rect 230992 166268 230998 166320
rect 231670 166268 231676 166320
rect 231728 166308 231734 166320
rect 232130 166308 232136 166320
rect 231728 166280 232136 166308
rect 231728 166268 231734 166280
rect 232130 166268 232136 166280
rect 232188 166268 232194 166320
rect 239674 165656 239680 165708
rect 239732 165696 239738 165708
rect 264974 165696 264980 165708
rect 239732 165668 264980 165696
rect 239732 165656 239738 165668
rect 264974 165656 264980 165668
rect 265032 165656 265038 165708
rect 232774 165588 232780 165640
rect 232832 165628 232838 165640
rect 265066 165628 265072 165640
rect 232832 165600 265072 165628
rect 232832 165588 232838 165600
rect 265066 165588 265072 165600
rect 265124 165588 265130 165640
rect 166350 165520 166356 165572
rect 166408 165560 166414 165572
rect 214006 165560 214012 165572
rect 166408 165532 214012 165560
rect 166408 165520 166414 165532
rect 214006 165520 214012 165532
rect 214064 165520 214070 165572
rect 231118 165520 231124 165572
rect 231176 165560 231182 165572
rect 234706 165560 234712 165572
rect 231176 165532 234712 165560
rect 231176 165520 231182 165532
rect 234706 165520 234712 165532
rect 234764 165520 234770 165572
rect 282822 165520 282828 165572
rect 282880 165560 282886 165572
rect 302418 165560 302424 165572
rect 282880 165532 302424 165560
rect 282880 165520 282886 165532
rect 302418 165520 302424 165532
rect 302476 165520 302482 165572
rect 191282 165452 191288 165504
rect 191340 165492 191346 165504
rect 213914 165492 213920 165504
rect 191340 165464 213920 165492
rect 191340 165452 191346 165464
rect 213914 165452 213920 165464
rect 213972 165452 213978 165504
rect 236914 164840 236920 164892
rect 236972 164880 236978 164892
rect 265158 164880 265164 164892
rect 236972 164852 265164 164880
rect 236972 164840 236978 164852
rect 265158 164840 265164 164852
rect 265216 164840 265222 164892
rect 236638 164228 236644 164280
rect 236696 164268 236702 164280
rect 264974 164268 264980 164280
rect 236696 164240 264980 164268
rect 236696 164228 236702 164240
rect 264974 164228 264980 164240
rect 265032 164228 265038 164280
rect 3234 164160 3240 164212
rect 3292 164200 3298 164212
rect 15838 164200 15844 164212
rect 3292 164172 15844 164200
rect 3292 164160 3298 164172
rect 15838 164160 15844 164172
rect 15896 164160 15902 164212
rect 171778 164160 171784 164212
rect 171836 164200 171842 164212
rect 214006 164200 214012 164212
rect 171836 164172 214012 164200
rect 171836 164160 171842 164172
rect 214006 164160 214012 164172
rect 214064 164160 214070 164212
rect 231578 164160 231584 164212
rect 231636 164200 231642 164212
rect 249886 164200 249892 164212
rect 231636 164172 249892 164200
rect 231636 164160 231642 164172
rect 249886 164160 249892 164172
rect 249944 164160 249950 164212
rect 282822 164160 282828 164212
rect 282880 164200 282886 164212
rect 299750 164200 299756 164212
rect 282880 164172 299756 164200
rect 282880 164160 282886 164172
rect 299750 164160 299756 164172
rect 299808 164160 299814 164212
rect 177482 164092 177488 164144
rect 177540 164132 177546 164144
rect 213914 164132 213920 164144
rect 177540 164104 213920 164132
rect 177540 164092 177546 164104
rect 213914 164092 213920 164104
rect 213972 164092 213978 164144
rect 231486 163956 231492 164008
rect 231544 163996 231550 164008
rect 235994 163996 236000 164008
rect 231544 163968 236000 163996
rect 231544 163956 231550 163968
rect 235994 163956 236000 163968
rect 236052 163956 236058 164008
rect 282822 163140 282828 163192
rect 282880 163180 282886 163192
rect 288618 163180 288624 163192
rect 282880 163152 288624 163180
rect 282880 163140 282886 163152
rect 288618 163140 288624 163152
rect 288676 163140 288682 163192
rect 250622 162936 250628 162988
rect 250680 162976 250686 162988
rect 264974 162976 264980 162988
rect 250680 162948 264980 162976
rect 250680 162936 250686 162948
rect 264974 162936 264980 162948
rect 265032 162936 265038 162988
rect 245194 162868 245200 162920
rect 245252 162908 245258 162920
rect 265066 162908 265072 162920
rect 245252 162880 265072 162908
rect 245252 162868 245258 162880
rect 265066 162868 265072 162880
rect 265124 162868 265130 162920
rect 171962 162800 171968 162852
rect 172020 162840 172026 162852
rect 213914 162840 213920 162852
rect 172020 162812 213920 162840
rect 172020 162800 172026 162812
rect 213914 162800 213920 162812
rect 213972 162800 213978 162852
rect 231762 162800 231768 162852
rect 231820 162840 231826 162852
rect 247218 162840 247224 162852
rect 231820 162812 247224 162840
rect 231820 162800 231826 162812
rect 247218 162800 247224 162812
rect 247276 162800 247282 162852
rect 282730 162800 282736 162852
rect 282788 162840 282794 162852
rect 306558 162840 306564 162852
rect 282788 162812 306564 162840
rect 282788 162800 282794 162812
rect 306558 162800 306564 162812
rect 306616 162800 306622 162852
rect 185670 162732 185676 162784
rect 185728 162772 185734 162784
rect 214006 162772 214012 162784
rect 185728 162744 214012 162772
rect 185728 162732 185734 162744
rect 214006 162732 214012 162744
rect 214064 162732 214070 162784
rect 282822 162732 282828 162784
rect 282880 162772 282886 162784
rect 301130 162772 301136 162784
rect 282880 162744 301136 162772
rect 282880 162732 282886 162744
rect 301130 162732 301136 162744
rect 301188 162732 301194 162784
rect 232590 162120 232596 162172
rect 232648 162160 232654 162172
rect 241698 162160 241704 162172
rect 232648 162132 241704 162160
rect 232648 162120 232654 162132
rect 241698 162120 241704 162132
rect 241756 162120 241762 162172
rect 257338 161508 257344 161560
rect 257396 161548 257402 161560
rect 264974 161548 264980 161560
rect 257396 161520 264980 161548
rect 257396 161508 257402 161520
rect 264974 161508 264980 161520
rect 265032 161508 265038 161560
rect 246482 161440 246488 161492
rect 246540 161480 246546 161492
rect 265066 161480 265072 161492
rect 246540 161452 265072 161480
rect 246540 161440 246546 161452
rect 265066 161440 265072 161452
rect 265124 161440 265130 161492
rect 169202 161372 169208 161424
rect 169260 161412 169266 161424
rect 214006 161412 214012 161424
rect 169260 161384 214012 161412
rect 169260 161372 169266 161384
rect 214006 161372 214012 161384
rect 214064 161372 214070 161424
rect 231762 161372 231768 161424
rect 231820 161412 231826 161424
rect 240226 161412 240232 161424
rect 231820 161384 240232 161412
rect 231820 161372 231826 161384
rect 240226 161372 240232 161384
rect 240284 161372 240290 161424
rect 282730 161372 282736 161424
rect 282788 161412 282794 161424
rect 299566 161412 299572 161424
rect 282788 161384 299572 161412
rect 282788 161372 282794 161384
rect 299566 161372 299572 161384
rect 299624 161372 299630 161424
rect 193950 161304 193956 161356
rect 194008 161344 194014 161356
rect 213914 161344 213920 161356
rect 194008 161316 213920 161344
rect 194008 161304 194014 161316
rect 213914 161304 213920 161316
rect 213972 161304 213978 161356
rect 282822 161304 282828 161356
rect 282880 161344 282886 161356
rect 296990 161344 296996 161356
rect 282880 161316 296996 161344
rect 282880 161304 282886 161316
rect 296990 161304 296996 161316
rect 297048 161304 297054 161356
rect 231302 160964 231308 161016
rect 231360 161004 231366 161016
rect 233510 161004 233516 161016
rect 231360 160976 233516 161004
rect 231360 160964 231366 160976
rect 233510 160964 233516 160976
rect 233568 160964 233574 161016
rect 246390 160148 246396 160200
rect 246448 160188 246454 160200
rect 264974 160188 264980 160200
rect 246448 160160 264980 160188
rect 246448 160148 246454 160160
rect 264974 160148 264980 160160
rect 265032 160148 265038 160200
rect 240778 160080 240784 160132
rect 240836 160120 240842 160132
rect 265066 160120 265072 160132
rect 240836 160092 265072 160120
rect 240836 160080 240842 160092
rect 265066 160080 265072 160092
rect 265124 160080 265130 160132
rect 182910 160012 182916 160064
rect 182968 160052 182974 160064
rect 213914 160052 213920 160064
rect 182968 160024 213920 160052
rect 182968 160012 182974 160024
rect 213914 160012 213920 160024
rect 213972 160012 213978 160064
rect 231762 160012 231768 160064
rect 231820 160052 231826 160064
rect 251266 160052 251272 160064
rect 231820 160024 251272 160052
rect 231820 160012 231826 160024
rect 251266 160012 251272 160024
rect 251324 160012 251330 160064
rect 282454 160012 282460 160064
rect 282512 160052 282518 160064
rect 302510 160052 302516 160064
rect 282512 160024 302516 160052
rect 282512 160012 282518 160024
rect 302510 160012 302516 160024
rect 302568 160012 302574 160064
rect 195514 159944 195520 159996
rect 195572 159984 195578 159996
rect 214006 159984 214012 159996
rect 195572 159956 214012 159984
rect 195572 159944 195578 159956
rect 214006 159944 214012 159956
rect 214064 159944 214070 159996
rect 231670 159944 231676 159996
rect 231728 159984 231734 159996
rect 244550 159984 244556 159996
rect 231728 159956 244556 159984
rect 231728 159944 231734 159956
rect 244550 159944 244556 159956
rect 244608 159944 244614 159996
rect 282546 159740 282552 159792
rect 282604 159780 282610 159792
rect 285950 159780 285956 159792
rect 282604 159752 285956 159780
rect 282604 159740 282610 159752
rect 285950 159740 285956 159752
rect 286008 159740 286014 159792
rect 171870 159332 171876 159384
rect 171928 159372 171934 159384
rect 188338 159372 188344 159384
rect 171928 159344 188344 159372
rect 171928 159332 171934 159344
rect 188338 159332 188344 159344
rect 188396 159332 188402 159384
rect 244918 159332 244924 159384
rect 244976 159372 244982 159384
rect 265158 159372 265164 159384
rect 244976 159344 265164 159372
rect 244976 159332 244982 159344
rect 265158 159332 265164 159344
rect 265216 159332 265222 159384
rect 167730 158992 167736 159044
rect 167788 159032 167794 159044
rect 169202 159032 169208 159044
rect 167788 159004 169208 159032
rect 167788 158992 167794 159004
rect 169202 158992 169208 159004
rect 169260 158992 169266 159044
rect 260190 158720 260196 158772
rect 260248 158760 260254 158772
rect 264974 158760 264980 158772
rect 260248 158732 264980 158760
rect 260248 158720 260254 158732
rect 264974 158720 264980 158732
rect 265032 158720 265038 158772
rect 169018 158652 169024 158704
rect 169076 158692 169082 158704
rect 213914 158692 213920 158704
rect 169076 158664 213920 158692
rect 169076 158652 169082 158664
rect 213914 158652 213920 158664
rect 213972 158652 213978 158704
rect 282086 158652 282092 158704
rect 282144 158692 282150 158704
rect 292850 158692 292856 158704
rect 282144 158664 292856 158692
rect 282144 158652 282150 158664
rect 292850 158652 292856 158664
rect 292908 158652 292914 158704
rect 181530 158584 181536 158636
rect 181588 158624 181594 158636
rect 214006 158624 214012 158636
rect 181588 158596 214012 158624
rect 181588 158584 181594 158596
rect 214006 158584 214012 158596
rect 214064 158584 214070 158636
rect 231486 158108 231492 158160
rect 231544 158148 231550 158160
rect 233878 158148 233884 158160
rect 231544 158120 233884 158148
rect 231544 158108 231550 158120
rect 233878 158108 233884 158120
rect 233936 158108 233942 158160
rect 233878 157972 233884 158024
rect 233936 158012 233942 158024
rect 242250 158012 242256 158024
rect 233936 157984 242256 158012
rect 233936 157972 233942 157984
rect 242250 157972 242256 157984
rect 242308 157972 242314 158024
rect 253290 157972 253296 158024
rect 253348 158012 253354 158024
rect 265066 158012 265072 158024
rect 253348 157984 265072 158012
rect 253348 157972 253354 157984
rect 265066 157972 265072 157984
rect 265124 157972 265130 158024
rect 282270 157972 282276 158024
rect 282328 158012 282334 158024
rect 298370 158012 298376 158024
rect 282328 157984 298376 158012
rect 282328 157972 282334 157984
rect 298370 157972 298376 157984
rect 298428 157972 298434 158024
rect 251910 157360 251916 157412
rect 251968 157400 251974 157412
rect 264974 157400 264980 157412
rect 251968 157372 264980 157400
rect 251968 157360 251974 157372
rect 264974 157360 264980 157372
rect 265032 157360 265038 157412
rect 166534 157292 166540 157344
rect 166592 157332 166598 157344
rect 213914 157332 213920 157344
rect 166592 157304 213920 157332
rect 166592 157292 166598 157304
rect 213914 157292 213920 157304
rect 213972 157292 213978 157344
rect 231762 157292 231768 157344
rect 231820 157332 231826 157344
rect 242986 157332 242992 157344
rect 231820 157304 242992 157332
rect 231820 157292 231826 157304
rect 242986 157292 242992 157304
rect 243044 157292 243050 157344
rect 180334 157224 180340 157276
rect 180392 157264 180398 157276
rect 214006 157264 214012 157276
rect 180392 157236 214012 157264
rect 180392 157224 180398 157236
rect 214006 157224 214012 157236
rect 214064 157224 214070 157276
rect 231486 156612 231492 156664
rect 231544 156652 231550 156664
rect 240318 156652 240324 156664
rect 231544 156624 240324 156652
rect 231544 156612 231550 156624
rect 240318 156612 240324 156624
rect 240376 156612 240382 156664
rect 250438 156000 250444 156052
rect 250496 156040 250502 156052
rect 264974 156040 264980 156052
rect 250496 156012 264980 156040
rect 250496 156000 250502 156012
rect 264974 156000 264980 156012
rect 265032 156000 265038 156052
rect 241054 155932 241060 155984
rect 241112 155972 241118 155984
rect 265066 155972 265072 155984
rect 241112 155944 265072 155972
rect 241112 155932 241118 155944
rect 265066 155932 265072 155944
rect 265124 155932 265130 155984
rect 178862 155864 178868 155916
rect 178920 155904 178926 155916
rect 213914 155904 213920 155916
rect 178920 155876 213920 155904
rect 178920 155864 178926 155876
rect 213914 155864 213920 155876
rect 213972 155864 213978 155916
rect 282178 155864 282184 155916
rect 282236 155904 282242 155916
rect 309226 155904 309232 155916
rect 282236 155876 309232 155904
rect 282236 155864 282242 155876
rect 309226 155864 309232 155876
rect 309284 155864 309290 155916
rect 230750 155796 230756 155848
rect 230808 155836 230814 155848
rect 232498 155836 232504 155848
rect 230808 155808 232504 155836
rect 230808 155796 230814 155808
rect 232498 155796 232504 155808
rect 232556 155796 232562 155848
rect 282822 155796 282828 155848
rect 282880 155836 282886 155848
rect 303798 155836 303804 155848
rect 282880 155808 303804 155836
rect 282880 155796 282886 155808
rect 303798 155796 303804 155808
rect 303856 155796 303862 155848
rect 231762 155388 231768 155440
rect 231820 155428 231826 155440
rect 237466 155428 237472 155440
rect 231820 155400 237472 155428
rect 231820 155388 231826 155400
rect 237466 155388 237472 155400
rect 237524 155388 237530 155440
rect 239490 154640 239496 154692
rect 239548 154680 239554 154692
rect 264974 154680 264980 154692
rect 239548 154652 264980 154680
rect 239548 154640 239554 154652
rect 264974 154640 264980 154652
rect 265032 154640 265038 154692
rect 238202 154572 238208 154624
rect 238260 154612 238266 154624
rect 265158 154612 265164 154624
rect 238260 154584 265164 154612
rect 238260 154572 238266 154584
rect 265158 154572 265164 154584
rect 265216 154572 265222 154624
rect 231578 154504 231584 154556
rect 231636 154544 231642 154556
rect 245838 154544 245844 154556
rect 231636 154516 245844 154544
rect 231636 154504 231642 154516
rect 245838 154504 245844 154516
rect 245896 154504 245902 154556
rect 282362 154504 282368 154556
rect 282420 154544 282426 154556
rect 295610 154544 295616 154556
rect 282420 154516 295616 154544
rect 282420 154504 282426 154516
rect 295610 154504 295616 154516
rect 295668 154504 295674 154556
rect 282086 154436 282092 154488
rect 282144 154476 282150 154488
rect 294230 154476 294236 154488
rect 282144 154448 294236 154476
rect 282144 154436 282150 154448
rect 294230 154436 294236 154448
rect 294288 154436 294294 154488
rect 231670 154300 231676 154352
rect 231728 154340 231734 154352
rect 234062 154340 234068 154352
rect 231728 154312 234068 154340
rect 231728 154300 231734 154312
rect 234062 154300 234068 154312
rect 234120 154300 234126 154352
rect 234154 153824 234160 153876
rect 234212 153864 234218 153876
rect 265618 153864 265624 153876
rect 234212 153836 265624 153864
rect 234212 153824 234218 153836
rect 265618 153824 265624 153836
rect 265676 153824 265682 153876
rect 264514 153416 264520 153468
rect 264572 153456 264578 153468
rect 265802 153456 265808 153468
rect 264572 153428 265808 153456
rect 264572 153416 264578 153428
rect 265802 153416 265808 153428
rect 265860 153416 265866 153468
rect 203610 153212 203616 153264
rect 203668 153252 203674 153264
rect 213914 153252 213920 153264
rect 203668 153224 213920 153252
rect 203668 153212 203674 153224
rect 213914 153212 213920 153224
rect 213972 153212 213978 153264
rect 211890 152056 211896 152108
rect 211948 152096 211954 152108
rect 214006 152096 214012 152108
rect 211948 152068 214012 152096
rect 211948 152056 211954 152068
rect 214006 152056 214012 152068
rect 214064 152056 214070 152108
rect 238386 151892 238392 151904
rect 230768 151864 238392 151892
rect 230768 151836 230796 151864
rect 238386 151852 238392 151864
rect 238444 151852 238450 151904
rect 247862 151852 247868 151904
rect 247920 151892 247926 151904
rect 264974 151892 264980 151904
rect 247920 151864 264980 151892
rect 247920 151852 247926 151864
rect 264974 151852 264980 151864
rect 265032 151852 265038 151904
rect 166258 151784 166264 151836
rect 166316 151824 166322 151836
rect 213914 151824 213920 151836
rect 166316 151796 213920 151824
rect 166316 151784 166322 151796
rect 213914 151784 213920 151796
rect 213972 151784 213978 151836
rect 230750 151784 230756 151836
rect 230808 151784 230814 151836
rect 238018 151784 238024 151836
rect 238076 151824 238082 151836
rect 265066 151824 265072 151836
rect 238076 151796 265072 151824
rect 238076 151784 238082 151796
rect 265066 151784 265072 151796
rect 265124 151784 265130 151836
rect 231762 151716 231768 151768
rect 231820 151756 231826 151768
rect 244458 151756 244464 151768
rect 231820 151728 244464 151756
rect 231820 151716 231826 151728
rect 244458 151716 244464 151728
rect 244516 151716 244522 151768
rect 282822 151716 282828 151768
rect 282880 151756 282886 151768
rect 305178 151756 305184 151768
rect 282880 151728 305184 151756
rect 282880 151716 282886 151728
rect 305178 151716 305184 151728
rect 305236 151716 305242 151768
rect 184290 150492 184296 150544
rect 184348 150532 184354 150544
rect 214006 150532 214012 150544
rect 184348 150504 214012 150532
rect 184348 150492 184354 150504
rect 214006 150492 214012 150504
rect 214064 150492 214070 150544
rect 264514 150492 264520 150544
rect 264572 150532 264578 150544
rect 266262 150532 266268 150544
rect 264572 150504 266268 150532
rect 264572 150492 264578 150504
rect 266262 150492 266268 150504
rect 266320 150492 266326 150544
rect 169110 150424 169116 150476
rect 169168 150464 169174 150476
rect 213914 150464 213920 150476
rect 169168 150436 213920 150464
rect 169168 150424 169174 150436
rect 213914 150424 213920 150436
rect 213972 150424 213978 150476
rect 242434 150424 242440 150476
rect 242492 150464 242498 150476
rect 264974 150464 264980 150476
rect 242492 150436 264980 150464
rect 242492 150424 242498 150436
rect 264974 150424 264980 150436
rect 265032 150424 265038 150476
rect 169202 150356 169208 150408
rect 169260 150396 169266 150408
rect 214006 150396 214012 150408
rect 169260 150368 214012 150396
rect 169260 150356 169266 150368
rect 214006 150356 214012 150368
rect 214064 150356 214070 150408
rect 231762 150356 231768 150408
rect 231820 150396 231826 150408
rect 247126 150396 247132 150408
rect 231820 150368 247132 150396
rect 231820 150356 231826 150368
rect 247126 150356 247132 150368
rect 247184 150356 247190 150408
rect 2774 150288 2780 150340
rect 2832 150328 2838 150340
rect 4798 150328 4804 150340
rect 2832 150300 4804 150328
rect 2832 150288 2838 150300
rect 4798 150288 4804 150300
rect 4856 150288 4862 150340
rect 231486 150288 231492 150340
rect 231544 150328 231550 150340
rect 244274 150328 244280 150340
rect 231544 150300 244280 150328
rect 231544 150288 231550 150300
rect 244274 150288 244280 150300
rect 244332 150288 244338 150340
rect 203518 149676 203524 149728
rect 203576 149716 203582 149728
rect 213914 149716 213920 149728
rect 203576 149688 213920 149716
rect 203576 149676 203582 149688
rect 213914 149676 213920 149688
rect 213972 149676 213978 149728
rect 252002 149676 252008 149728
rect 252060 149716 252066 149728
rect 265066 149716 265072 149728
rect 252060 149688 265072 149716
rect 252060 149676 252066 149688
rect 265066 149676 265072 149688
rect 265124 149676 265130 149728
rect 245102 149064 245108 149116
rect 245160 149104 245166 149116
rect 264974 149104 264980 149116
rect 245160 149076 264980 149104
rect 245160 149064 245166 149076
rect 264974 149064 264980 149076
rect 265032 149064 265038 149116
rect 231762 148996 231768 149048
rect 231820 149036 231826 149048
rect 255314 149036 255320 149048
rect 231820 149008 255320 149036
rect 231820 148996 231826 149008
rect 255314 148996 255320 149008
rect 255372 148996 255378 149048
rect 282822 148928 282828 148980
rect 282880 148968 282886 148980
rect 290090 148968 290096 148980
rect 282880 148940 290096 148968
rect 282880 148928 282886 148940
rect 290090 148928 290096 148940
rect 290148 148928 290154 148980
rect 281534 148860 281540 148912
rect 281592 148900 281598 148912
rect 283190 148900 283196 148912
rect 281592 148872 283196 148900
rect 281592 148860 281598 148872
rect 283190 148860 283196 148872
rect 283248 148860 283254 148912
rect 231302 148316 231308 148368
rect 231360 148356 231366 148368
rect 248414 148356 248420 148368
rect 231360 148328 248420 148356
rect 231360 148316 231366 148328
rect 248414 148316 248420 148328
rect 248472 148316 248478 148368
rect 263134 147704 263140 147756
rect 263192 147744 263198 147756
rect 265710 147744 265716 147756
rect 263192 147716 265716 147744
rect 263192 147704 263198 147716
rect 265710 147704 265716 147716
rect 265768 147704 265774 147756
rect 166350 147636 166356 147688
rect 166408 147676 166414 147688
rect 213914 147676 213920 147688
rect 166408 147648 213920 147676
rect 166408 147636 166414 147648
rect 213914 147636 213920 147648
rect 213972 147636 213978 147688
rect 253474 147636 253480 147688
rect 253532 147676 253538 147688
rect 264974 147676 264980 147688
rect 253532 147648 264980 147676
rect 253532 147636 253538 147648
rect 264974 147636 264980 147648
rect 265032 147636 265038 147688
rect 282822 147568 282828 147620
rect 282880 147608 282886 147620
rect 307938 147608 307944 147620
rect 282880 147580 307944 147608
rect 282880 147568 282886 147580
rect 307938 147568 307944 147580
rect 307996 147568 308002 147620
rect 231118 146956 231124 147008
rect 231176 146996 231182 147008
rect 240962 146996 240968 147008
rect 231176 146968 240968 146996
rect 231176 146956 231182 146968
rect 240962 146956 240968 146968
rect 241020 146956 241026 147008
rect 232866 146888 232872 146940
rect 232924 146928 232930 146940
rect 254670 146928 254676 146940
rect 232924 146900 254676 146928
rect 232924 146888 232930 146900
rect 254670 146888 254676 146900
rect 254728 146888 254734 146940
rect 256234 146888 256240 146940
rect 256292 146928 256298 146940
rect 265158 146928 265164 146940
rect 256292 146900 265164 146928
rect 256292 146888 256298 146900
rect 265158 146888 265164 146900
rect 265216 146888 265222 146940
rect 258994 146820 259000 146872
rect 259052 146860 259058 146872
rect 265250 146860 265256 146872
rect 259052 146832 265256 146860
rect 259052 146820 259058 146832
rect 265250 146820 265256 146832
rect 265308 146820 265314 146872
rect 249426 146616 249432 146668
rect 249484 146656 249490 146668
rect 257338 146656 257344 146668
rect 249484 146628 257344 146656
rect 249484 146616 249490 146628
rect 257338 146616 257344 146628
rect 257396 146616 257402 146668
rect 185670 146276 185676 146328
rect 185728 146316 185734 146328
rect 213914 146316 213920 146328
rect 185728 146288 213920 146316
rect 185728 146276 185734 146288
rect 213914 146276 213920 146288
rect 213972 146276 213978 146328
rect 230750 146140 230756 146192
rect 230808 146180 230814 146192
rect 232590 146180 232596 146192
rect 230808 146152 232596 146180
rect 230808 146140 230814 146152
rect 232590 146140 232596 146152
rect 232648 146140 232654 146192
rect 170398 145528 170404 145580
rect 170456 145568 170462 145580
rect 209038 145568 209044 145580
rect 170456 145540 209044 145568
rect 170456 145528 170462 145540
rect 209038 145528 209044 145540
rect 209096 145528 209102 145580
rect 234062 144984 234068 145036
rect 234120 145024 234126 145036
rect 265066 145024 265072 145036
rect 234120 144996 265072 145024
rect 234120 144984 234126 144996
rect 265066 144984 265072 144996
rect 265124 144984 265130 145036
rect 203518 144916 203524 144968
rect 203576 144956 203582 144968
rect 213914 144956 213920 144968
rect 203576 144928 213920 144956
rect 203576 144916 203582 144928
rect 213914 144916 213920 144928
rect 213972 144916 213978 144968
rect 232498 144916 232504 144968
rect 232556 144956 232562 144968
rect 264974 144956 264980 144968
rect 232556 144928 264980 144956
rect 232556 144916 232562 144928
rect 264974 144916 264980 144928
rect 265032 144916 265038 144968
rect 282454 144848 282460 144900
rect 282512 144888 282518 144900
rect 310606 144888 310612 144900
rect 282512 144860 310612 144888
rect 282512 144848 282518 144860
rect 310606 144848 310612 144860
rect 310664 144848 310670 144900
rect 281902 144780 281908 144832
rect 281960 144820 281966 144832
rect 298278 144820 298284 144832
rect 281960 144792 298284 144820
rect 281960 144780 281966 144792
rect 298278 144780 298284 144792
rect 298336 144780 298342 144832
rect 230290 144168 230296 144220
rect 230348 144208 230354 144220
rect 242894 144208 242900 144220
rect 230348 144180 242900 144208
rect 230348 144168 230354 144180
rect 242894 144168 242900 144180
rect 242952 144168 242958 144220
rect 243814 144168 243820 144220
rect 243872 144208 243878 144220
rect 265158 144208 265164 144220
rect 243872 144180 265164 144208
rect 243872 144168 243878 144180
rect 265158 144168 265164 144180
rect 265216 144168 265222 144220
rect 204898 143624 204904 143676
rect 204956 143664 204962 143676
rect 213914 143664 213920 143676
rect 204956 143636 213920 143664
rect 204956 143624 204962 143636
rect 213914 143624 213920 143636
rect 213972 143624 213978 143676
rect 177482 143556 177488 143608
rect 177540 143596 177546 143608
rect 214006 143596 214012 143608
rect 177540 143568 214012 143596
rect 177540 143556 177546 143568
rect 214006 143556 214012 143568
rect 214064 143556 214070 143608
rect 240962 143556 240968 143608
rect 241020 143596 241026 143608
rect 264974 143596 264980 143608
rect 241020 143568 264980 143596
rect 241020 143556 241026 143568
rect 264974 143556 264980 143568
rect 265032 143556 265038 143608
rect 231762 143488 231768 143540
rect 231820 143528 231826 143540
rect 250070 143528 250076 143540
rect 231820 143500 250076 143528
rect 231820 143488 231826 143500
rect 250070 143488 250076 143500
rect 250128 143488 250134 143540
rect 282086 143488 282092 143540
rect 282144 143528 282150 143540
rect 295334 143528 295340 143540
rect 282144 143500 295340 143528
rect 282144 143488 282150 143500
rect 295334 143488 295340 143500
rect 295392 143488 295398 143540
rect 185578 142808 185584 142860
rect 185636 142848 185642 142860
rect 200758 142848 200764 142860
rect 185636 142820 200764 142848
rect 185636 142808 185642 142820
rect 200758 142808 200764 142820
rect 200816 142808 200822 142860
rect 230658 142808 230664 142860
rect 230716 142848 230722 142860
rect 251174 142848 251180 142860
rect 230716 142820 251180 142848
rect 230716 142808 230722 142820
rect 251174 142808 251180 142820
rect 251232 142808 251238 142860
rect 260282 142196 260288 142248
rect 260340 142236 260346 142248
rect 265066 142236 265072 142248
rect 260340 142208 265072 142236
rect 260340 142196 260346 142208
rect 265066 142196 265072 142208
rect 265124 142196 265130 142248
rect 207750 142128 207756 142180
rect 207808 142168 207814 142180
rect 213914 142168 213920 142180
rect 207808 142140 213920 142168
rect 207808 142128 207814 142140
rect 213914 142128 213920 142140
rect 213972 142128 213978 142180
rect 254670 142128 254676 142180
rect 254728 142168 254734 142180
rect 264974 142168 264980 142180
rect 254728 142140 264980 142168
rect 254728 142128 254734 142140
rect 264974 142128 264980 142140
rect 265032 142128 265038 142180
rect 281902 142060 281908 142112
rect 281960 142100 281966 142112
rect 284570 142100 284576 142112
rect 281960 142072 284576 142100
rect 281960 142060 281966 142072
rect 284570 142060 284576 142072
rect 284628 142060 284634 142112
rect 186958 141448 186964 141500
rect 187016 141488 187022 141500
rect 195238 141488 195244 141500
rect 187016 141460 195244 141488
rect 187016 141448 187022 141460
rect 195238 141448 195244 141460
rect 195296 141448 195302 141500
rect 231210 141448 231216 141500
rect 231268 141488 231274 141500
rect 254578 141488 254584 141500
rect 231268 141460 254584 141488
rect 231268 141448 231274 141460
rect 254578 141448 254584 141460
rect 254636 141448 254642 141500
rect 192570 141380 192576 141432
rect 192628 141420 192634 141432
rect 214006 141420 214012 141432
rect 192628 141392 214012 141420
rect 192628 141380 192634 141392
rect 214006 141380 214012 141392
rect 214064 141380 214070 141432
rect 230934 141380 230940 141432
rect 230992 141420 230998 141432
rect 255958 141420 255964 141432
rect 230992 141392 255964 141420
rect 230992 141380 230998 141392
rect 255958 141380 255964 141392
rect 256016 141380 256022 141432
rect 282270 141312 282276 141364
rect 282328 141352 282334 141364
rect 285858 141352 285864 141364
rect 282328 141324 285864 141352
rect 282328 141312 282334 141324
rect 285858 141312 285864 141324
rect 285916 141312 285922 141364
rect 261662 140836 261668 140888
rect 261720 140876 261726 140888
rect 265158 140876 265164 140888
rect 261720 140848 265164 140876
rect 261720 140836 261726 140848
rect 265158 140836 265164 140848
rect 265216 140836 265222 140888
rect 256050 140768 256056 140820
rect 256108 140808 256114 140820
rect 264974 140808 264980 140820
rect 256108 140780 264980 140808
rect 256108 140768 256114 140780
rect 264974 140768 264980 140780
rect 265032 140768 265038 140820
rect 231302 140700 231308 140752
rect 231360 140740 231366 140752
rect 236086 140740 236092 140752
rect 231360 140712 236092 140740
rect 231360 140700 231366 140712
rect 236086 140700 236092 140712
rect 236144 140700 236150 140752
rect 282270 140700 282276 140752
rect 282328 140740 282334 140752
rect 311986 140740 311992 140752
rect 282328 140712 311992 140740
rect 282328 140700 282334 140712
rect 311986 140700 311992 140712
rect 312044 140700 312050 140752
rect 281718 140632 281724 140684
rect 281776 140672 281782 140684
rect 300946 140672 300952 140684
rect 281776 140644 300952 140672
rect 281776 140632 281782 140644
rect 300946 140632 300952 140644
rect 301004 140632 301010 140684
rect 234338 140020 234344 140072
rect 234396 140060 234402 140072
rect 260190 140060 260196 140072
rect 234396 140032 260196 140060
rect 234396 140020 234402 140032
rect 260190 140020 260196 140032
rect 260248 140020 260254 140072
rect 210418 139476 210424 139528
rect 210476 139516 210482 139528
rect 214006 139516 214012 139528
rect 210476 139488 214012 139516
rect 210476 139476 210482 139488
rect 214006 139476 214012 139488
rect 214064 139476 214070 139528
rect 260374 139476 260380 139528
rect 260432 139516 260438 139528
rect 265894 139516 265900 139528
rect 260432 139488 265900 139516
rect 260432 139476 260438 139488
rect 265894 139476 265900 139488
rect 265952 139476 265958 139528
rect 206278 139408 206284 139460
rect 206336 139448 206342 139460
rect 213914 139448 213920 139460
rect 206336 139420 213920 139448
rect 206336 139408 206342 139420
rect 213914 139408 213920 139420
rect 213972 139408 213978 139460
rect 256142 139408 256148 139460
rect 256200 139448 256206 139460
rect 264974 139448 264980 139460
rect 256200 139420 264980 139448
rect 256200 139408 256206 139420
rect 264974 139408 264980 139420
rect 265032 139408 265038 139460
rect 231762 139340 231768 139392
rect 231820 139380 231826 139392
rect 255406 139380 255412 139392
rect 231820 139352 255412 139380
rect 231820 139340 231826 139352
rect 255406 139340 255412 139352
rect 255464 139340 255470 139392
rect 282270 139340 282276 139392
rect 282328 139380 282334 139392
rect 302234 139380 302240 139392
rect 282328 139352 302240 139380
rect 282328 139340 282334 139352
rect 302234 139340 302240 139352
rect 302292 139340 302298 139392
rect 282822 139272 282828 139324
rect 282880 139312 282886 139324
rect 296898 139312 296904 139324
rect 282880 139284 296904 139312
rect 282880 139272 282886 139284
rect 296898 139272 296904 139284
rect 296956 139272 296962 139324
rect 173158 138660 173164 138712
rect 173216 138700 173222 138712
rect 214466 138700 214472 138712
rect 173216 138672 214472 138700
rect 173216 138660 173222 138672
rect 214466 138660 214472 138672
rect 214524 138660 214530 138712
rect 250714 138660 250720 138712
rect 250772 138700 250778 138712
rect 265618 138700 265624 138712
rect 250772 138672 265624 138700
rect 250772 138660 250778 138672
rect 265618 138660 265624 138672
rect 265676 138660 265682 138712
rect 211798 137980 211804 138032
rect 211856 138020 211862 138032
rect 213914 138020 213920 138032
rect 211856 137992 213920 138020
rect 211856 137980 211862 137992
rect 213914 137980 213920 137992
rect 213972 137980 213978 138032
rect 257614 137980 257620 138032
rect 257672 138020 257678 138032
rect 264974 138020 264980 138032
rect 257672 137992 264980 138020
rect 257672 137980 257678 137992
rect 264974 137980 264980 137992
rect 265032 137980 265038 138032
rect 3510 137912 3516 137964
rect 3568 137952 3574 137964
rect 32398 137952 32404 137964
rect 3568 137924 32404 137952
rect 3568 137912 3574 137924
rect 32398 137912 32404 137924
rect 32456 137912 32462 137964
rect 231578 137912 231584 137964
rect 231636 137952 231642 137964
rect 252646 137952 252652 137964
rect 231636 137924 252652 137952
rect 231636 137912 231642 137924
rect 252646 137912 252652 137924
rect 252704 137912 252710 137964
rect 281718 137912 281724 137964
rect 281776 137952 281782 137964
rect 291470 137952 291476 137964
rect 281776 137924 291476 137952
rect 281776 137912 281782 137924
rect 291470 137912 291476 137924
rect 291528 137912 291534 137964
rect 231670 137572 231676 137624
rect 231728 137612 231734 137624
rect 238294 137612 238300 137624
rect 231728 137584 238300 137612
rect 231728 137572 231734 137584
rect 238294 137572 238300 137584
rect 238352 137572 238358 137624
rect 167730 137232 167736 137284
rect 167788 137272 167794 137284
rect 215938 137272 215944 137284
rect 167788 137244 215944 137272
rect 167788 137232 167794 137244
rect 215938 137232 215944 137244
rect 215996 137232 216002 137284
rect 178862 136620 178868 136672
rect 178920 136660 178926 136672
rect 213914 136660 213920 136672
rect 178920 136632 213920 136660
rect 178920 136620 178926 136632
rect 213914 136620 213920 136632
rect 213972 136620 213978 136672
rect 254578 136620 254584 136672
rect 254636 136660 254642 136672
rect 264974 136660 264980 136672
rect 254636 136632 264980 136660
rect 254636 136620 254642 136632
rect 264974 136620 264980 136632
rect 265032 136620 265038 136672
rect 231394 136552 231400 136604
rect 231452 136592 231458 136604
rect 247770 136592 247776 136604
rect 231452 136564 247776 136592
rect 231452 136552 231458 136564
rect 247770 136552 247776 136564
rect 247828 136552 247834 136604
rect 281902 136484 281908 136536
rect 281960 136524 281966 136536
rect 301038 136524 301044 136536
rect 281960 136496 301044 136524
rect 281960 136484 281966 136496
rect 301038 136484 301044 136496
rect 301096 136484 301102 136536
rect 231302 135940 231308 135992
rect 231360 135980 231366 135992
rect 239674 135980 239680 135992
rect 231360 135952 239680 135980
rect 231360 135940 231366 135952
rect 239674 135940 239680 135952
rect 239732 135940 239738 135992
rect 177390 135872 177396 135924
rect 177448 135912 177454 135924
rect 198182 135912 198188 135924
rect 177448 135884 198188 135912
rect 177448 135872 177454 135884
rect 198182 135872 198188 135884
rect 198240 135872 198246 135924
rect 239582 135872 239588 135924
rect 239640 135912 239646 135924
rect 265250 135912 265256 135924
rect 239640 135884 265256 135912
rect 239640 135872 239646 135884
rect 265250 135872 265256 135884
rect 265308 135872 265314 135924
rect 207658 135328 207664 135380
rect 207716 135368 207722 135380
rect 214006 135368 214012 135380
rect 207716 135340 214012 135368
rect 207716 135328 207722 135340
rect 214006 135328 214012 135340
rect 214064 135328 214070 135380
rect 202782 135260 202788 135312
rect 202840 135300 202846 135312
rect 213914 135300 213920 135312
rect 202840 135272 213920 135300
rect 202840 135260 202846 135272
rect 213914 135260 213920 135272
rect 213972 135260 213978 135312
rect 258718 135260 258724 135312
rect 258776 135300 258782 135312
rect 265066 135300 265072 135312
rect 258776 135272 265072 135300
rect 258776 135260 258782 135272
rect 265066 135260 265072 135272
rect 265124 135260 265130 135312
rect 231762 135192 231768 135244
rect 231820 135232 231826 135244
rect 260098 135232 260104 135244
rect 231820 135204 260104 135232
rect 231820 135192 231826 135204
rect 260098 135192 260104 135204
rect 260156 135192 260162 135244
rect 282086 135192 282092 135244
rect 282144 135232 282150 135244
rect 289814 135232 289820 135244
rect 282144 135204 289820 135232
rect 282144 135192 282150 135204
rect 289814 135192 289820 135204
rect 289872 135192 289878 135244
rect 231486 135124 231492 135176
rect 231544 135164 231550 135176
rect 247678 135164 247684 135176
rect 231544 135136 247684 135164
rect 231544 135124 231550 135136
rect 247678 135124 247684 135136
rect 247736 135124 247742 135176
rect 169018 134580 169024 134632
rect 169076 134620 169082 134632
rect 202782 134620 202788 134632
rect 169076 134592 202788 134620
rect 169076 134580 169082 134592
rect 202782 134580 202788 134592
rect 202840 134580 202846 134632
rect 177390 134512 177396 134564
rect 177448 134552 177454 134564
rect 211890 134552 211896 134564
rect 177448 134524 211896 134552
rect 177448 134512 177454 134524
rect 211890 134512 211896 134524
rect 211948 134512 211954 134564
rect 209314 133900 209320 133952
rect 209372 133940 209378 133952
rect 213914 133940 213920 133952
rect 209372 133912 213920 133940
rect 209372 133900 209378 133912
rect 213914 133900 213920 133912
rect 213972 133900 213978 133952
rect 257338 133900 257344 133952
rect 257396 133940 257402 133952
rect 264974 133940 264980 133952
rect 257396 133912 264980 133940
rect 257396 133900 257402 133912
rect 264974 133900 264980 133912
rect 265032 133900 265038 133952
rect 282270 133832 282276 133884
rect 282328 133872 282334 133884
rect 294138 133872 294144 133884
rect 282328 133844 294144 133872
rect 282328 133832 282334 133844
rect 294138 133832 294144 133844
rect 294196 133832 294202 133884
rect 282822 133764 282828 133816
rect 282880 133804 282886 133816
rect 292666 133804 292672 133816
rect 282880 133776 292672 133804
rect 282880 133764 282886 133776
rect 292666 133764 292672 133776
rect 292724 133764 292730 133816
rect 230566 133560 230572 133612
rect 230624 133600 230630 133612
rect 233970 133600 233976 133612
rect 230624 133572 233976 133600
rect 230624 133560 230630 133572
rect 233970 133560 233976 133572
rect 234028 133560 234034 133612
rect 231670 133220 231676 133272
rect 231728 133260 231734 133272
rect 238110 133260 238116 133272
rect 231728 133232 238116 133260
rect 231728 133220 231734 133232
rect 238110 133220 238116 133232
rect 238168 133220 238174 133272
rect 247678 132540 247684 132592
rect 247736 132580 247742 132592
rect 264974 132580 264980 132592
rect 247736 132552 264980 132580
rect 247736 132540 247742 132552
rect 264974 132540 264980 132552
rect 265032 132540 265038 132592
rect 206462 132472 206468 132524
rect 206520 132512 206526 132524
rect 213914 132512 213920 132524
rect 206520 132484 213920 132512
rect 206520 132472 206526 132484
rect 213914 132472 213920 132484
rect 213972 132472 213978 132524
rect 233878 132472 233884 132524
rect 233936 132512 233942 132524
rect 265066 132512 265072 132524
rect 233936 132484 265072 132512
rect 233936 132472 233942 132484
rect 265066 132472 265072 132484
rect 265124 132472 265130 132524
rect 231762 132404 231768 132456
rect 231820 132444 231826 132456
rect 257430 132444 257436 132456
rect 231820 132416 257436 132444
rect 231820 132404 231826 132416
rect 257430 132404 257436 132416
rect 257488 132404 257494 132456
rect 282730 132404 282736 132456
rect 282788 132444 282794 132456
rect 306650 132444 306656 132456
rect 282788 132416 306656 132444
rect 282788 132404 282794 132416
rect 306650 132404 306656 132416
rect 306708 132404 306714 132456
rect 282822 132336 282828 132388
rect 282880 132376 282886 132388
rect 299658 132376 299664 132388
rect 282880 132348 299664 132376
rect 282880 132336 282886 132348
rect 299658 132336 299664 132348
rect 299716 132336 299722 132388
rect 181530 131724 181536 131776
rect 181588 131764 181594 131776
rect 214650 131764 214656 131776
rect 181588 131736 214656 131764
rect 181588 131724 181594 131736
rect 214650 131724 214656 131736
rect 214708 131724 214714 131776
rect 232590 131180 232596 131232
rect 232648 131220 232654 131232
rect 232648 131192 238754 131220
rect 232648 131180 232654 131192
rect 191282 131112 191288 131164
rect 191340 131152 191346 131164
rect 213914 131152 213920 131164
rect 191340 131124 213920 131152
rect 191340 131112 191346 131124
rect 213914 131112 213920 131124
rect 213972 131112 213978 131164
rect 230934 131112 230940 131164
rect 230992 131152 230998 131164
rect 232774 131152 232780 131164
rect 230992 131124 232780 131152
rect 230992 131112 230998 131124
rect 232774 131112 232780 131124
rect 232832 131112 232838 131164
rect 238726 131152 238754 131192
rect 261570 131180 261576 131232
rect 261628 131220 261634 131232
rect 265066 131220 265072 131232
rect 261628 131192 265072 131220
rect 261628 131180 261634 131192
rect 265066 131180 265072 131192
rect 265124 131180 265130 131232
rect 264974 131152 264980 131164
rect 238726 131124 264980 131152
rect 264974 131112 264980 131124
rect 265032 131112 265038 131164
rect 231762 131044 231768 131096
rect 231820 131084 231826 131096
rect 249242 131084 249248 131096
rect 231820 131056 249248 131084
rect 231820 131044 231826 131056
rect 249242 131044 249248 131056
rect 249300 131044 249306 131096
rect 282270 131044 282276 131096
rect 282328 131084 282334 131096
rect 313366 131084 313372 131096
rect 282328 131056 313372 131084
rect 282328 131044 282334 131056
rect 313366 131044 313372 131056
rect 313424 131044 313430 131096
rect 281534 130568 281540 130620
rect 281592 130608 281598 130620
rect 284478 130608 284484 130620
rect 281592 130580 284484 130608
rect 281592 130568 281598 130580
rect 284478 130568 284484 130580
rect 284536 130568 284542 130620
rect 202322 129820 202328 129872
rect 202380 129860 202386 129872
rect 214006 129860 214012 129872
rect 202380 129832 214012 129860
rect 202380 129820 202386 129832
rect 214006 129820 214012 129832
rect 214064 129820 214070 129872
rect 171778 129752 171784 129804
rect 171836 129792 171842 129804
rect 213914 129792 213920 129804
rect 171836 129764 213920 129792
rect 171836 129752 171842 129764
rect 213914 129752 213920 129764
rect 213972 129752 213978 129804
rect 235350 129752 235356 129804
rect 235408 129792 235414 129804
rect 264974 129792 264980 129804
rect 235408 129764 264980 129792
rect 235408 129752 235414 129764
rect 264974 129752 264980 129764
rect 265032 129752 265038 129804
rect 231762 129684 231768 129736
rect 231820 129724 231826 129736
rect 264238 129724 264244 129736
rect 231820 129696 264244 129724
rect 231820 129684 231826 129696
rect 264238 129684 264244 129696
rect 264296 129684 264302 129736
rect 282086 129684 282092 129736
rect 282144 129724 282150 129736
rect 309410 129724 309416 129736
rect 282144 129696 309416 129724
rect 282144 129684 282150 129696
rect 309410 129684 309416 129696
rect 309468 129684 309474 129736
rect 230750 129548 230756 129600
rect 230808 129588 230814 129600
rect 236914 129588 236920 129600
rect 230808 129560 236920 129588
rect 230808 129548 230814 129560
rect 236914 129548 236920 129560
rect 236972 129548 236978 129600
rect 209222 128392 209228 128444
rect 209280 128432 209286 128444
rect 214006 128432 214012 128444
rect 209280 128404 214012 128432
rect 209280 128392 209286 128404
rect 214006 128392 214012 128404
rect 214064 128392 214070 128444
rect 178770 128324 178776 128376
rect 178828 128364 178834 128376
rect 213914 128364 213920 128376
rect 178828 128336 213920 128364
rect 178828 128324 178834 128336
rect 213914 128324 213920 128336
rect 213972 128324 213978 128376
rect 237006 128324 237012 128376
rect 237064 128364 237070 128376
rect 264974 128364 264980 128376
rect 237064 128336 264980 128364
rect 237064 128324 237070 128336
rect 264974 128324 264980 128336
rect 265032 128324 265038 128376
rect 231762 128256 231768 128308
rect 231820 128296 231826 128308
rect 242158 128296 242164 128308
rect 231820 128268 242164 128296
rect 231820 128256 231826 128268
rect 242158 128256 242164 128268
rect 242216 128256 242222 128308
rect 282822 128256 282828 128308
rect 282880 128296 282886 128308
rect 313274 128296 313280 128308
rect 282880 128268 313280 128296
rect 282880 128256 282886 128268
rect 313274 128256 313280 128268
rect 313332 128256 313338 128308
rect 282730 128188 282736 128240
rect 282788 128228 282794 128240
rect 287238 128228 287244 128240
rect 282788 128200 287244 128228
rect 282788 128188 282794 128200
rect 287238 128188 287244 128200
rect 287296 128188 287302 128240
rect 231118 127712 231124 127764
rect 231176 127752 231182 127764
rect 235258 127752 235264 127764
rect 231176 127724 235264 127752
rect 231176 127712 231182 127724
rect 235258 127712 235264 127724
rect 235316 127712 235322 127764
rect 250806 127576 250812 127628
rect 250864 127616 250870 127628
rect 258718 127616 258724 127628
rect 250864 127588 258724 127616
rect 250864 127576 250870 127588
rect 258718 127576 258724 127588
rect 258776 127576 258782 127628
rect 185762 127032 185768 127084
rect 185820 127072 185826 127084
rect 213914 127072 213920 127084
rect 185820 127044 213920 127072
rect 185820 127032 185826 127044
rect 213914 127032 213920 127044
rect 213972 127032 213978 127084
rect 173250 126964 173256 127016
rect 173308 127004 173314 127016
rect 214006 127004 214012 127016
rect 173308 126976 214012 127004
rect 173308 126964 173314 126976
rect 214006 126964 214012 126976
rect 214064 126964 214070 127016
rect 246298 126964 246304 127016
rect 246356 127004 246362 127016
rect 264974 127004 264980 127016
rect 246356 126976 264980 127004
rect 246356 126964 246362 126976
rect 264974 126964 264980 126976
rect 265032 126964 265038 127016
rect 231762 126896 231768 126948
rect 231820 126936 231826 126948
rect 239398 126936 239404 126948
rect 231820 126908 239404 126936
rect 231820 126896 231826 126908
rect 239398 126896 239404 126908
rect 239456 126896 239462 126948
rect 282270 126896 282276 126948
rect 282328 126936 282334 126948
rect 288526 126936 288532 126948
rect 282328 126908 288532 126936
rect 282328 126896 282334 126908
rect 288526 126896 288532 126908
rect 288584 126896 288590 126948
rect 249334 126284 249340 126336
rect 249392 126324 249398 126336
rect 265894 126324 265900 126336
rect 249392 126296 265900 126324
rect 249392 126284 249398 126296
rect 265894 126284 265900 126296
rect 265952 126284 265958 126336
rect 231394 126216 231400 126268
rect 231452 126256 231458 126268
rect 249426 126256 249432 126268
rect 231452 126228 249432 126256
rect 231452 126216 231458 126228
rect 249426 126216 249432 126228
rect 249484 126216 249490 126268
rect 196802 125672 196808 125724
rect 196860 125712 196866 125724
rect 214006 125712 214012 125724
rect 196860 125684 214012 125712
rect 196860 125672 196866 125684
rect 214006 125672 214012 125684
rect 214064 125672 214070 125724
rect 169202 125604 169208 125656
rect 169260 125644 169266 125656
rect 213914 125644 213920 125656
rect 169260 125616 213920 125644
rect 169260 125604 169266 125616
rect 213914 125604 213920 125616
rect 213972 125604 213978 125656
rect 258718 125604 258724 125656
rect 258776 125644 258782 125656
rect 264974 125644 264980 125656
rect 258776 125616 264980 125644
rect 258776 125604 258782 125616
rect 264974 125604 264980 125616
rect 265032 125604 265038 125656
rect 230474 125536 230480 125588
rect 230532 125576 230538 125588
rect 234154 125576 234160 125588
rect 230532 125548 234160 125576
rect 230532 125536 230538 125548
rect 234154 125536 234160 125548
rect 234212 125536 234218 125588
rect 282822 125536 282828 125588
rect 282880 125576 282886 125588
rect 314654 125576 314660 125588
rect 282880 125548 314660 125576
rect 282880 125536 282886 125548
rect 314654 125536 314660 125548
rect 314712 125536 314718 125588
rect 282086 125468 282092 125520
rect 282144 125508 282150 125520
rect 298186 125508 298192 125520
rect 282144 125480 298192 125508
rect 282144 125468 282150 125480
rect 298186 125468 298192 125480
rect 298244 125468 298250 125520
rect 186958 124856 186964 124908
rect 187016 124896 187022 124908
rect 206278 124896 206284 124908
rect 187016 124868 206284 124896
rect 187016 124856 187022 124868
rect 206278 124856 206284 124868
rect 206336 124856 206342 124908
rect 230658 124856 230664 124908
rect 230716 124896 230722 124908
rect 240778 124896 240784 124908
rect 230716 124868 240784 124896
rect 230716 124856 230722 124868
rect 240778 124856 240784 124868
rect 240836 124856 240842 124908
rect 176010 124176 176016 124228
rect 176068 124216 176074 124228
rect 213914 124216 213920 124228
rect 176068 124188 213920 124216
rect 176068 124176 176074 124188
rect 213914 124176 213920 124188
rect 213972 124176 213978 124228
rect 235258 124176 235264 124228
rect 235316 124216 235322 124228
rect 264974 124216 264980 124228
rect 235316 124188 264980 124216
rect 235316 124176 235322 124188
rect 264974 124176 264980 124188
rect 265032 124176 265038 124228
rect 231762 124108 231768 124160
rect 231820 124148 231826 124160
rect 261754 124148 261760 124160
rect 231820 124120 261760 124148
rect 231820 124108 231826 124120
rect 261754 124108 261760 124120
rect 261812 124108 261818 124160
rect 282270 124108 282276 124160
rect 282328 124148 282334 124160
rect 307754 124148 307760 124160
rect 282328 124120 307760 124148
rect 282328 124108 282334 124120
rect 307754 124108 307760 124120
rect 307812 124108 307818 124160
rect 231394 124040 231400 124092
rect 231452 124080 231458 124092
rect 250622 124080 250628 124092
rect 231452 124052 250628 124080
rect 231452 124040 231458 124052
rect 250622 124040 250628 124052
rect 250680 124040 250686 124092
rect 282822 124040 282828 124092
rect 282880 124080 282886 124092
rect 294046 124080 294052 124092
rect 282880 124052 294052 124080
rect 282880 124040 282886 124052
rect 294046 124040 294052 124052
rect 294104 124040 294110 124092
rect 210602 123088 210608 123140
rect 210660 123128 210666 123140
rect 214006 123128 214012 123140
rect 210660 123100 214012 123128
rect 210660 123088 210666 123100
rect 214006 123088 214012 123100
rect 214064 123088 214070 123140
rect 262122 123020 262128 123072
rect 262180 123060 262186 123072
rect 265066 123060 265072 123072
rect 262180 123032 265072 123060
rect 262180 123020 262186 123032
rect 265066 123020 265072 123032
rect 265124 123020 265130 123072
rect 174630 122816 174636 122868
rect 174688 122856 174694 122868
rect 213914 122856 213920 122868
rect 174688 122828 213920 122856
rect 174688 122816 174694 122828
rect 213914 122816 213920 122828
rect 213972 122816 213978 122868
rect 257522 122816 257528 122868
rect 257580 122856 257586 122868
rect 264974 122856 264980 122868
rect 257580 122828 264980 122856
rect 257580 122816 257586 122828
rect 264974 122816 264980 122828
rect 265032 122816 265038 122868
rect 231762 122748 231768 122800
rect 231820 122788 231826 122800
rect 263042 122788 263048 122800
rect 231820 122760 263048 122788
rect 231820 122748 231826 122760
rect 263042 122748 263048 122760
rect 263100 122748 263106 122800
rect 282454 122748 282460 122800
rect 282512 122788 282518 122800
rect 303614 122788 303620 122800
rect 282512 122760 303620 122788
rect 282512 122748 282518 122760
rect 303614 122748 303620 122760
rect 303672 122748 303678 122800
rect 231486 122680 231492 122732
rect 231544 122720 231550 122732
rect 244918 122720 244924 122732
rect 231544 122692 244924 122720
rect 231544 122680 231550 122692
rect 244918 122680 244924 122692
rect 244976 122680 244982 122732
rect 282638 122068 282644 122120
rect 282696 122108 282702 122120
rect 295518 122108 295524 122120
rect 282696 122080 295524 122108
rect 282696 122068 282702 122080
rect 295518 122068 295524 122080
rect 295576 122068 295582 122120
rect 199470 121524 199476 121576
rect 199528 121564 199534 121576
rect 214006 121564 214012 121576
rect 199528 121536 214012 121564
rect 199528 121524 199534 121536
rect 214006 121524 214012 121536
rect 214064 121524 214070 121576
rect 178954 121456 178960 121508
rect 179012 121496 179018 121508
rect 213914 121496 213920 121508
rect 179012 121468 213920 121496
rect 179012 121456 179018 121468
rect 213914 121456 213920 121468
rect 213972 121456 213978 121508
rect 252094 121456 252100 121508
rect 252152 121496 252158 121508
rect 264974 121496 264980 121508
rect 252152 121468 264980 121496
rect 252152 121456 252158 121468
rect 264974 121456 264980 121468
rect 265032 121456 265038 121508
rect 231762 121388 231768 121440
rect 231820 121428 231826 121440
rect 246482 121428 246488 121440
rect 231820 121400 246488 121428
rect 231820 121388 231826 121400
rect 246482 121388 246488 121400
rect 246540 121388 246546 121440
rect 282822 121388 282828 121440
rect 282880 121428 282886 121440
rect 305270 121428 305276 121440
rect 282880 121400 305276 121428
rect 282880 121388 282886 121400
rect 305270 121388 305276 121400
rect 305328 121388 305334 121440
rect 169294 120708 169300 120760
rect 169352 120748 169358 120760
rect 214834 120748 214840 120760
rect 169352 120720 214840 120748
rect 169352 120708 169358 120720
rect 214834 120708 214840 120720
rect 214892 120708 214898 120760
rect 191374 120096 191380 120148
rect 191432 120136 191438 120148
rect 213914 120136 213920 120148
rect 191432 120108 213920 120136
rect 191432 120096 191438 120108
rect 213914 120096 213920 120108
rect 213972 120096 213978 120148
rect 231394 120096 231400 120148
rect 231452 120136 231458 120148
rect 238018 120136 238024 120148
rect 231452 120108 238024 120136
rect 231452 120096 231458 120108
rect 238018 120096 238024 120108
rect 238076 120096 238082 120148
rect 240778 120096 240784 120148
rect 240836 120136 240842 120148
rect 264974 120136 264980 120148
rect 240836 120108 264980 120136
rect 240836 120096 240842 120108
rect 264974 120096 264980 120108
rect 265032 120096 265038 120148
rect 231486 120028 231492 120080
rect 231544 120068 231550 120080
rect 253290 120068 253296 120080
rect 231544 120040 253296 120068
rect 231544 120028 231550 120040
rect 253290 120028 253296 120040
rect 253348 120028 253354 120080
rect 282086 120028 282092 120080
rect 282144 120068 282150 120080
rect 285766 120068 285772 120080
rect 282144 120040 285772 120068
rect 282144 120028 282150 120040
rect 285766 120028 285772 120040
rect 285824 120028 285830 120080
rect 282178 119348 282184 119400
rect 282236 119388 282242 119400
rect 307846 119388 307852 119400
rect 282236 119360 307852 119388
rect 282236 119348 282242 119360
rect 307846 119348 307852 119360
rect 307904 119348 307910 119400
rect 206278 118736 206284 118788
rect 206336 118776 206342 118788
rect 213914 118776 213920 118788
rect 206336 118748 213920 118776
rect 206336 118736 206342 118748
rect 213914 118736 213920 118748
rect 213972 118736 213978 118788
rect 181622 118668 181628 118720
rect 181680 118708 181686 118720
rect 214006 118708 214012 118720
rect 181680 118680 214012 118708
rect 181680 118668 181686 118680
rect 214006 118668 214012 118680
rect 214064 118668 214070 118720
rect 230934 118668 230940 118720
rect 230992 118708 230998 118720
rect 234338 118708 234344 118720
rect 230992 118680 234344 118708
rect 230992 118668 230998 118680
rect 234338 118668 234344 118680
rect 234396 118668 234402 118720
rect 231578 118600 231584 118652
rect 231636 118640 231642 118652
rect 251910 118640 251916 118652
rect 231636 118612 251916 118640
rect 231636 118600 231642 118612
rect 251910 118600 251916 118612
rect 251968 118600 251974 118652
rect 281810 118396 281816 118448
rect 281868 118436 281874 118448
rect 284386 118436 284392 118448
rect 281868 118408 284392 118436
rect 281868 118396 281874 118408
rect 284386 118396 284392 118408
rect 284444 118396 284450 118448
rect 264330 117988 264336 118040
rect 264388 118028 264394 118040
rect 264606 118028 264612 118040
rect 264388 118000 264612 118028
rect 264388 117988 264394 118000
rect 264606 117988 264612 118000
rect 264664 117988 264670 118040
rect 230750 117920 230756 117972
rect 230808 117960 230814 117972
rect 241054 117960 241060 117972
rect 230808 117932 241060 117960
rect 230808 117920 230814 117932
rect 241054 117920 241060 117932
rect 241112 117920 241118 117972
rect 207842 117376 207848 117428
rect 207900 117416 207906 117428
rect 213914 117416 213920 117428
rect 207900 117388 213920 117416
rect 207900 117376 207906 117388
rect 213914 117376 213920 117388
rect 213972 117376 213978 117428
rect 253198 117376 253204 117428
rect 253256 117416 253262 117428
rect 265066 117416 265072 117428
rect 253256 117388 265072 117416
rect 253256 117376 253262 117388
rect 265066 117376 265072 117388
rect 265124 117376 265130 117428
rect 170582 117308 170588 117360
rect 170640 117348 170646 117360
rect 214006 117348 214012 117360
rect 170640 117320 214012 117348
rect 170640 117308 170646 117320
rect 214006 117308 214012 117320
rect 214064 117308 214070 117360
rect 242158 117308 242164 117360
rect 242216 117348 242222 117360
rect 264974 117348 264980 117360
rect 242216 117320 264980 117348
rect 242216 117308 242222 117320
rect 264974 117308 264980 117320
rect 265032 117308 265038 117360
rect 231762 117240 231768 117292
rect 231820 117280 231826 117292
rect 242250 117280 242256 117292
rect 231820 117252 242256 117280
rect 231820 117240 231826 117252
rect 242250 117240 242256 117252
rect 242308 117240 242314 117292
rect 282822 117240 282828 117292
rect 282880 117280 282886 117292
rect 292758 117280 292764 117292
rect 282880 117252 292764 117280
rect 282880 117240 282886 117252
rect 292758 117240 292764 117252
rect 292816 117240 292822 117292
rect 231486 117172 231492 117224
rect 231544 117212 231550 117224
rect 236822 117212 236828 117224
rect 231544 117184 236828 117212
rect 231544 117172 231550 117184
rect 236822 117172 236828 117184
rect 236880 117172 236886 117224
rect 282362 117104 282368 117156
rect 282420 117144 282426 117156
rect 287146 117144 287152 117156
rect 282420 117116 287152 117144
rect 282420 117104 282426 117116
rect 287146 117104 287152 117116
rect 287204 117104 287210 117156
rect 206370 116016 206376 116068
rect 206428 116056 206434 116068
rect 214006 116056 214012 116068
rect 206428 116028 214012 116056
rect 206428 116016 206434 116028
rect 214006 116016 214012 116028
rect 214064 116016 214070 116068
rect 263226 116016 263232 116068
rect 263284 116056 263290 116068
rect 265066 116056 265072 116068
rect 263284 116028 265072 116056
rect 263284 116016 263290 116028
rect 265066 116016 265072 116028
rect 265124 116016 265130 116068
rect 189810 115948 189816 116000
rect 189868 115988 189874 116000
rect 213914 115988 213920 116000
rect 189868 115960 213920 115988
rect 189868 115948 189874 115960
rect 213914 115948 213920 115960
rect 213972 115948 213978 116000
rect 253290 115948 253296 116000
rect 253348 115988 253354 116000
rect 264974 115988 264980 116000
rect 253348 115960 264980 115988
rect 253348 115948 253354 115960
rect 264974 115948 264980 115960
rect 265032 115948 265038 116000
rect 203702 115880 203708 115932
rect 203760 115920 203766 115932
rect 204990 115920 204996 115932
rect 203760 115892 204996 115920
rect 203760 115880 203766 115892
rect 204990 115880 204996 115892
rect 205048 115880 205054 115932
rect 231486 115880 231492 115932
rect 231544 115920 231550 115932
rect 263134 115920 263140 115932
rect 231544 115892 263140 115920
rect 231544 115880 231550 115892
rect 263134 115880 263140 115892
rect 263192 115880 263198 115932
rect 282822 115880 282828 115932
rect 282880 115920 282886 115932
rect 302326 115920 302332 115932
rect 282880 115892 302332 115920
rect 282880 115880 282886 115892
rect 302326 115880 302332 115892
rect 302384 115880 302390 115932
rect 230934 115812 230940 115864
rect 230992 115852 230998 115864
rect 238202 115852 238208 115864
rect 230992 115824 238208 115852
rect 230992 115812 230998 115824
rect 238202 115812 238208 115824
rect 238260 115812 238266 115864
rect 282270 115336 282276 115388
rect 282328 115376 282334 115388
rect 285674 115376 285680 115388
rect 282328 115348 285680 115376
rect 282328 115336 282334 115348
rect 285674 115336 285680 115348
rect 285732 115336 285738 115388
rect 195330 115200 195336 115252
rect 195388 115240 195394 115252
rect 214926 115240 214932 115252
rect 195388 115212 214932 115240
rect 195388 115200 195394 115212
rect 214926 115200 214932 115212
rect 214984 115200 214990 115252
rect 205082 114520 205088 114572
rect 205140 114560 205146 114572
rect 213914 114560 213920 114572
rect 205140 114532 213920 114560
rect 205140 114520 205146 114532
rect 213914 114520 213920 114532
rect 213972 114520 213978 114572
rect 242342 114520 242348 114572
rect 242400 114560 242406 114572
rect 264974 114560 264980 114572
rect 242400 114532 264980 114560
rect 242400 114520 242406 114532
rect 264974 114520 264980 114532
rect 265032 114520 265038 114572
rect 231670 114452 231676 114504
rect 231728 114492 231734 114504
rect 239490 114492 239496 114504
rect 231728 114464 239496 114492
rect 231728 114452 231734 114464
rect 239490 114452 239496 114464
rect 239548 114452 239554 114504
rect 230566 114112 230572 114164
rect 230624 114152 230630 114164
rect 232682 114152 232688 114164
rect 230624 114124 232688 114152
rect 230624 114112 230630 114124
rect 232682 114112 232688 114124
rect 232740 114112 232746 114164
rect 188430 113228 188436 113280
rect 188488 113268 188494 113280
rect 214006 113268 214012 113280
rect 188488 113240 214012 113268
rect 188488 113228 188494 113240
rect 214006 113228 214012 113240
rect 214064 113228 214070 113280
rect 249242 113228 249248 113280
rect 249300 113268 249306 113280
rect 265066 113268 265072 113280
rect 249300 113240 265072 113268
rect 249300 113228 249306 113240
rect 265066 113228 265072 113240
rect 265124 113228 265130 113280
rect 176194 113160 176200 113212
rect 176252 113200 176258 113212
rect 213914 113200 213920 113212
rect 176252 113172 213920 113200
rect 176252 113160 176258 113172
rect 213914 113160 213920 113172
rect 213972 113160 213978 113212
rect 234154 113160 234160 113212
rect 234212 113200 234218 113212
rect 264974 113200 264980 113212
rect 234212 113172 264980 113200
rect 234212 113160 234218 113172
rect 264974 113160 264980 113172
rect 265032 113160 265038 113212
rect 231762 113092 231768 113144
rect 231820 113132 231826 113144
rect 264514 113132 264520 113144
rect 231820 113104 264520 113132
rect 231820 113092 231826 113104
rect 264514 113092 264520 113104
rect 264572 113092 264578 113144
rect 282822 113092 282828 113144
rect 282880 113132 282886 113144
rect 303706 113132 303712 113144
rect 282880 113104 303712 113132
rect 282880 113092 282886 113104
rect 303706 113092 303712 113104
rect 303764 113092 303770 113144
rect 231302 113024 231308 113076
rect 231360 113064 231366 113076
rect 258994 113064 259000 113076
rect 231360 113036 259000 113064
rect 231360 113024 231366 113036
rect 258994 113024 259000 113036
rect 259052 113024 259058 113076
rect 281994 113024 282000 113076
rect 282052 113064 282058 113076
rect 291194 113064 291200 113076
rect 282052 113036 291200 113064
rect 282052 113024 282058 113036
rect 291194 113024 291200 113036
rect 291252 113024 291258 113076
rect 184382 112412 184388 112464
rect 184440 112452 184446 112464
rect 214834 112452 214840 112464
rect 184440 112424 214840 112452
rect 184440 112412 184446 112424
rect 214834 112412 214840 112424
rect 214892 112412 214898 112464
rect 187050 111800 187056 111852
rect 187108 111840 187114 111852
rect 213914 111840 213920 111852
rect 187108 111812 213920 111840
rect 187108 111800 187114 111812
rect 213914 111800 213920 111812
rect 213972 111800 213978 111852
rect 260466 111800 260472 111852
rect 260524 111840 260530 111852
rect 264974 111840 264980 111852
rect 260524 111812 264980 111840
rect 260524 111800 260530 111812
rect 264974 111800 264980 111812
rect 265032 111800 265038 111852
rect 168282 111732 168288 111784
rect 168340 111772 168346 111784
rect 169110 111772 169116 111784
rect 168340 111744 169116 111772
rect 168340 111732 168346 111744
rect 169110 111732 169116 111744
rect 169168 111732 169174 111784
rect 231762 111732 231768 111784
rect 231820 111772 231826 111784
rect 247862 111772 247868 111784
rect 231820 111744 247868 111772
rect 231820 111732 231826 111744
rect 247862 111732 247868 111744
rect 247920 111732 247926 111784
rect 282822 111732 282828 111784
rect 282880 111772 282886 111784
rect 289998 111772 290004 111784
rect 282880 111744 290004 111772
rect 282880 111732 282886 111744
rect 289998 111732 290004 111744
rect 290056 111732 290062 111784
rect 231670 111664 231676 111716
rect 231728 111704 231734 111716
rect 235442 111704 235448 111716
rect 231728 111676 235448 111704
rect 231728 111664 231734 111676
rect 235442 111664 235448 111676
rect 235500 111664 235506 111716
rect 209130 110508 209136 110560
rect 209188 110548 209194 110560
rect 213914 110548 213920 110560
rect 209188 110520 213920 110548
rect 209188 110508 209194 110520
rect 213914 110508 213920 110520
rect 213972 110508 213978 110560
rect 255958 110508 255964 110560
rect 256016 110548 256022 110560
rect 264974 110548 264980 110560
rect 256016 110520 264980 110548
rect 256016 110508 256022 110520
rect 264974 110508 264980 110520
rect 265032 110508 265038 110560
rect 170490 110440 170496 110492
rect 170548 110480 170554 110492
rect 214006 110480 214012 110492
rect 170548 110452 214012 110480
rect 170548 110440 170554 110452
rect 214006 110440 214012 110452
rect 214064 110440 214070 110492
rect 244918 110440 244924 110492
rect 244976 110480 244982 110492
rect 265066 110480 265072 110492
rect 244976 110452 265072 110480
rect 244976 110440 244982 110452
rect 265066 110440 265072 110452
rect 265124 110440 265130 110492
rect 167822 110372 167828 110424
rect 167880 110412 167886 110424
rect 184290 110412 184296 110424
rect 167880 110384 184296 110412
rect 167880 110372 167886 110384
rect 184290 110372 184296 110384
rect 184348 110372 184354 110424
rect 231762 110372 231768 110424
rect 231820 110412 231826 110424
rect 252002 110412 252008 110424
rect 231820 110384 252008 110412
rect 231820 110372 231826 110384
rect 252002 110372 252008 110384
rect 252060 110372 252066 110424
rect 282270 110372 282276 110424
rect 282328 110412 282334 110424
rect 296806 110412 296812 110424
rect 282328 110384 296812 110412
rect 282328 110372 282334 110384
rect 296806 110372 296812 110384
rect 296864 110372 296870 110424
rect 231210 110304 231216 110356
rect 231268 110344 231274 110356
rect 242434 110344 242440 110356
rect 231268 110316 242440 110344
rect 231268 110304 231274 110316
rect 242434 110304 242440 110316
rect 242492 110304 242498 110356
rect 282822 109760 282828 109812
rect 282880 109800 282886 109812
rect 287330 109800 287336 109812
rect 282880 109772 287336 109800
rect 282880 109760 282886 109772
rect 287330 109760 287336 109772
rect 287388 109760 287394 109812
rect 200850 109080 200856 109132
rect 200908 109120 200914 109132
rect 202322 109120 202328 109132
rect 200908 109092 202328 109120
rect 200908 109080 200914 109092
rect 202322 109080 202328 109092
rect 202380 109080 202386 109132
rect 173342 109012 173348 109064
rect 173400 109052 173406 109064
rect 213914 109052 213920 109064
rect 173400 109024 213920 109052
rect 173400 109012 173406 109024
rect 213914 109012 213920 109024
rect 213972 109012 213978 109064
rect 257430 109012 257436 109064
rect 257488 109052 257494 109064
rect 264974 109052 264980 109064
rect 257488 109024 264980 109052
rect 257488 109012 257494 109024
rect 264974 109012 264980 109024
rect 265032 109012 265038 109064
rect 231394 108944 231400 108996
rect 231452 108984 231458 108996
rect 256234 108984 256240 108996
rect 231452 108956 256240 108984
rect 231452 108944 231458 108956
rect 256234 108944 256240 108956
rect 256292 108944 256298 108996
rect 231762 108876 231768 108928
rect 231820 108916 231826 108928
rect 245102 108916 245108 108928
rect 231820 108888 245108 108916
rect 231820 108876 231826 108888
rect 245102 108876 245108 108888
rect 245160 108876 245166 108928
rect 281718 108876 281724 108928
rect 281776 108916 281782 108928
rect 284294 108916 284300 108928
rect 281776 108888 284300 108916
rect 281776 108876 281782 108888
rect 284294 108876 284300 108888
rect 284352 108876 284358 108928
rect 282270 108264 282276 108316
rect 282328 108304 282334 108316
rect 296714 108304 296720 108316
rect 282328 108276 296720 108304
rect 282328 108264 282334 108276
rect 296714 108264 296720 108276
rect 296772 108264 296778 108316
rect 210510 107720 210516 107772
rect 210568 107760 210574 107772
rect 214006 107760 214012 107772
rect 210568 107732 214012 107760
rect 210568 107720 210574 107732
rect 214006 107720 214012 107732
rect 214064 107720 214070 107772
rect 258994 107720 259000 107772
rect 259052 107760 259058 107772
rect 264974 107760 264980 107772
rect 259052 107732 264980 107760
rect 259052 107720 259058 107732
rect 264974 107720 264980 107732
rect 265032 107720 265038 107772
rect 202322 107652 202328 107704
rect 202380 107692 202386 107704
rect 213914 107692 213920 107704
rect 202380 107664 213920 107692
rect 202380 107652 202386 107664
rect 213914 107652 213920 107664
rect 213972 107652 213978 107704
rect 250530 107652 250536 107704
rect 250588 107692 250594 107704
rect 265066 107692 265072 107704
rect 250588 107664 265072 107692
rect 250588 107652 250594 107664
rect 265066 107652 265072 107664
rect 265124 107652 265130 107704
rect 231210 107584 231216 107636
rect 231268 107624 231274 107636
rect 253474 107624 253480 107636
rect 231268 107596 253480 107624
rect 231268 107584 231274 107596
rect 253474 107584 253480 107596
rect 253532 107584 253538 107636
rect 231762 107516 231768 107568
rect 231820 107556 231826 107568
rect 250714 107556 250720 107568
rect 231820 107528 250720 107556
rect 231820 107516 231826 107528
rect 250714 107516 250720 107528
rect 250772 107516 250778 107568
rect 184474 106360 184480 106412
rect 184532 106400 184538 106412
rect 213914 106400 213920 106412
rect 184532 106372 213920 106400
rect 184532 106360 184538 106372
rect 213914 106360 213920 106372
rect 213972 106360 213978 106412
rect 253382 106360 253388 106412
rect 253440 106400 253446 106412
rect 264974 106400 264980 106412
rect 253440 106372 264980 106400
rect 253440 106360 253446 106372
rect 264974 106360 264980 106372
rect 265032 106360 265038 106412
rect 167822 106292 167828 106344
rect 167880 106332 167886 106344
rect 214006 106332 214012 106344
rect 167880 106304 214012 106332
rect 167880 106292 167886 106304
rect 214006 106292 214012 106304
rect 214064 106292 214070 106344
rect 251910 106292 251916 106344
rect 251968 106332 251974 106344
rect 265066 106332 265072 106344
rect 251968 106304 265072 106332
rect 251968 106292 251974 106304
rect 265066 106292 265072 106304
rect 265124 106292 265130 106344
rect 231762 106224 231768 106276
rect 231820 106264 231826 106276
rect 260374 106264 260380 106276
rect 231820 106236 260380 106264
rect 231820 106224 231826 106236
rect 260374 106224 260380 106236
rect 260432 106224 260438 106276
rect 282822 106224 282828 106276
rect 282880 106264 282886 106276
rect 291286 106264 291292 106276
rect 282880 106236 291292 106264
rect 282880 106224 282886 106236
rect 291286 106224 291292 106236
rect 291344 106224 291350 106276
rect 166534 105544 166540 105596
rect 166592 105584 166598 105596
rect 204898 105584 204904 105596
rect 166592 105556 204904 105584
rect 166592 105544 166598 105556
rect 204898 105544 204904 105556
rect 204956 105544 204962 105596
rect 230750 105544 230756 105596
rect 230808 105584 230814 105596
rect 253934 105584 253940 105596
rect 230808 105556 253940 105584
rect 230808 105544 230814 105556
rect 253934 105544 253940 105556
rect 253992 105544 253998 105596
rect 204990 104932 204996 104984
rect 205048 104972 205054 104984
rect 213914 104972 213920 104984
rect 205048 104944 213920 104972
rect 205048 104932 205054 104944
rect 213914 104932 213920 104944
rect 213972 104932 213978 104984
rect 258810 104932 258816 104984
rect 258868 104972 258874 104984
rect 265066 104972 265072 104984
rect 258868 104944 265072 104972
rect 258868 104932 258874 104944
rect 265066 104932 265072 104944
rect 265124 104932 265130 104984
rect 174722 104864 174728 104916
rect 174780 104904 174786 104916
rect 214006 104904 214012 104916
rect 174780 104876 214012 104904
rect 174780 104864 174786 104876
rect 214006 104864 214012 104876
rect 214064 104864 214070 104916
rect 260190 104864 260196 104916
rect 260248 104904 260254 104916
rect 264974 104904 264980 104916
rect 260248 104876 264980 104904
rect 260248 104864 260254 104876
rect 264974 104864 264980 104876
rect 265032 104864 265038 104916
rect 231302 104796 231308 104848
rect 231360 104836 231366 104848
rect 243814 104836 243820 104848
rect 231360 104808 243820 104836
rect 231360 104796 231366 104808
rect 243814 104796 243820 104808
rect 243872 104796 243878 104848
rect 254854 104796 254860 104848
rect 254912 104836 254918 104848
rect 257614 104836 257620 104848
rect 254912 104808 257620 104836
rect 254912 104796 254918 104808
rect 257614 104796 257620 104808
rect 257672 104796 257678 104848
rect 282822 104796 282828 104848
rect 282880 104836 282886 104848
rect 310514 104836 310520 104848
rect 282880 104808 310520 104836
rect 282880 104796 282886 104808
rect 310514 104796 310520 104808
rect 310572 104796 310578 104848
rect 281994 104728 282000 104780
rect 282052 104768 282058 104780
rect 292574 104768 292580 104780
rect 282052 104740 292580 104768
rect 282052 104728 282058 104740
rect 292574 104728 292580 104740
rect 292632 104728 292638 104780
rect 231302 103912 231308 103964
rect 231360 103952 231366 103964
rect 234062 103952 234068 103964
rect 231360 103924 234068 103952
rect 231360 103912 231366 103924
rect 234062 103912 234068 103924
rect 234120 103912 234126 103964
rect 191190 103504 191196 103556
rect 191248 103544 191254 103556
rect 213914 103544 213920 103556
rect 191248 103516 213920 103544
rect 191248 103504 191254 103516
rect 213914 103504 213920 103516
rect 213972 103504 213978 103556
rect 233970 103504 233976 103556
rect 234028 103544 234034 103556
rect 264974 103544 264980 103556
rect 234028 103516 264980 103544
rect 234028 103504 234034 103516
rect 264974 103504 264980 103516
rect 265032 103504 265038 103556
rect 282822 103436 282828 103488
rect 282880 103476 282886 103488
rect 289906 103476 289912 103488
rect 282880 103448 289912 103476
rect 282880 103436 282886 103448
rect 289906 103436 289912 103448
rect 289964 103436 289970 103488
rect 231578 103368 231584 103420
rect 231636 103408 231642 103420
rect 240962 103408 240968 103420
rect 231636 103380 240968 103408
rect 231636 103368 231642 103380
rect 240962 103368 240968 103380
rect 241020 103368 241026 103420
rect 282730 103096 282736 103148
rect 282788 103136 282794 103148
rect 288434 103136 288440 103148
rect 282788 103108 288440 103136
rect 282788 103096 282794 103108
rect 288434 103096 288440 103108
rect 288492 103096 288498 103148
rect 230566 102824 230572 102876
rect 230624 102864 230630 102876
rect 232498 102864 232504 102876
rect 230624 102836 232504 102864
rect 230624 102824 230630 102836
rect 232498 102824 232504 102836
rect 232556 102824 232562 102876
rect 173434 102756 173440 102808
rect 173492 102796 173498 102808
rect 191374 102796 191380 102808
rect 173492 102768 191380 102796
rect 173492 102756 173498 102768
rect 191374 102756 191380 102768
rect 191432 102756 191438 102808
rect 192662 102212 192668 102264
rect 192720 102252 192726 102264
rect 213914 102252 213920 102264
rect 192720 102224 213920 102252
rect 192720 102212 192726 102224
rect 213914 102212 213920 102224
rect 213972 102212 213978 102264
rect 171962 102144 171968 102196
rect 172020 102184 172026 102196
rect 214006 102184 214012 102196
rect 172020 102156 214012 102184
rect 172020 102144 172026 102156
rect 214006 102144 214012 102156
rect 214064 102144 214070 102196
rect 250622 102144 250628 102196
rect 250680 102184 250686 102196
rect 264974 102184 264980 102196
rect 250680 102156 264980 102184
rect 250680 102144 250686 102156
rect 264974 102144 264980 102156
rect 265032 102144 265038 102196
rect 231670 102076 231676 102128
rect 231728 102116 231734 102128
rect 254670 102116 254676 102128
rect 231728 102088 254676 102116
rect 231728 102076 231734 102088
rect 254670 102076 254676 102088
rect 254728 102076 254734 102128
rect 282822 102076 282828 102128
rect 282880 102116 282886 102128
rect 309318 102116 309324 102128
rect 282880 102088 309324 102116
rect 282880 102076 282886 102088
rect 309318 102076 309324 102088
rect 309376 102076 309382 102128
rect 231394 102008 231400 102060
rect 231452 102048 231458 102060
rect 239582 102048 239588 102060
rect 231452 102020 239588 102048
rect 231452 102008 231458 102020
rect 239582 102008 239588 102020
rect 239640 102008 239646 102060
rect 260374 100784 260380 100836
rect 260432 100824 260438 100836
rect 265066 100824 265072 100836
rect 260432 100796 265072 100824
rect 260432 100784 260438 100796
rect 265066 100784 265072 100796
rect 265124 100784 265130 100836
rect 177574 100716 177580 100768
rect 177632 100756 177638 100768
rect 213914 100756 213920 100768
rect 177632 100728 213920 100756
rect 177632 100716 177638 100728
rect 213914 100716 213920 100728
rect 213972 100716 213978 100768
rect 246390 100716 246396 100768
rect 246448 100756 246454 100768
rect 264974 100756 264980 100768
rect 246448 100728 264980 100756
rect 246448 100716 246454 100728
rect 264974 100716 264980 100728
rect 265032 100716 265038 100768
rect 231762 100648 231768 100700
rect 231820 100688 231826 100700
rect 261662 100688 261668 100700
rect 231820 100660 261668 100688
rect 231820 100648 231826 100660
rect 261662 100648 261668 100660
rect 261720 100648 261726 100700
rect 281718 100648 281724 100700
rect 281776 100688 281782 100700
rect 295426 100688 295432 100700
rect 281776 100660 295432 100688
rect 281776 100648 281782 100660
rect 295426 100648 295432 100660
rect 295484 100648 295490 100700
rect 231670 100580 231676 100632
rect 231728 100620 231734 100632
rect 245010 100620 245016 100632
rect 231728 100592 245016 100620
rect 231728 100580 231734 100592
rect 245010 100580 245016 100592
rect 245068 100580 245074 100632
rect 167730 99968 167736 100020
rect 167788 100008 167794 100020
rect 211798 100008 211804 100020
rect 167788 99980 211804 100008
rect 167788 99968 167794 99980
rect 211798 99968 211804 99980
rect 211856 99968 211862 100020
rect 211890 99424 211896 99476
rect 211948 99464 211954 99476
rect 214006 99464 214012 99476
rect 211948 99436 214012 99464
rect 211948 99424 211954 99436
rect 214006 99424 214012 99436
rect 214064 99424 214070 99476
rect 169110 99356 169116 99408
rect 169168 99396 169174 99408
rect 213914 99396 213920 99408
rect 169168 99368 213920 99396
rect 169168 99356 169174 99368
rect 213914 99356 213920 99368
rect 213972 99356 213978 99408
rect 245194 99356 245200 99408
rect 245252 99396 245258 99408
rect 264974 99396 264980 99408
rect 245252 99368 264980 99396
rect 245252 99356 245258 99368
rect 264974 99356 264980 99368
rect 265032 99356 265038 99408
rect 231394 99288 231400 99340
rect 231452 99328 231458 99340
rect 246574 99328 246580 99340
rect 231452 99300 246580 99328
rect 231452 99288 231458 99300
rect 246574 99288 246580 99300
rect 246632 99288 246638 99340
rect 231210 99220 231216 99272
rect 231268 99260 231274 99272
rect 243538 99260 243544 99272
rect 231268 99232 243544 99260
rect 231268 99220 231274 99232
rect 243538 99220 243544 99232
rect 243596 99220 243602 99272
rect 253474 98336 253480 98388
rect 253532 98376 253538 98388
rect 256142 98376 256148 98388
rect 253532 98348 256148 98376
rect 253532 98336 253538 98348
rect 256142 98336 256148 98348
rect 256200 98336 256206 98388
rect 211798 98064 211804 98116
rect 211856 98104 211862 98116
rect 214006 98104 214012 98116
rect 211856 98076 214012 98104
rect 211856 98064 211862 98076
rect 214006 98064 214012 98076
rect 214064 98064 214070 98116
rect 167914 97996 167920 98048
rect 167972 98036 167978 98048
rect 213914 98036 213920 98048
rect 167972 98008 213920 98036
rect 167972 97996 167978 98008
rect 213914 97996 213920 98008
rect 213972 97996 213978 98048
rect 256234 97996 256240 98048
rect 256292 98036 256298 98048
rect 264974 98036 264980 98048
rect 256292 98008 264980 98036
rect 256292 97996 256298 98008
rect 264974 97996 264980 98008
rect 265032 97996 265038 98048
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 17218 97968 17224 97980
rect 3476 97940 17224 97968
rect 3476 97928 3482 97940
rect 17218 97928 17224 97940
rect 17276 97928 17282 97980
rect 169570 97928 169576 97980
rect 169628 97968 169634 97980
rect 232774 97968 232780 97980
rect 169628 97940 232780 97968
rect 169628 97928 169634 97940
rect 232774 97928 232780 97940
rect 232832 97928 232838 97980
rect 231210 97860 231216 97912
rect 231268 97900 231274 97912
rect 256050 97900 256056 97912
rect 231268 97872 256056 97900
rect 231268 97860 231274 97872
rect 256050 97860 256056 97872
rect 256108 97860 256114 97912
rect 184658 97248 184664 97300
rect 184716 97288 184722 97300
rect 213270 97288 213276 97300
rect 184716 97260 213276 97288
rect 184716 97248 184722 97260
rect 213270 97248 213276 97260
rect 213328 97248 213334 97300
rect 263134 96704 263140 96756
rect 263192 96744 263198 96756
rect 265066 96744 265072 96756
rect 263192 96716 265072 96744
rect 263192 96704 263198 96716
rect 265066 96704 265072 96716
rect 265124 96704 265130 96756
rect 229002 96676 229008 96688
rect 223684 96648 229008 96676
rect 223684 96076 223712 96648
rect 229002 96636 229008 96648
rect 229060 96636 229066 96688
rect 256142 96636 256148 96688
rect 256200 96676 256206 96688
rect 264974 96676 264980 96688
rect 256200 96648 264980 96676
rect 256200 96636 256206 96648
rect 264974 96636 264980 96648
rect 265032 96636 265038 96688
rect 223666 96024 223672 96076
rect 223724 96024 223730 96076
rect 164970 95956 164976 96008
rect 165028 95996 165034 96008
rect 185670 95996 185676 96008
rect 165028 95968 185676 95996
rect 165028 95956 165034 95968
rect 185670 95956 185676 95968
rect 185728 95956 185734 96008
rect 165890 95888 165896 95940
rect 165948 95928 165954 95940
rect 210602 95928 210608 95940
rect 165948 95900 210608 95928
rect 165948 95888 165954 95900
rect 210602 95888 210608 95900
rect 210660 95888 210666 95940
rect 244274 95616 244280 95668
rect 244332 95656 244338 95668
rect 249794 95656 249800 95668
rect 244332 95628 249800 95656
rect 244332 95616 244338 95628
rect 249794 95616 249800 95628
rect 249852 95616 249858 95668
rect 230474 95480 230480 95532
rect 230532 95520 230538 95532
rect 232498 95520 232504 95532
rect 230532 95492 232504 95520
rect 230532 95480 230538 95492
rect 232498 95480 232504 95492
rect 232556 95480 232562 95532
rect 225598 95276 225604 95328
rect 225656 95316 225662 95328
rect 225656 95288 238754 95316
rect 225656 95276 225662 95288
rect 187970 95208 187976 95260
rect 188028 95248 188034 95260
rect 213914 95248 213920 95260
rect 188028 95220 213920 95248
rect 188028 95208 188034 95220
rect 213914 95208 213920 95220
rect 213972 95208 213978 95260
rect 227070 95208 227076 95260
rect 227128 95248 227134 95260
rect 229094 95248 229100 95260
rect 227128 95220 229100 95248
rect 227128 95208 227134 95220
rect 229094 95208 229100 95220
rect 229152 95208 229158 95260
rect 238726 95248 238754 95288
rect 262674 95248 262680 95260
rect 238726 95220 262680 95248
rect 262674 95208 262680 95220
rect 262732 95208 262738 95260
rect 213362 95140 213368 95192
rect 213420 95180 213426 95192
rect 281534 95180 281540 95192
rect 213420 95152 281540 95180
rect 213420 95140 213426 95152
rect 281534 95140 281540 95152
rect 281592 95140 281598 95192
rect 67450 94528 67456 94580
rect 67508 94568 67514 94580
rect 108298 94568 108304 94580
rect 67508 94540 108304 94568
rect 67508 94528 67514 94540
rect 108298 94528 108304 94540
rect 108356 94528 108362 94580
rect 64690 94460 64696 94512
rect 64748 94500 64754 94512
rect 111058 94500 111064 94512
rect 64748 94472 111064 94500
rect 64748 94460 64754 94472
rect 111058 94460 111064 94472
rect 111116 94460 111122 94512
rect 222930 94460 222936 94512
rect 222988 94500 222994 94512
rect 234246 94500 234252 94512
rect 222988 94472 234252 94500
rect 222988 94460 222994 94472
rect 234246 94460 234252 94472
rect 234304 94460 234310 94512
rect 125410 93916 125416 93968
rect 125468 93956 125474 93968
rect 169202 93956 169208 93968
rect 125468 93928 169208 93956
rect 125468 93916 125474 93928
rect 169202 93916 169208 93928
rect 169260 93916 169266 93968
rect 110138 93848 110144 93900
rect 110196 93888 110202 93900
rect 207842 93888 207848 93900
rect 110196 93860 207848 93888
rect 110196 93848 110202 93860
rect 207842 93848 207848 93860
rect 207900 93848 207906 93900
rect 249794 93780 249800 93832
rect 249852 93820 249858 93832
rect 273990 93820 273996 93832
rect 249852 93792 273996 93820
rect 249852 93780 249858 93792
rect 273990 93780 273996 93792
rect 274048 93780 274054 93832
rect 261478 93712 261484 93764
rect 261536 93752 261542 93764
rect 281718 93752 281724 93764
rect 261536 93724 281724 93752
rect 261536 93712 261542 93724
rect 281718 93712 281724 93724
rect 281776 93712 281782 93764
rect 162762 93168 162768 93220
rect 162820 93208 162826 93220
rect 177390 93208 177396 93220
rect 162820 93180 177396 93208
rect 162820 93168 162826 93180
rect 177390 93168 177396 93180
rect 177448 93168 177454 93220
rect 179046 93168 179052 93220
rect 179104 93208 179110 93220
rect 214558 93208 214564 93220
rect 179104 93180 214564 93208
rect 179104 93168 179110 93180
rect 214558 93168 214564 93180
rect 214616 93168 214622 93220
rect 108114 93100 108120 93152
rect 108172 93140 108178 93152
rect 121454 93140 121460 93152
rect 108172 93112 121460 93140
rect 108172 93100 108178 93112
rect 121454 93100 121460 93112
rect 121512 93100 121518 93152
rect 121730 93100 121736 93152
rect 121788 93140 121794 93152
rect 174630 93140 174636 93152
rect 121788 93112 174636 93140
rect 121788 93100 121794 93112
rect 174630 93100 174636 93112
rect 174688 93100 174694 93152
rect 209130 93100 209136 93152
rect 209188 93140 209194 93152
rect 258994 93140 259000 93152
rect 209188 93112 259000 93140
rect 209188 93100 209194 93112
rect 258994 93100 259000 93112
rect 259052 93100 259058 93152
rect 105722 92488 105728 92540
rect 105780 92528 105786 92540
rect 112438 92528 112444 92540
rect 105780 92500 112444 92528
rect 105780 92488 105786 92500
rect 112438 92488 112444 92500
rect 112496 92488 112502 92540
rect 222838 92488 222844 92540
rect 222896 92528 222902 92540
rect 230014 92528 230020 92540
rect 222896 92500 230020 92528
rect 222896 92488 222902 92500
rect 230014 92488 230020 92500
rect 230072 92488 230078 92540
rect 136082 92420 136088 92472
rect 136140 92460 136146 92472
rect 166350 92460 166356 92472
rect 136140 92432 166356 92460
rect 136140 92420 136146 92432
rect 166350 92420 166356 92432
rect 166408 92420 166414 92472
rect 152090 92352 152096 92404
rect 152148 92392 152154 92404
rect 162762 92392 162768 92404
rect 152148 92364 162768 92392
rect 152148 92352 152154 92364
rect 162762 92352 162768 92364
rect 162820 92352 162826 92404
rect 166442 91808 166448 91860
rect 166500 91848 166506 91860
rect 178862 91848 178868 91860
rect 166500 91820 178868 91848
rect 166500 91808 166506 91820
rect 178862 91808 178868 91820
rect 178920 91808 178926 91860
rect 208394 91808 208400 91860
rect 208452 91848 208458 91860
rect 253474 91848 253480 91860
rect 208452 91820 253480 91848
rect 208452 91808 208458 91820
rect 253474 91808 253480 91820
rect 253532 91808 253538 91860
rect 67358 91740 67364 91792
rect 67416 91780 67422 91792
rect 106918 91780 106924 91792
rect 67416 91752 106924 91780
rect 67416 91740 67422 91752
rect 106918 91740 106924 91752
rect 106976 91740 106982 91792
rect 164878 91740 164884 91792
rect 164936 91780 164942 91792
rect 207658 91780 207664 91792
rect 164936 91752 207664 91780
rect 164936 91740 164942 91752
rect 207658 91740 207664 91752
rect 207716 91740 207722 91792
rect 214558 91740 214564 91792
rect 214616 91780 214622 91792
rect 265802 91780 265808 91792
rect 214616 91752 265808 91780
rect 214616 91740 214622 91752
rect 265802 91740 265808 91752
rect 265860 91740 265866 91792
rect 115474 91128 115480 91180
rect 115532 91168 115538 91180
rect 133138 91168 133144 91180
rect 115532 91140 133144 91168
rect 115532 91128 115538 91140
rect 133138 91128 133144 91140
rect 133196 91128 133202 91180
rect 100018 91060 100024 91112
rect 100076 91100 100082 91112
rect 104250 91100 104256 91112
rect 100076 91072 104256 91100
rect 100076 91060 100082 91072
rect 104250 91060 104256 91072
rect 104308 91060 104314 91112
rect 118050 91060 118056 91112
rect 118108 91100 118114 91112
rect 135898 91100 135904 91112
rect 118108 91072 135904 91100
rect 118108 91060 118114 91072
rect 135898 91060 135904 91072
rect 135956 91060 135962 91112
rect 113450 90992 113456 91044
rect 113508 91032 113514 91044
rect 206278 91032 206284 91044
rect 113508 91004 206284 91032
rect 113508 90992 113514 91004
rect 206278 90992 206284 91004
rect 206336 90992 206342 91044
rect 111610 90924 111616 90976
rect 111668 90964 111674 90976
rect 170582 90964 170588 90976
rect 111668 90936 170588 90964
rect 111668 90924 111674 90936
rect 170582 90924 170588 90936
rect 170640 90924 170646 90976
rect 176102 90380 176108 90432
rect 176160 90420 176166 90432
rect 209314 90420 209320 90432
rect 176160 90392 209320 90420
rect 176160 90380 176166 90392
rect 209314 90380 209320 90392
rect 209372 90380 209378 90432
rect 218698 90380 218704 90432
rect 218756 90420 218762 90432
rect 239674 90420 239680 90432
rect 218756 90392 239680 90420
rect 218756 90380 218762 90392
rect 239674 90380 239680 90392
rect 239732 90380 239738 90432
rect 66162 90312 66168 90364
rect 66220 90352 66226 90364
rect 104158 90352 104164 90364
rect 66220 90324 104164 90352
rect 66220 90312 66226 90324
rect 104158 90312 104164 90324
rect 104216 90312 104222 90364
rect 207658 90312 207664 90364
rect 207716 90352 207722 90364
rect 267274 90352 267280 90364
rect 207716 90324 267280 90352
rect 207716 90312 207722 90324
rect 267274 90312 267280 90324
rect 267332 90312 267338 90364
rect 115566 89632 115572 89684
rect 115624 89672 115630 89684
rect 181622 89672 181628 89684
rect 115624 89644 181628 89672
rect 115624 89632 115630 89644
rect 181622 89632 181628 89644
rect 181680 89632 181686 89684
rect 121178 89564 121184 89616
rect 121236 89604 121242 89616
rect 165890 89604 165896 89616
rect 121236 89576 165896 89604
rect 121236 89564 121242 89576
rect 165890 89564 165896 89576
rect 165948 89564 165954 89616
rect 221458 89020 221464 89072
rect 221516 89060 221522 89072
rect 245102 89060 245108 89072
rect 221516 89032 245108 89060
rect 221516 89020 221522 89032
rect 245102 89020 245108 89032
rect 245160 89020 245166 89072
rect 67542 88952 67548 89004
rect 67600 88992 67606 89004
rect 115198 88992 115204 89004
rect 67600 88964 115204 88992
rect 67600 88952 67606 88964
rect 115198 88952 115204 88964
rect 115256 88952 115262 89004
rect 213270 88952 213276 89004
rect 213328 88992 213334 89004
rect 260466 88992 260472 89004
rect 213328 88964 260472 88992
rect 213328 88952 213334 88964
rect 260466 88952 260472 88964
rect 260524 88952 260530 89004
rect 203518 88340 203524 88392
rect 203576 88380 203582 88392
rect 208394 88380 208400 88392
rect 203576 88352 208400 88380
rect 203576 88340 203582 88352
rect 208394 88340 208400 88352
rect 208452 88340 208458 88392
rect 119706 88272 119712 88324
rect 119764 88312 119770 88324
rect 199470 88312 199476 88324
rect 119764 88284 199476 88312
rect 119764 88272 119770 88284
rect 199470 88272 199476 88284
rect 199528 88272 199534 88324
rect 206278 87660 206284 87712
rect 206336 87700 206342 87712
rect 229830 87700 229836 87712
rect 206336 87672 229836 87700
rect 206336 87660 206342 87672
rect 229830 87660 229836 87672
rect 229888 87660 229894 87712
rect 165062 87592 165068 87644
rect 165120 87632 165126 87644
rect 203610 87632 203616 87644
rect 165120 87604 203616 87632
rect 165120 87592 165126 87604
rect 203610 87592 203616 87604
rect 203668 87592 203674 87644
rect 214742 87592 214748 87644
rect 214800 87632 214806 87644
rect 247954 87632 247960 87644
rect 214800 87604 247960 87632
rect 214800 87592 214806 87604
rect 247954 87592 247960 87604
rect 248012 87592 248018 87644
rect 93210 86912 93216 86964
rect 93268 86952 93274 86964
rect 167822 86952 167828 86964
rect 93268 86924 167828 86952
rect 93268 86912 93274 86924
rect 167822 86912 167828 86924
rect 167880 86912 167886 86964
rect 151538 86844 151544 86896
rect 151596 86884 151602 86896
rect 166258 86884 166264 86896
rect 151596 86856 166264 86884
rect 151596 86844 151602 86856
rect 166258 86844 166264 86856
rect 166316 86844 166322 86896
rect 220078 86300 220084 86352
rect 220136 86340 220142 86352
rect 254854 86340 254860 86352
rect 220136 86312 254860 86340
rect 220136 86300 220142 86312
rect 254854 86300 254860 86312
rect 254912 86300 254918 86352
rect 184290 86232 184296 86284
rect 184348 86272 184354 86284
rect 235534 86272 235540 86284
rect 184348 86244 235540 86272
rect 184348 86232 184354 86244
rect 235534 86232 235540 86244
rect 235592 86232 235598 86284
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 11698 85524 11704 85536
rect 3200 85496 11704 85524
rect 3200 85484 3206 85496
rect 11698 85484 11704 85496
rect 11756 85484 11762 85536
rect 105538 85484 105544 85536
rect 105596 85524 105602 85536
rect 205082 85524 205088 85536
rect 105596 85496 205088 85524
rect 105596 85484 105602 85496
rect 205082 85484 205088 85496
rect 205140 85484 205146 85536
rect 126514 85416 126520 85468
rect 126572 85456 126578 85468
rect 196802 85456 196808 85468
rect 126572 85428 196808 85456
rect 126572 85416 126578 85428
rect 196802 85416 196808 85428
rect 196860 85416 196866 85468
rect 215938 84872 215944 84924
rect 215996 84912 216002 84924
rect 231302 84912 231308 84924
rect 215996 84884 231308 84912
rect 215996 84872 216002 84884
rect 231302 84872 231308 84884
rect 231360 84872 231366 84924
rect 226978 84804 226984 84856
rect 227036 84844 227042 84856
rect 245194 84844 245200 84856
rect 227036 84816 245200 84844
rect 227036 84804 227042 84816
rect 245194 84804 245200 84816
rect 245252 84804 245258 84856
rect 96522 84124 96528 84176
rect 96580 84164 96586 84176
rect 182910 84164 182916 84176
rect 96580 84136 182916 84164
rect 96580 84124 96586 84136
rect 182910 84124 182916 84136
rect 182968 84124 182974 84176
rect 97810 84056 97816 84108
rect 97868 84096 97874 84108
rect 173342 84096 173348 84108
rect 97868 84068 173348 84096
rect 97868 84056 97874 84068
rect 173342 84056 173348 84068
rect 173400 84056 173406 84108
rect 195238 83512 195244 83564
rect 195296 83552 195302 83564
rect 232866 83552 232872 83564
rect 195296 83524 232872 83552
rect 195296 83512 195302 83524
rect 232866 83512 232872 83524
rect 232924 83512 232930 83564
rect 178678 83444 178684 83496
rect 178736 83484 178742 83496
rect 281534 83484 281540 83496
rect 178736 83456 281540 83484
rect 178736 83444 178742 83456
rect 281534 83444 281540 83456
rect 281592 83444 281598 83496
rect 100570 82764 100576 82816
rect 100628 82804 100634 82816
rect 187050 82804 187056 82816
rect 100628 82776 187056 82804
rect 100628 82764 100634 82776
rect 187050 82764 187056 82776
rect 187108 82764 187114 82816
rect 107562 82696 107568 82748
rect 107620 82736 107626 82748
rect 184382 82736 184388 82748
rect 107620 82708 184388 82736
rect 107620 82696 107626 82708
rect 184382 82696 184388 82708
rect 184440 82696 184446 82748
rect 95142 81336 95148 81388
rect 95200 81376 95206 81388
rect 202322 81376 202328 81388
rect 95200 81348 202328 81376
rect 95200 81336 95206 81348
rect 202322 81336 202328 81348
rect 202380 81336 202386 81388
rect 129642 81268 129648 81320
rect 129700 81308 129706 81320
rect 177482 81308 177488 81320
rect 129700 81280 177488 81308
rect 129700 81268 129706 81280
rect 177482 81268 177488 81280
rect 177540 81268 177546 81320
rect 133782 79976 133788 80028
rect 133840 80016 133846 80028
rect 216030 80016 216036 80028
rect 133840 79988 216036 80016
rect 133840 79976 133846 79988
rect 216030 79976 216036 79988
rect 216088 79976 216094 80028
rect 117222 79908 117228 79960
rect 117280 79948 117286 79960
rect 173434 79948 173440 79960
rect 117280 79920 173440 79948
rect 117280 79908 117286 79920
rect 173434 79908 173440 79920
rect 173492 79908 173498 79960
rect 118510 78616 118516 78668
rect 118568 78656 118574 78668
rect 169202 78656 169208 78668
rect 118568 78628 169208 78656
rect 118568 78616 118574 78628
rect 169202 78616 169208 78628
rect 169260 78616 169266 78668
rect 151630 78548 151636 78600
rect 151688 78588 151694 78600
rect 165062 78588 165068 78600
rect 151688 78560 165068 78588
rect 151688 78548 151694 78560
rect 165062 78548 165068 78560
rect 165120 78548 165126 78600
rect 174538 77936 174544 77988
rect 174596 77976 174602 77988
rect 241514 77976 241520 77988
rect 174596 77948 241520 77976
rect 174596 77936 174602 77948
rect 241514 77936 241520 77948
rect 241572 77936 241578 77988
rect 91002 77188 91008 77240
rect 91060 77228 91066 77240
rect 174722 77228 174728 77240
rect 91060 77200 174728 77228
rect 91060 77188 91066 77200
rect 174722 77188 174728 77200
rect 174780 77188 174786 77240
rect 126238 76508 126244 76560
rect 126296 76548 126302 76560
rect 265710 76548 265716 76560
rect 126296 76520 265716 76548
rect 126296 76508 126302 76520
rect 265710 76508 265716 76520
rect 265768 76508 265774 76560
rect 104250 75828 104256 75880
rect 104308 75868 104314 75880
rect 170490 75868 170496 75880
rect 104308 75840 170496 75868
rect 104308 75828 104314 75840
rect 170490 75828 170496 75840
rect 170548 75828 170554 75880
rect 119982 75148 119988 75200
rect 120040 75188 120046 75200
rect 254762 75188 254768 75200
rect 120040 75160 254768 75188
rect 120040 75148 120046 75160
rect 254762 75148 254768 75160
rect 254820 75148 254826 75200
rect 124858 74468 124864 74520
rect 124916 74508 124922 74520
rect 206462 74508 206468 74520
rect 124916 74480 206468 74508
rect 124916 74468 124922 74480
rect 206462 74468 206468 74480
rect 206520 74468 206526 74520
rect 114278 74400 114284 74452
rect 114336 74440 114342 74452
rect 164878 74440 164884 74452
rect 114336 74412 164884 74440
rect 114336 74400 114342 74412
rect 164878 74400 164884 74412
rect 164936 74400 164942 74452
rect 117130 73108 117136 73160
rect 117188 73148 117194 73160
rect 162118 73148 162124 73160
rect 117188 73120 162124 73148
rect 117188 73108 117194 73120
rect 162118 73108 162124 73120
rect 162176 73108 162182 73160
rect 151722 73040 151728 73092
rect 151780 73080 151786 73092
rect 181530 73080 181536 73092
rect 151780 73052 181536 73080
rect 151780 73040 151786 73052
rect 181530 73040 181536 73052
rect 181588 73040 181594 73092
rect 3418 71680 3424 71732
rect 3476 71720 3482 71732
rect 39298 71720 39304 71732
rect 3476 71692 39304 71720
rect 3476 71680 3482 71692
rect 39298 71680 39304 71692
rect 39356 71680 39362 71732
rect 64782 71680 64788 71732
rect 64840 71720 64846 71732
rect 204990 71720 204996 71732
rect 64840 71692 204996 71720
rect 64840 71680 64846 71692
rect 204990 71680 204996 71692
rect 205048 71680 205054 71732
rect 119890 71612 119896 71664
rect 119948 71652 119954 71664
rect 167730 71652 167736 71664
rect 119948 71624 167736 71652
rect 119948 71612 119954 71624
rect 167730 71612 167736 71624
rect 167788 71612 167794 71664
rect 102042 70320 102048 70372
rect 102100 70360 102106 70372
rect 179046 70360 179052 70372
rect 102100 70332 179052 70360
rect 102100 70320 102106 70332
rect 179046 70320 179052 70332
rect 179104 70320 179110 70372
rect 131022 70252 131028 70304
rect 131080 70292 131086 70304
rect 173158 70292 173164 70304
rect 131080 70264 173164 70292
rect 131080 70252 131086 70264
rect 173158 70252 173164 70264
rect 173216 70252 173222 70304
rect 122742 68960 122748 69012
rect 122800 69000 122806 69012
rect 210418 69000 210424 69012
rect 122800 68972 210424 69000
rect 122800 68960 122806 68972
rect 210418 68960 210424 68972
rect 210476 68960 210482 69012
rect 130378 68280 130384 68332
rect 130436 68320 130442 68332
rect 169754 68320 169760 68332
rect 130436 68292 169760 68320
rect 130436 68280 130442 68292
rect 169754 68280 169760 68292
rect 169812 68280 169818 68332
rect 110230 67532 110236 67584
rect 110288 67572 110294 67584
rect 176102 67572 176108 67584
rect 110288 67544 176108 67572
rect 110288 67532 110294 67544
rect 176102 67532 176108 67544
rect 176160 67532 176166 67584
rect 133138 67464 133144 67516
rect 133196 67504 133202 67516
rect 166442 67504 166448 67516
rect 133196 67476 166448 67504
rect 133196 67464 133202 67476
rect 166442 67464 166448 67476
rect 166500 67464 166506 67516
rect 104710 66172 104716 66224
rect 104768 66212 104774 66224
rect 180150 66212 180156 66224
rect 104768 66184 180156 66212
rect 104768 66172 104774 66184
rect 180150 66172 180156 66184
rect 180208 66172 180214 66224
rect 124030 66104 124036 66156
rect 124088 66144 124094 66156
rect 195330 66144 195336 66156
rect 124088 66116 195336 66144
rect 124088 66104 124094 66116
rect 195330 66104 195336 66116
rect 195388 66104 195394 66156
rect 103330 64812 103336 64864
rect 103388 64852 103394 64864
rect 200850 64852 200856 64864
rect 103388 64824 200856 64852
rect 103388 64812 103394 64824
rect 200850 64812 200856 64824
rect 200908 64812 200914 64864
rect 122098 64744 122104 64796
rect 122156 64784 122162 64796
rect 192662 64784 192668 64796
rect 122156 64756 192668 64784
rect 122156 64744 122162 64756
rect 192662 64744 192668 64756
rect 192720 64744 192726 64796
rect 228450 64132 228456 64184
rect 228508 64172 228514 64184
rect 267734 64172 267740 64184
rect 228508 64144 267740 64172
rect 228508 64132 228514 64144
rect 267734 64132 267740 64144
rect 267792 64132 267798 64184
rect 111702 63452 111708 63504
rect 111760 63492 111766 63504
rect 199378 63492 199384 63504
rect 111760 63464 199384 63492
rect 111760 63452 111766 63464
rect 199378 63452 199384 63464
rect 199436 63452 199442 63504
rect 93762 62772 93768 62824
rect 93820 62812 93826 62824
rect 267090 62812 267096 62824
rect 93820 62784 267096 62812
rect 93820 62772 93826 62784
rect 267090 62772 267096 62784
rect 267148 62772 267154 62824
rect 121362 62024 121368 62076
rect 121420 62064 121426 62076
rect 186958 62064 186964 62076
rect 121420 62036 186964 62064
rect 121420 62024 121426 62036
rect 186958 62024 186964 62036
rect 187016 62024 187022 62076
rect 77202 61344 77208 61396
rect 77260 61384 77266 61396
rect 253382 61384 253388 61396
rect 77260 61356 253388 61384
rect 77260 61344 77266 61356
rect 253382 61344 253388 61356
rect 253440 61344 253446 61396
rect 107562 60052 107568 60104
rect 107620 60092 107626 60104
rect 229738 60092 229744 60104
rect 107620 60064 229744 60092
rect 107620 60052 107626 60064
rect 229738 60052 229744 60064
rect 229796 60052 229802 60104
rect 79962 59984 79968 60036
rect 80020 60024 80026 60036
rect 251910 60024 251916 60036
rect 80020 59996 251916 60024
rect 80020 59984 80026 59996
rect 251910 59984 251916 59996
rect 251968 59984 251974 60036
rect 3050 59304 3056 59356
rect 3108 59344 3114 59356
rect 33778 59344 33784 59356
rect 3108 59316 33784 59344
rect 3108 59304 3114 59316
rect 33778 59304 33784 59316
rect 33836 59304 33842 59356
rect 112438 59304 112444 59356
rect 112496 59344 112502 59356
rect 191282 59344 191288 59356
rect 112496 59316 191288 59344
rect 112496 59304 112502 59316
rect 191282 59304 191288 59316
rect 191340 59304 191346 59356
rect 86862 58624 86868 58676
rect 86920 58664 86926 58676
rect 250438 58664 250444 58676
rect 86920 58636 250444 58664
rect 86920 58624 86926 58636
rect 250438 58624 250444 58636
rect 250496 58624 250502 58676
rect 99190 57876 99196 57928
rect 99248 57916 99254 57928
rect 178770 57916 178776 57928
rect 99248 57888 178776 57916
rect 99248 57876 99254 57888
rect 178770 57876 178776 57888
rect 178828 57876 178834 57928
rect 100662 57196 100668 57248
rect 100720 57236 100726 57248
rect 236730 57236 236736 57248
rect 100720 57208 236736 57236
rect 100720 57196 100726 57208
rect 236730 57196 236736 57208
rect 236788 57196 236794 57248
rect 115658 56516 115664 56568
rect 115716 56556 115722 56568
rect 216122 56556 216128 56568
rect 115716 56528 216128 56556
rect 115716 56516 115722 56528
rect 216122 56516 216128 56528
rect 216180 56516 216186 56568
rect 91002 55836 91008 55888
rect 91060 55876 91066 55888
rect 243722 55876 243728 55888
rect 91060 55848 243728 55876
rect 91060 55836 91066 55848
rect 243722 55836 243728 55848
rect 243780 55836 243786 55888
rect 110322 55156 110328 55208
rect 110380 55196 110386 55208
rect 206370 55196 206376 55208
rect 110380 55168 206376 55196
rect 110380 55156 110386 55168
rect 206370 55156 206376 55168
rect 206428 55156 206434 55208
rect 97902 54476 97908 54528
rect 97960 54516 97966 54528
rect 242250 54516 242256 54528
rect 97960 54488 242256 54516
rect 97960 54476 97966 54488
rect 242250 54476 242256 54488
rect 242308 54476 242314 54528
rect 85482 53728 85488 53780
rect 85540 53768 85546 53780
rect 214650 53768 214656 53780
rect 85540 53740 214656 53768
rect 85540 53728 85546 53740
rect 214650 53728 214656 53740
rect 214708 53728 214714 53780
rect 102042 53048 102048 53100
rect 102100 53088 102106 53100
rect 257430 53088 257436 53100
rect 102100 53060 257436 53088
rect 102100 53048 102106 53060
rect 257430 53048 257436 53060
rect 257488 53048 257494 53100
rect 86770 52368 86776 52420
rect 86828 52408 86834 52420
rect 211798 52408 211804 52420
rect 86828 52380 211804 52408
rect 86828 52368 86834 52380
rect 211798 52368 211804 52380
rect 211856 52368 211862 52420
rect 124122 52300 124128 52352
rect 124180 52340 124186 52352
rect 176010 52340 176016 52352
rect 124180 52312 176016 52340
rect 124180 52300 124186 52312
rect 176010 52300 176016 52312
rect 176068 52300 176074 52352
rect 95050 51008 95056 51060
rect 95108 51048 95114 51060
rect 210510 51048 210516 51060
rect 95108 51020 210516 51048
rect 95108 51008 95114 51020
rect 210510 51008 210516 51020
rect 210568 51008 210574 51060
rect 111702 50328 111708 50380
rect 111760 50368 111766 50380
rect 255958 50368 255964 50380
rect 111760 50340 255964 50368
rect 111760 50328 111766 50340
rect 255958 50328 255964 50340
rect 256016 50328 256022 50380
rect 70302 48968 70308 49020
rect 70360 49008 70366 49020
rect 260190 49008 260196 49020
rect 70360 48980 260196 49008
rect 70360 48968 70366 48980
rect 260190 48968 260196 48980
rect 260248 48968 260254 49020
rect 115842 47608 115848 47660
rect 115900 47648 115906 47660
rect 244918 47648 244924 47660
rect 115900 47620 244924 47648
rect 115900 47608 115906 47620
rect 244918 47608 244924 47620
rect 244976 47608 244982 47660
rect 31662 47540 31668 47592
rect 31720 47580 31726 47592
rect 254578 47580 254584 47592
rect 31720 47552 254584 47580
rect 31720 47540 31726 47552
rect 254578 47540 254584 47552
rect 254636 47540 254642 47592
rect 98638 46248 98644 46300
rect 98696 46288 98702 46300
rect 207658 46288 207664 46300
rect 98696 46260 207664 46288
rect 98696 46248 98702 46260
rect 207658 46248 207664 46260
rect 207716 46248 207722 46300
rect 22002 46180 22008 46232
rect 22060 46220 22066 46232
rect 245010 46220 245016 46232
rect 22060 46192 245016 46220
rect 22060 46180 22066 46192
rect 245010 46180 245016 46192
rect 245068 46180 245074 46232
rect 3418 45500 3424 45552
rect 3476 45540 3482 45552
rect 36538 45540 36544 45552
rect 3476 45512 36544 45540
rect 3476 45500 3482 45512
rect 36538 45500 36544 45512
rect 36596 45500 36602 45552
rect 66162 44888 66168 44940
rect 66220 44928 66226 44940
rect 258810 44928 258816 44940
rect 66220 44900 258816 44928
rect 66220 44888 66226 44900
rect 258810 44888 258816 44900
rect 258868 44888 258874 44940
rect 50982 44820 50988 44872
rect 51040 44860 51046 44872
rect 249794 44860 249800 44872
rect 51040 44832 249800 44860
rect 51040 44820 51046 44832
rect 249794 44820 249800 44832
rect 249852 44820 249858 44872
rect 124858 43460 124864 43512
rect 124916 43500 124922 43512
rect 209222 43500 209228 43512
rect 124916 43472 209228 43500
rect 124916 43460 124922 43472
rect 209222 43460 209228 43472
rect 209280 43460 209286 43512
rect 217226 43460 217232 43512
rect 217284 43500 217290 43512
rect 259454 43500 259460 43512
rect 217284 43472 259460 43500
rect 217284 43460 217290 43472
rect 259454 43460 259460 43472
rect 259512 43460 259518 43512
rect 34422 43392 34428 43444
rect 34480 43432 34486 43444
rect 246390 43432 246396 43444
rect 34480 43404 246396 43432
rect 34480 43392 34486 43404
rect 246390 43392 246396 43404
rect 246448 43392 246454 43444
rect 122742 42100 122748 42152
rect 122800 42140 122806 42152
rect 213270 42140 213276 42152
rect 122800 42112 213276 42140
rect 122800 42100 122806 42112
rect 213270 42100 213276 42112
rect 213328 42100 213334 42152
rect 45462 42032 45468 42084
rect 45520 42072 45526 42084
rect 239490 42072 239496 42084
rect 45520 42044 239496 42072
rect 45520 42032 45526 42044
rect 239490 42032 239496 42044
rect 239548 42032 239554 42084
rect 85482 40740 85488 40792
rect 85540 40780 85546 40792
rect 260098 40780 260104 40792
rect 85540 40752 260104 40780
rect 85540 40740 85546 40752
rect 260098 40740 260104 40752
rect 260156 40740 260162 40792
rect 46842 40672 46848 40724
rect 46900 40712 46906 40724
rect 235350 40712 235356 40724
rect 46900 40684 235356 40712
rect 46900 40672 46906 40684
rect 235350 40672 235356 40684
rect 235408 40672 235414 40724
rect 99282 37952 99288 38004
rect 99340 37992 99346 38004
rect 184290 37992 184296 38004
rect 99340 37964 184296 37992
rect 99340 37952 99346 37964
rect 184290 37952 184296 37964
rect 184348 37952 184354 38004
rect 49602 37884 49608 37936
rect 49660 37924 49666 37936
rect 253290 37924 253296 37936
rect 49660 37896 253296 37924
rect 49660 37884 49666 37896
rect 253290 37884 253296 37896
rect 253348 37884 253354 37936
rect 200758 36592 200764 36644
rect 200816 36632 200822 36644
rect 269114 36632 269120 36644
rect 200816 36604 269120 36632
rect 200816 36592 200822 36604
rect 269114 36592 269120 36604
rect 269172 36592 269178 36644
rect 56502 36524 56508 36576
rect 56560 36564 56566 36576
rect 242158 36564 242164 36576
rect 56560 36536 242164 36564
rect 56560 36524 56566 36536
rect 242158 36524 242164 36536
rect 242216 36524 242222 36576
rect 4062 35232 4068 35284
rect 4120 35272 4126 35284
rect 185578 35272 185584 35284
rect 4120 35244 185584 35272
rect 4120 35232 4126 35244
rect 185578 35232 185584 35244
rect 185636 35232 185642 35284
rect 53558 35164 53564 35216
rect 53616 35204 53622 35216
rect 251818 35204 251824 35216
rect 53616 35176 251824 35204
rect 53616 35164 53622 35176
rect 251818 35164 251824 35176
rect 251876 35164 251882 35216
rect 61930 33804 61936 33856
rect 61988 33844 61994 33856
rect 267182 33844 267188 33856
rect 61988 33816 267188 33844
rect 61988 33804 61994 33816
rect 267182 33804 267188 33816
rect 267240 33804 267246 33856
rect 53742 33736 53748 33788
rect 53800 33776 53806 33788
rect 278774 33776 278780 33788
rect 53800 33748 278780 33776
rect 53800 33736 53806 33748
rect 278774 33736 278780 33748
rect 278832 33736 278838 33788
rect 3142 33056 3148 33108
rect 3200 33096 3206 33108
rect 35158 33096 35164 33108
rect 3200 33068 35164 33096
rect 3200 33056 3206 33068
rect 35158 33056 35164 33068
rect 35216 33056 35222 33108
rect 124122 32444 124128 32496
rect 124180 32484 124186 32496
rect 258718 32484 258724 32496
rect 124180 32456 258724 32484
rect 124180 32444 124186 32456
rect 258718 32444 258724 32456
rect 258776 32444 258782 32496
rect 44082 32376 44088 32428
rect 44140 32416 44146 32428
rect 296714 32416 296720 32428
rect 44140 32388 296720 32416
rect 44140 32376 44146 32388
rect 296714 32376 296720 32388
rect 296772 32376 296778 32428
rect 54938 31084 54944 31136
rect 54996 31124 55002 31136
rect 218698 31124 218704 31136
rect 54996 31096 218704 31124
rect 54996 31084 55002 31096
rect 218698 31084 218704 31096
rect 218756 31084 218762 31136
rect 37090 31016 37096 31068
rect 37148 31056 37154 31068
rect 243630 31056 243636 31068
rect 37148 31028 243636 31056
rect 37148 31016 37154 31028
rect 243630 31016 243636 31028
rect 243688 31016 243694 31068
rect 59170 29656 59176 29708
rect 59228 29696 59234 29708
rect 233970 29696 233976 29708
rect 59228 29668 233976 29696
rect 59228 29656 59234 29668
rect 233970 29656 233976 29668
rect 234028 29656 234034 29708
rect 62022 29588 62028 29640
rect 62080 29628 62086 29640
rect 324406 29628 324412 29640
rect 62080 29600 324412 29628
rect 62080 29588 62086 29600
rect 324406 29588 324412 29600
rect 324464 29588 324470 29640
rect 84102 28296 84108 28348
rect 84160 28336 84166 28348
rect 209130 28336 209136 28348
rect 84160 28308 209136 28336
rect 84160 28296 84166 28308
rect 209130 28296 209136 28308
rect 209188 28296 209194 28348
rect 1394 28228 1400 28280
rect 1452 28268 1458 28280
rect 231210 28268 231216 28280
rect 1452 28240 231216 28268
rect 1452 28228 1458 28240
rect 231210 28228 231216 28240
rect 231268 28228 231274 28280
rect 90358 26868 90364 26920
rect 90416 26908 90422 26920
rect 221458 26908 221464 26920
rect 90416 26880 221464 26908
rect 90416 26868 90422 26880
rect 221458 26868 221464 26880
rect 221516 26868 221522 26920
rect 113082 25508 113088 25560
rect 113140 25548 113146 25560
rect 235258 25548 235264 25560
rect 113140 25520 235264 25548
rect 113140 25508 113146 25520
rect 235258 25508 235264 25520
rect 235316 25508 235322 25560
rect 111610 24080 111616 24132
rect 111668 24120 111674 24132
rect 262858 24120 262864 24132
rect 111668 24092 262864 24120
rect 111668 24080 111674 24092
rect 262858 24080 262864 24092
rect 262916 24080 262922 24132
rect 123478 22788 123484 22840
rect 123536 22828 123542 22840
rect 160738 22828 160744 22840
rect 123536 22800 160744 22828
rect 123536 22788 123542 22800
rect 160738 22788 160744 22800
rect 160796 22788 160802 22840
rect 39942 22720 39948 22772
rect 40000 22760 40006 22772
rect 232682 22760 232688 22772
rect 40000 22732 232688 22760
rect 40000 22720 40006 22732
rect 232682 22720 232688 22732
rect 232740 22720 232746 22772
rect 188338 21428 188344 21480
rect 188396 21468 188402 21480
rect 269114 21468 269120 21480
rect 188396 21440 269120 21468
rect 188396 21428 188402 21440
rect 269114 21428 269120 21440
rect 269172 21428 269178 21480
rect 92382 21360 92388 21412
rect 92440 21400 92446 21412
rect 204898 21400 204904 21412
rect 92440 21372 204904 21400
rect 92440 21360 92446 21372
rect 204898 21360 204904 21372
rect 204956 21360 204962 21412
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 51718 20652 51724 20664
rect 3476 20624 51724 20652
rect 3476 20612 3482 20624
rect 51718 20612 51724 20624
rect 51776 20612 51782 20664
rect 48222 19932 48228 19984
rect 48280 19972 48286 19984
rect 289814 19972 289820 19984
rect 48280 19944 289820 19972
rect 48280 19932 48286 19944
rect 289814 19932 289820 19944
rect 289872 19932 289878 19984
rect 103422 18640 103428 18692
rect 103480 18680 103486 18692
rect 222930 18680 222936 18692
rect 103480 18652 222936 18680
rect 103480 18640 103486 18652
rect 222930 18640 222936 18652
rect 222988 18640 222994 18692
rect 55122 18572 55128 18624
rect 55180 18612 55186 18624
rect 310514 18612 310520 18624
rect 55180 18584 310520 18612
rect 55180 18572 55186 18584
rect 310514 18572 310520 18584
rect 310572 18572 310578 18624
rect 209038 17280 209044 17332
rect 209096 17320 209102 17332
rect 302234 17320 302240 17332
rect 209096 17292 302240 17320
rect 209096 17280 209102 17292
rect 302234 17280 302240 17292
rect 302292 17280 302298 17332
rect 81342 17212 81348 17264
rect 81400 17252 81406 17264
rect 240778 17252 240784 17264
rect 81400 17224 240784 17252
rect 81400 17212 81406 17224
rect 240778 17212 240784 17224
rect 240836 17212 240842 17264
rect 181438 15920 181444 15972
rect 181496 15960 181502 15972
rect 269758 15960 269764 15972
rect 181496 15932 269764 15960
rect 181496 15920 181502 15932
rect 269758 15920 269764 15932
rect 269816 15920 269822 15972
rect 110322 15852 110328 15904
rect 110380 15892 110386 15904
rect 239398 15892 239404 15904
rect 110380 15864 239404 15892
rect 110380 15852 110386 15864
rect 239398 15852 239404 15864
rect 239456 15852 239462 15904
rect 135254 14696 135260 14748
rect 135312 14736 135318 14748
rect 136450 14736 136456 14748
rect 135312 14708 136456 14736
rect 135312 14696 135318 14708
rect 136450 14696 136456 14708
rect 136508 14696 136514 14748
rect 121086 14492 121092 14544
rect 121144 14532 121150 14544
rect 203518 14532 203524 14544
rect 121144 14504 203524 14532
rect 121144 14492 121150 14504
rect 203518 14492 203524 14504
rect 203576 14492 203582 14544
rect 12158 14424 12164 14476
rect 12216 14464 12222 14476
rect 226978 14464 226984 14476
rect 12216 14436 226984 14464
rect 12216 14424 12222 14436
rect 226978 14424 226984 14436
rect 227036 14424 227042 14476
rect 118602 13132 118608 13184
rect 118660 13172 118666 13184
rect 231118 13172 231124 13184
rect 118660 13144 231124 13172
rect 118660 13132 118666 13144
rect 231118 13132 231124 13144
rect 231176 13132 231182 13184
rect 60642 13064 60648 13116
rect 60700 13104 60706 13116
rect 253198 13104 253204 13116
rect 60700 13076 253204 13104
rect 60700 13064 60706 13076
rect 253198 13064 253204 13076
rect 253256 13064 253262 13116
rect 197998 11772 198004 11824
rect 198056 11812 198062 11824
rect 245194 11812 245200 11824
rect 198056 11784 245200 11812
rect 198056 11772 198062 11784
rect 245194 11772 245200 11784
rect 245252 11772 245258 11824
rect 96246 11704 96252 11756
rect 96304 11744 96310 11756
rect 215938 11744 215944 11756
rect 96304 11716 215944 11744
rect 96304 11704 96310 11716
rect 215938 11704 215944 11716
rect 215996 11704 216002 11756
rect 259454 11704 259460 11756
rect 259512 11744 259518 11756
rect 260650 11744 260656 11756
rect 259512 11716 260656 11744
rect 259512 11704 259518 11716
rect 260650 11704 260656 11716
rect 260708 11704 260714 11756
rect 307846 11704 307852 11756
rect 307904 11744 307910 11756
rect 309042 11744 309048 11756
rect 307904 11716 309048 11744
rect 307904 11704 307910 11716
rect 309042 11704 309048 11716
rect 309100 11704 309106 11756
rect 332686 11704 332692 11756
rect 332744 11744 332750 11756
rect 333882 11744 333888 11756
rect 332744 11716 333888 11744
rect 332744 11704 332750 11716
rect 333882 11704 333888 11716
rect 333940 11704 333946 11756
rect 114462 10344 114468 10396
rect 114520 10384 114526 10396
rect 220078 10384 220084 10396
rect 114520 10356 220084 10384
rect 114520 10344 114526 10356
rect 220078 10344 220084 10356
rect 220136 10344 220142 10396
rect 9582 10276 9588 10328
rect 9640 10316 9646 10328
rect 180058 10316 180064 10328
rect 9640 10288 180064 10316
rect 9640 10276 9646 10288
rect 180058 10276 180064 10288
rect 180116 10276 180122 10328
rect 184198 10276 184204 10328
rect 184256 10316 184262 10328
rect 244090 10316 244096 10328
rect 184256 10288 244096 10316
rect 184256 10276 184262 10288
rect 244090 10276 244096 10288
rect 244148 10276 244154 10328
rect 77386 8984 77392 9036
rect 77444 9024 77450 9036
rect 98638 9024 98644 9036
rect 77444 8996 98644 9024
rect 77444 8984 77450 8996
rect 98638 8984 98644 8996
rect 98696 8984 98702 9036
rect 177298 8984 177304 9036
rect 177356 9024 177362 9036
rect 242894 9024 242900 9036
rect 177356 8996 242900 9024
rect 177356 8984 177362 8996
rect 242894 8984 242900 8996
rect 242952 8984 242958 9036
rect 97810 8916 97816 8968
rect 97868 8956 97874 8968
rect 264238 8956 264244 8968
rect 97868 8928 264244 8956
rect 97868 8916 97874 8928
rect 264238 8916 264244 8928
rect 264296 8916 264302 8968
rect 224218 7556 224224 7608
rect 224276 7596 224282 7608
rect 253474 7596 253480 7608
rect 224276 7568 253480 7596
rect 224276 7556 224282 7568
rect 253474 7556 253480 7568
rect 253532 7556 253538 7608
rect 71498 6196 71504 6248
rect 71556 6236 71562 6248
rect 233878 6236 233884 6248
rect 71556 6208 233884 6236
rect 71556 6196 71562 6208
rect 233878 6196 233884 6208
rect 233936 6196 233942 6248
rect 47854 6128 47860 6180
rect 47912 6168 47918 6180
rect 228358 6168 228364 6180
rect 47912 6140 228364 6168
rect 47912 6128 47918 6140
rect 228358 6128 228364 6140
rect 228416 6128 228422 6180
rect 238018 6128 238024 6180
rect 238076 6168 238082 6180
rect 267734 6168 267740 6180
rect 238076 6140 267740 6168
rect 238076 6128 238082 6140
rect 267734 6128 267740 6140
rect 267792 6128 267798 6180
rect 340966 6128 340972 6180
rect 341024 6168 341030 6180
rect 349154 6168 349160 6180
rect 341024 6140 349160 6168
rect 341024 6128 341030 6140
rect 349154 6128 349160 6140
rect 349212 6128 349218 6180
rect 304350 5516 304356 5568
rect 304408 5556 304414 5568
rect 305086 5556 305092 5568
rect 304408 5528 305092 5556
rect 304408 5516 304414 5528
rect 305086 5516 305092 5528
rect 305144 5516 305150 5568
rect 95142 4836 95148 4888
rect 95200 4876 95206 4888
rect 266998 4876 267004 4888
rect 95200 4848 267004 4876
rect 95200 4836 95206 4848
rect 266998 4836 267004 4848
rect 267056 4836 267062 4888
rect 20622 4768 20628 4820
rect 20680 4808 20686 4820
rect 228450 4808 228456 4820
rect 20680 4780 228456 4808
rect 20680 4768 20686 4780
rect 228450 4768 228456 4780
rect 228508 4768 228514 4820
rect 318058 4768 318064 4820
rect 318116 4808 318122 4820
rect 329190 4808 329196 4820
rect 318116 4780 329196 4808
rect 318116 4768 318122 4780
rect 329190 4768 329196 4780
rect 329248 4768 329254 4820
rect 232498 4156 232504 4208
rect 232556 4196 232562 4208
rect 235810 4196 235816 4208
rect 232556 4168 235816 4196
rect 232556 4156 232562 4168
rect 235810 4156 235816 4168
rect 235868 4156 235874 4208
rect 296070 4088 296076 4140
rect 296128 4128 296134 4140
rect 298094 4128 298100 4140
rect 296128 4100 298100 4128
rect 296128 4088 296134 4100
rect 298094 4088 298100 4100
rect 298152 4088 298158 4140
rect 304258 3952 304264 4004
rect 304316 3992 304322 4004
rect 307938 3992 307944 4004
rect 304316 3964 307944 3992
rect 304316 3952 304322 3964
rect 307938 3952 307944 3964
rect 307996 3952 308002 4004
rect 11146 3544 11152 3596
rect 11204 3584 11210 3596
rect 12250 3584 12256 3596
rect 11204 3556 12256 3584
rect 11204 3544 11210 3556
rect 12250 3544 12256 3556
rect 12308 3544 12314 3596
rect 35986 3544 35992 3596
rect 36044 3584 36050 3596
rect 37090 3584 37096 3596
rect 36044 3556 37096 3584
rect 36044 3544 36050 3556
rect 37090 3544 37096 3556
rect 37148 3544 37154 3596
rect 44266 3544 44272 3596
rect 44324 3584 44330 3596
rect 45370 3584 45376 3596
rect 44324 3556 45376 3584
rect 44324 3544 44330 3556
rect 45370 3544 45376 3556
rect 45428 3544 45434 3596
rect 64322 3544 64328 3596
rect 64380 3584 64386 3596
rect 64782 3584 64788 3596
rect 64380 3556 64788 3584
rect 64380 3544 64386 3556
rect 64782 3544 64788 3556
rect 64840 3544 64846 3596
rect 69106 3544 69112 3596
rect 69164 3584 69170 3596
rect 70210 3584 70216 3596
rect 69164 3556 70216 3584
rect 69164 3544 69170 3556
rect 70210 3544 70216 3556
rect 70268 3544 70274 3596
rect 119890 3544 119896 3596
rect 119948 3584 119954 3596
rect 126238 3584 126244 3596
rect 119948 3556 126244 3584
rect 119948 3544 119954 3556
rect 126238 3544 126244 3556
rect 126296 3544 126302 3596
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3970 3516 3976 3528
rect 2924 3488 3976 3516
rect 2924 3476 2930 3488
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 8754 3476 8760 3528
rect 8812 3516 8818 3528
rect 9582 3516 9588 3528
rect 8812 3488 9588 3516
rect 8812 3476 8818 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 9950 3476 9956 3528
rect 10008 3516 10014 3528
rect 10962 3516 10968 3528
rect 10008 3488 10968 3516
rect 10008 3476 10014 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 17034 3476 17040 3528
rect 17092 3516 17098 3528
rect 17862 3516 17868 3528
rect 17092 3488 17868 3516
rect 17092 3476 17098 3488
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 18230 3476 18236 3528
rect 18288 3516 18294 3528
rect 19242 3516 19248 3528
rect 18288 3488 19248 3516
rect 18288 3476 18294 3488
rect 19242 3476 19248 3488
rect 19300 3476 19306 3528
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 20530 3516 20536 3528
rect 19484 3488 20536 3516
rect 19484 3476 19490 3488
rect 20530 3476 20536 3488
rect 20588 3476 20594 3528
rect 24210 3476 24216 3528
rect 24268 3516 24274 3528
rect 24762 3516 24768 3528
rect 24268 3488 24768 3516
rect 24268 3476 24274 3488
rect 24762 3476 24768 3488
rect 24820 3476 24826 3528
rect 25314 3476 25320 3528
rect 25372 3516 25378 3528
rect 26142 3516 26148 3528
rect 25372 3488 26148 3516
rect 25372 3476 25378 3488
rect 26142 3476 26148 3488
rect 26200 3476 26206 3528
rect 27706 3476 27712 3528
rect 27764 3516 27770 3528
rect 28810 3516 28816 3528
rect 27764 3488 28816 3516
rect 27764 3476 27770 3488
rect 28810 3476 28816 3488
rect 28868 3476 28874 3528
rect 32398 3476 32404 3528
rect 32456 3516 32462 3528
rect 33042 3516 33048 3528
rect 32456 3488 33048 3516
rect 32456 3476 32462 3488
rect 33042 3476 33048 3488
rect 33100 3476 33106 3528
rect 33594 3476 33600 3528
rect 33652 3516 33658 3528
rect 34422 3516 34428 3528
rect 33652 3488 34428 3516
rect 33652 3476 33658 3488
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
rect 34790 3476 34796 3528
rect 34848 3516 34854 3528
rect 35802 3516 35808 3528
rect 34848 3488 35808 3516
rect 34848 3476 34854 3488
rect 35802 3476 35808 3488
rect 35860 3476 35866 3528
rect 40678 3476 40684 3528
rect 40736 3516 40742 3528
rect 41230 3516 41236 3528
rect 40736 3488 41236 3516
rect 40736 3476 40742 3488
rect 41230 3476 41236 3488
rect 41288 3476 41294 3528
rect 43070 3476 43076 3528
rect 43128 3516 43134 3528
rect 43990 3516 43996 3528
rect 43128 3488 43996 3516
rect 43128 3476 43134 3488
rect 43990 3476 43996 3488
rect 44048 3476 44054 3528
rect 48958 3476 48964 3528
rect 49016 3516 49022 3528
rect 49602 3516 49608 3528
rect 49016 3488 49608 3516
rect 49016 3476 49022 3488
rect 49602 3476 49608 3488
rect 49660 3476 49666 3528
rect 50154 3476 50160 3528
rect 50212 3516 50218 3528
rect 50890 3516 50896 3528
rect 50212 3488 50896 3516
rect 50212 3476 50218 3488
rect 50890 3476 50896 3488
rect 50948 3476 50954 3528
rect 52546 3476 52552 3528
rect 52604 3516 52610 3528
rect 53558 3516 53564 3528
rect 52604 3488 53564 3516
rect 52604 3476 52610 3488
rect 53558 3476 53564 3488
rect 53616 3476 53622 3528
rect 56042 3476 56048 3528
rect 56100 3516 56106 3528
rect 56502 3516 56508 3528
rect 56100 3488 56508 3516
rect 56100 3476 56106 3488
rect 56502 3476 56508 3488
rect 56560 3476 56566 3528
rect 57238 3476 57244 3528
rect 57296 3516 57302 3528
rect 57882 3516 57888 3528
rect 57296 3488 57888 3516
rect 57296 3476 57302 3488
rect 57882 3476 57888 3488
rect 57940 3476 57946 3528
rect 58434 3476 58440 3528
rect 58492 3516 58498 3528
rect 59170 3516 59176 3528
rect 58492 3488 59176 3516
rect 58492 3476 58498 3488
rect 59170 3476 59176 3488
rect 59228 3476 59234 3528
rect 59630 3476 59636 3528
rect 59688 3516 59694 3528
rect 60642 3516 60648 3528
rect 59688 3488 60648 3516
rect 59688 3476 59694 3488
rect 60642 3476 60648 3488
rect 60700 3476 60706 3528
rect 63218 3476 63224 3528
rect 63276 3516 63282 3528
rect 97810 3516 97816 3528
rect 63276 3488 97816 3516
rect 63276 3476 63282 3488
rect 97810 3476 97816 3488
rect 97868 3476 97874 3528
rect 98638 3476 98644 3528
rect 98696 3516 98702 3528
rect 99282 3516 99288 3528
rect 98696 3488 99288 3516
rect 98696 3476 98702 3488
rect 99282 3476 99288 3488
rect 99340 3476 99346 3528
rect 99834 3476 99840 3528
rect 99892 3516 99898 3528
rect 100662 3516 100668 3528
rect 99892 3488 100668 3516
rect 99892 3476 99898 3488
rect 100662 3476 100668 3488
rect 100720 3476 100726 3528
rect 101030 3476 101036 3528
rect 101088 3516 101094 3528
rect 102042 3516 102048 3528
rect 101088 3488 102048 3516
rect 101088 3476 101094 3488
rect 102042 3476 102048 3488
rect 102100 3476 102106 3528
rect 105722 3476 105728 3528
rect 105780 3516 105786 3528
rect 106182 3516 106188 3528
rect 105780 3488 106188 3516
rect 105780 3476 105786 3488
rect 106182 3476 106188 3488
rect 106240 3476 106246 3528
rect 106918 3476 106924 3528
rect 106976 3516 106982 3528
rect 107562 3516 107568 3528
rect 106976 3488 107568 3516
rect 106976 3476 106982 3488
rect 107562 3476 107568 3488
rect 107620 3476 107626 3528
rect 108114 3476 108120 3528
rect 108172 3516 108178 3528
rect 108942 3516 108948 3528
rect 108172 3488 108948 3516
rect 108172 3476 108178 3488
rect 108942 3476 108948 3488
rect 109000 3476 109006 3528
rect 109310 3476 109316 3528
rect 109368 3516 109374 3528
rect 110322 3516 110328 3528
rect 109368 3488 110328 3516
rect 109368 3476 109374 3488
rect 110322 3476 110328 3488
rect 110380 3476 110386 3528
rect 110506 3476 110512 3528
rect 110564 3516 110570 3528
rect 111518 3516 111524 3528
rect 110564 3488 111524 3516
rect 110564 3476 110570 3488
rect 111518 3476 111524 3488
rect 111576 3476 111582 3528
rect 114002 3476 114008 3528
rect 114060 3516 114066 3528
rect 114462 3516 114468 3528
rect 114060 3488 114468 3516
rect 114060 3476 114066 3488
rect 114462 3476 114468 3488
rect 114520 3476 114526 3528
rect 115198 3476 115204 3528
rect 115256 3516 115262 3528
rect 115842 3516 115848 3528
rect 115256 3488 115848 3516
rect 115256 3476 115262 3488
rect 115842 3476 115848 3488
rect 115900 3476 115906 3528
rect 116394 3476 116400 3528
rect 116452 3516 116458 3528
rect 117038 3516 117044 3528
rect 116452 3488 117044 3516
rect 116452 3476 116458 3488
rect 117038 3476 117044 3488
rect 117096 3476 117102 3528
rect 117590 3476 117596 3528
rect 117648 3516 117654 3528
rect 118602 3516 118608 3528
rect 117648 3488 118608 3516
rect 117648 3476 117654 3488
rect 118602 3476 118608 3488
rect 118660 3476 118666 3528
rect 118786 3476 118792 3528
rect 118844 3516 118850 3528
rect 119982 3516 119988 3528
rect 118844 3488 119988 3516
rect 118844 3476 118850 3488
rect 119982 3476 119988 3488
rect 120040 3476 120046 3528
rect 123478 3476 123484 3528
rect 123536 3516 123542 3528
rect 124122 3516 124128 3528
rect 123536 3488 124128 3516
rect 123536 3476 123542 3488
rect 124122 3476 124128 3488
rect 124180 3476 124186 3528
rect 129366 3476 129372 3528
rect 129424 3516 129430 3528
rect 130378 3516 130384 3528
rect 129424 3488 130384 3516
rect 129424 3476 129430 3488
rect 130378 3476 130384 3488
rect 130436 3476 130442 3528
rect 202138 3476 202144 3528
rect 202196 3516 202202 3528
rect 257062 3516 257068 3528
rect 202196 3488 257068 3516
rect 202196 3476 202202 3488
rect 257062 3476 257068 3488
rect 257120 3476 257126 3528
rect 313918 3476 313924 3528
rect 313976 3516 313982 3528
rect 315022 3516 315028 3528
rect 313976 3488 315028 3516
rect 313976 3476 313982 3488
rect 315022 3476 315028 3488
rect 315080 3476 315086 3528
rect 316034 3476 316040 3528
rect 316092 3516 316098 3528
rect 317322 3516 317328 3528
rect 316092 3488 317328 3516
rect 316092 3476 316098 3488
rect 317322 3476 317328 3488
rect 317380 3476 317386 3528
rect 324314 3476 324320 3528
rect 324372 3516 324378 3528
rect 325602 3516 325608 3528
rect 324372 3488 325608 3516
rect 324372 3476 324378 3488
rect 325602 3476 325608 3488
rect 325660 3476 325666 3528
rect 335998 3476 336004 3528
rect 336056 3516 336062 3528
rect 337470 3516 337476 3528
rect 336056 3488 337476 3516
rect 336056 3476 336062 3488
rect 337470 3476 337476 3488
rect 337528 3476 337534 3528
rect 340874 3476 340880 3528
rect 340932 3516 340938 3528
rect 342162 3516 342168 3528
rect 340932 3488 342168 3516
rect 340932 3476 340938 3488
rect 342162 3476 342168 3488
rect 342220 3476 342226 3528
rect 350442 3476 350448 3528
rect 350500 3516 350506 3528
rect 353294 3516 353300 3528
rect 350500 3488 353300 3516
rect 350500 3476 350506 3488
rect 353294 3476 353300 3488
rect 353352 3476 353358 3528
rect 582190 3476 582196 3528
rect 582248 3516 582254 3528
rect 583478 3516 583484 3528
rect 582248 3488 583484 3516
rect 582248 3476 582254 3488
rect 583478 3476 583484 3488
rect 583536 3476 583542 3528
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 15838 3448 15844 3460
rect 6512 3420 15844 3448
rect 6512 3408 6518 3420
rect 15838 3408 15844 3420
rect 15896 3408 15902 3460
rect 26510 3408 26516 3460
rect 26568 3448 26574 3460
rect 26568 3420 64874 3448
rect 26568 3408 26574 3420
rect 64846 3380 64874 3420
rect 65518 3408 65524 3460
rect 65576 3448 65582 3460
rect 66162 3448 66168 3460
rect 65576 3420 66168 3448
rect 65576 3408 65582 3420
rect 66162 3408 66168 3420
rect 66220 3408 66226 3460
rect 67910 3408 67916 3460
rect 67968 3448 67974 3460
rect 68922 3448 68928 3460
rect 67968 3420 68928 3448
rect 67968 3408 67974 3420
rect 68922 3408 68928 3420
rect 68980 3408 68986 3460
rect 72602 3408 72608 3460
rect 72660 3448 72666 3460
rect 73062 3448 73068 3460
rect 72660 3420 73068 3448
rect 72660 3408 72666 3420
rect 73062 3408 73068 3420
rect 73120 3408 73126 3460
rect 74994 3408 75000 3460
rect 75052 3448 75058 3460
rect 75822 3448 75828 3460
rect 75052 3420 75828 3448
rect 75052 3408 75058 3420
rect 75822 3408 75828 3420
rect 75880 3408 75886 3460
rect 76190 3408 76196 3460
rect 76248 3448 76254 3460
rect 77202 3448 77208 3460
rect 76248 3420 77208 3448
rect 76248 3408 76254 3420
rect 77202 3408 77208 3420
rect 77260 3408 77266 3460
rect 80882 3408 80888 3460
rect 80940 3448 80946 3460
rect 81342 3448 81348 3460
rect 80940 3420 81348 3448
rect 80940 3408 80946 3420
rect 81342 3408 81348 3420
rect 81400 3408 81406 3460
rect 83274 3408 83280 3460
rect 83332 3448 83338 3460
rect 84102 3448 84108 3460
rect 83332 3420 84108 3448
rect 83332 3408 83338 3420
rect 84102 3408 84108 3420
rect 84160 3408 84166 3460
rect 84470 3408 84476 3460
rect 84528 3448 84534 3460
rect 85482 3448 85488 3460
rect 84528 3420 85488 3448
rect 84528 3408 84534 3420
rect 85482 3408 85488 3420
rect 85540 3408 85546 3460
rect 89162 3408 89168 3460
rect 89220 3448 89226 3460
rect 89622 3448 89628 3460
rect 89220 3420 89628 3448
rect 89220 3408 89226 3420
rect 89622 3408 89628 3420
rect 89680 3408 89686 3460
rect 91554 3408 91560 3460
rect 91612 3448 91618 3460
rect 92382 3448 92388 3460
rect 91612 3420 92388 3448
rect 91612 3408 91618 3420
rect 92382 3408 92388 3420
rect 92440 3408 92446 3460
rect 92750 3408 92756 3460
rect 92808 3448 92814 3460
rect 93762 3448 93768 3460
rect 92808 3420 93768 3448
rect 92808 3408 92814 3420
rect 93762 3408 93768 3420
rect 93820 3408 93826 3460
rect 97442 3408 97448 3460
rect 97500 3448 97506 3460
rect 97902 3448 97908 3460
rect 97500 3420 97908 3448
rect 97500 3408 97506 3420
rect 97902 3408 97908 3420
rect 97960 3408 97966 3460
rect 102226 3408 102232 3460
rect 102284 3448 102290 3460
rect 123386 3448 123392 3460
rect 102284 3420 123392 3448
rect 102284 3408 102290 3420
rect 123386 3408 123392 3420
rect 123444 3408 123450 3460
rect 124674 3408 124680 3460
rect 124732 3448 124738 3460
rect 214558 3448 214564 3460
rect 124732 3420 214564 3448
rect 124732 3408 124738 3420
rect 214558 3408 214564 3420
rect 214616 3408 214622 3460
rect 285398 3408 285404 3460
rect 285456 3448 285462 3460
rect 306466 3448 306472 3460
rect 285456 3420 306472 3448
rect 285456 3408 285462 3420
rect 306466 3408 306472 3420
rect 306524 3408 306530 3460
rect 323578 3408 323584 3460
rect 323636 3448 323642 3460
rect 332686 3448 332692 3460
rect 323636 3420 332692 3448
rect 323636 3408 323642 3420
rect 332686 3408 332692 3420
rect 332744 3408 332750 3460
rect 71038 3380 71044 3392
rect 64846 3352 71044 3380
rect 71038 3340 71044 3352
rect 71096 3340 71102 3392
rect 78582 3340 78588 3392
rect 78640 3380 78646 3392
rect 87598 3380 87604 3392
rect 78640 3352 87604 3380
rect 78640 3340 78646 3352
rect 87598 3340 87604 3352
rect 87656 3340 87662 3392
rect 122282 3272 122288 3324
rect 122340 3312 122346 3324
rect 122742 3312 122748 3324
rect 122340 3284 122748 3312
rect 122340 3272 122346 3284
rect 122742 3272 122748 3284
rect 122800 3272 122806 3324
rect 346946 3272 346952 3324
rect 347004 3312 347010 3324
rect 351914 3312 351920 3324
rect 347004 3284 351920 3312
rect 347004 3272 347010 3284
rect 351914 3272 351920 3284
rect 351972 3272 351978 3324
rect 280798 3136 280804 3188
rect 280856 3176 280862 3188
rect 283098 3176 283104 3188
rect 280856 3148 283104 3176
rect 280856 3136 280862 3148
rect 283098 3136 283104 3148
rect 283156 3136 283162 3188
rect 269758 3068 269764 3120
rect 269816 3108 269822 3120
rect 272426 3108 272432 3120
rect 269816 3080 272432 3108
rect 269816 3068 269822 3080
rect 272426 3068 272432 3080
rect 272484 3068 272490 3120
rect 347038 3068 347044 3120
rect 347096 3108 347102 3120
rect 349246 3108 349252 3120
rect 347096 3080 349252 3108
rect 347096 3068 347102 3080
rect 349246 3068 349252 3080
rect 349304 3068 349310 3120
rect 90358 3000 90364 3052
rect 90416 3040 90422 3052
rect 91002 3040 91008 3052
rect 90416 3012 91008 3040
rect 90416 3000 90422 3012
rect 91002 3000 91008 3012
rect 91060 3000 91066 3052
rect 580994 3000 581000 3052
rect 581052 3040 581058 3052
rect 583386 3040 583392 3052
rect 581052 3012 583392 3040
rect 581052 3000 581058 3012
rect 583386 3000 583392 3012
rect 583444 3000 583450 3052
rect 93946 2932 93952 2984
rect 94004 2972 94010 2984
rect 94958 2972 94964 2984
rect 94004 2944 94964 2972
rect 94004 2932 94010 2944
rect 94958 2932 94964 2944
rect 95016 2932 95022 2984
rect 51350 2116 51356 2168
rect 51408 2156 51414 2168
rect 90266 2156 90272 2168
rect 51408 2128 90272 2156
rect 51408 2116 51414 2128
rect 90266 2116 90272 2128
rect 90324 2116 90330 2168
rect 198090 2116 198096 2168
rect 198148 2156 198154 2168
rect 254670 2156 254676 2168
rect 198148 2128 254676 2156
rect 198148 2116 198154 2128
rect 254670 2116 254676 2128
rect 254728 2116 254734 2168
rect 7650 2048 7656 2100
rect 7708 2088 7714 2100
rect 32306 2088 32312 2100
rect 7708 2060 32312 2088
rect 7708 2048 7714 2060
rect 32306 2048 32312 2060
rect 32364 2048 32370 2100
rect 87966 2048 87972 2100
rect 88024 2088 88030 2100
rect 222838 2088 222844 2100
rect 88024 2060 222844 2088
rect 88024 2048 88030 2060
rect 222838 2048 222844 2060
rect 222896 2048 222902 2100
<< via1 >>
rect 122104 703604 122156 703656
rect 234988 703604 235040 703656
rect 75828 703536 75880 703588
rect 202604 703536 202656 703588
rect 67640 703468 67692 703520
rect 267464 703468 267516 703520
rect 93768 703400 93820 703452
rect 300124 703400 300176 703452
rect 59268 703332 59320 703384
rect 283840 703332 283892 703384
rect 73068 703264 73120 703316
rect 332508 703264 332560 703316
rect 130384 703196 130436 703248
rect 413652 703196 413704 703248
rect 61844 703128 61896 703180
rect 348792 703128 348844 703180
rect 101496 703060 101548 703112
rect 397460 703060 397512 703112
rect 124864 702992 124916 703044
rect 429844 702992 429896 703044
rect 57888 702924 57940 702976
rect 364984 702924 365036 702976
rect 126244 702856 126296 702908
rect 462320 702856 462372 702908
rect 71044 702788 71096 702840
rect 494796 702788 494848 702840
rect 97908 702720 97960 702772
rect 478512 702720 478564 702772
rect 129004 702652 129056 702704
rect 543464 702652 543516 702704
rect 8116 702584 8168 702636
rect 89812 702584 89864 702636
rect 94504 702584 94556 702636
rect 527180 702584 527232 702636
rect 53748 702516 53800 702568
rect 580264 702516 580316 702568
rect 66168 702448 66220 702500
rect 559656 702448 559708 702500
rect 83464 700340 83516 700392
rect 89168 700340 89220 700392
rect 40500 700272 40552 700324
rect 89076 700272 89128 700324
rect 133144 700272 133196 700324
rect 218980 700272 219032 700324
rect 24308 699660 24360 699712
rect 25504 699660 25556 699712
rect 3424 683136 3476 683188
rect 11704 683136 11756 683188
rect 3516 670692 3568 670744
rect 14464 670692 14516 670744
rect 3424 658112 3476 658164
rect 7564 658112 7616 658164
rect 3424 632068 3476 632120
rect 17224 632068 17276 632120
rect 2780 619080 2832 619132
rect 4804 619080 4856 619132
rect 3240 605820 3292 605872
rect 87604 605820 87656 605872
rect 67456 599564 67508 599616
rect 104900 599564 104952 599616
rect 79968 597524 80020 597576
rect 106924 597524 106976 597576
rect 67548 596776 67600 596828
rect 169760 596776 169812 596828
rect 25504 596096 25556 596148
rect 79968 596096 80020 596148
rect 108304 595416 108356 595468
rect 582748 595416 582800 595468
rect 77024 594804 77076 594856
rect 101404 594804 101456 594856
rect 87604 594532 87656 594584
rect 91192 594532 91244 594584
rect 83464 593376 83516 593428
rect 110420 593376 110472 593428
rect 7564 592628 7616 592680
rect 69020 592628 69072 592680
rect 75736 592084 75788 592136
rect 96620 592084 96672 592136
rect 79784 592016 79836 592068
rect 105544 592016 105596 592068
rect 78404 590792 78456 590844
rect 103520 590792 103572 590844
rect 61936 590656 61988 590708
rect 70860 590656 70912 590708
rect 71688 590656 71740 590708
rect 75000 590656 75052 590708
rect 75736 590656 75788 590708
rect 3424 589908 3476 589960
rect 71688 589908 71740 589960
rect 81348 589432 81400 589484
rect 70308 589364 70360 589416
rect 89720 589364 89772 589416
rect 108304 589296 108356 589348
rect 69480 588616 69532 588668
rect 88984 588616 89036 588668
rect 85580 588548 85632 588600
rect 114468 588548 114520 588600
rect 84384 588412 84436 588464
rect 86224 588412 86276 588464
rect 89168 588412 89220 588464
rect 63316 587868 63368 587920
rect 66812 587868 66864 587920
rect 92480 587800 92532 587852
rect 114468 587800 114520 587852
rect 122104 587800 122156 587852
rect 59176 586508 59228 586560
rect 66260 586508 66312 586560
rect 89168 585760 89220 585812
rect 116584 585760 116636 585812
rect 50896 585148 50948 585200
rect 67732 585148 67784 585200
rect 91928 584400 91980 584452
rect 93768 584400 93820 584452
rect 115204 584400 115256 584452
rect 91928 583652 91980 583704
rect 93768 583652 93820 583704
rect 94504 583652 94556 583704
rect 48136 582360 48188 582412
rect 66812 582360 66864 582412
rect 64696 581000 64748 581052
rect 66996 581000 67048 581052
rect 91100 581000 91152 581052
rect 102784 581000 102836 581052
rect 91100 578212 91152 578264
rect 121552 578212 121604 578264
rect 100668 577464 100720 577516
rect 582472 577464 582524 577516
rect 91100 576852 91152 576904
rect 100668 576852 100720 576904
rect 17224 576104 17276 576156
rect 34520 576104 34572 576156
rect 91192 576104 91244 576156
rect 105636 576104 105688 576156
rect 34520 575492 34572 575544
rect 35808 575492 35860 575544
rect 66904 575492 66956 575544
rect 89076 575492 89128 575544
rect 91284 575492 91336 575544
rect 55036 574744 55088 574796
rect 67456 574744 67508 574796
rect 91928 574744 91980 574796
rect 93768 574744 93820 574796
rect 101496 574744 101548 574796
rect 41328 572704 41380 572756
rect 66444 572704 66496 572756
rect 91100 572704 91152 572756
rect 120724 572704 120776 572756
rect 91100 571412 91152 571464
rect 94504 571412 94556 571464
rect 49608 571344 49660 571396
rect 66444 571344 66496 571396
rect 91192 571344 91244 571396
rect 126980 571344 127032 571396
rect 91100 569916 91152 569968
rect 128360 569916 128412 569968
rect 93768 569168 93820 569220
rect 123484 569168 123536 569220
rect 64788 568556 64840 568608
rect 66812 568556 66864 568608
rect 91284 567808 91336 567860
rect 124220 567808 124272 567860
rect 57704 567196 57756 567248
rect 66904 567196 66956 567248
rect 53656 566448 53708 566500
rect 67548 566448 67600 566500
rect 91100 565836 91152 565888
rect 101496 565836 101548 565888
rect 60648 564408 60700 564460
rect 66628 564408 66680 564460
rect 91100 564408 91152 564460
rect 120632 564408 120684 564460
rect 50988 564340 51040 564392
rect 53748 564340 53800 564392
rect 66444 564340 66496 564392
rect 91100 563048 91152 563100
rect 129740 563048 129792 563100
rect 37188 561688 37240 561740
rect 66444 561688 66496 561740
rect 44088 560260 44140 560312
rect 66628 560260 66680 560312
rect 56508 558900 56560 558952
rect 66628 558900 66680 558952
rect 48228 557540 48280 557592
rect 67640 557540 67692 557592
rect 91192 557540 91244 557592
rect 125600 557540 125652 557592
rect 91192 556180 91244 556232
rect 122104 556180 122156 556232
rect 58992 554752 59044 554804
rect 66352 554752 66404 554804
rect 91192 554752 91244 554804
rect 108948 554752 109000 554804
rect 582472 554752 582524 554804
rect 59268 554684 59320 554736
rect 65524 554684 65576 554736
rect 66260 554684 66312 554736
rect 3332 553392 3384 553444
rect 32404 553392 32456 553444
rect 107108 553052 107160 553104
rect 109040 553052 109092 553104
rect 91192 552100 91244 552152
rect 107016 552100 107068 552152
rect 91284 552032 91336 552084
rect 134524 552032 134576 552084
rect 63408 549244 63460 549296
rect 66536 549244 66588 549296
rect 91192 549244 91244 549296
rect 104256 549244 104308 549296
rect 91836 548496 91888 548548
rect 121460 548496 121512 548548
rect 62028 547884 62080 547936
rect 66536 547884 66588 547936
rect 61844 547748 61896 547800
rect 66812 547748 66864 547800
rect 53748 547136 53800 547188
rect 61844 547136 61896 547188
rect 91284 546456 91336 546508
rect 104164 546456 104216 546508
rect 57796 545708 57848 545760
rect 66168 545708 66220 545760
rect 91284 545708 91336 545760
rect 96436 545708 96488 545760
rect 126244 545708 126296 545760
rect 52368 545028 52420 545080
rect 57888 545028 57940 545080
rect 66812 545028 66864 545080
rect 91284 544348 91336 544400
rect 96528 544348 96580 544400
rect 129004 544348 129056 544400
rect 11704 542988 11756 543040
rect 39948 542988 40000 543040
rect 95884 542988 95936 543040
rect 117320 542988 117372 543040
rect 39948 542376 40000 542428
rect 66812 542376 66864 542428
rect 91284 542376 91336 542428
rect 97264 542376 97316 542428
rect 14464 541628 14516 541680
rect 67088 541628 67140 541680
rect 91284 541628 91336 541680
rect 136640 541628 136692 541680
rect 67548 540880 67600 540932
rect 68652 540880 68704 540932
rect 582656 540880 582708 540932
rect 3424 540200 3476 540252
rect 91284 539656 91336 539708
rect 93124 539656 93176 539708
rect 55128 539588 55180 539640
rect 67548 539588 67600 539640
rect 69848 539588 69900 539640
rect 67088 539452 67140 539504
rect 67548 539452 67600 539504
rect 67824 538908 67876 538960
rect 74724 538908 74776 538960
rect 3424 538840 3476 538892
rect 89904 538840 89956 538892
rect 80336 538228 80388 538280
rect 80796 538228 80848 538280
rect 582564 538228 582616 538280
rect 32404 538160 32456 538212
rect 70676 538160 70728 538212
rect 86868 538160 86920 538212
rect 133144 538160 133196 538212
rect 72424 537480 72476 537532
rect 579804 537480 579856 537532
rect 76012 536732 76064 536784
rect 124864 536732 124916 536784
rect 85488 536188 85540 536240
rect 86224 536188 86276 536240
rect 66168 536120 66220 536172
rect 76012 536120 76064 536172
rect 4804 536052 4856 536104
rect 45468 536052 45520 536104
rect 73160 536052 73212 536104
rect 73160 535440 73212 535492
rect 73988 535440 74040 535492
rect 7564 534692 7616 534744
rect 91376 534692 91428 534744
rect 56416 534012 56468 534064
rect 580264 534012 580316 534064
rect 78680 533400 78732 533452
rect 79508 533400 79560 533452
rect 5448 533332 5500 533384
rect 91192 533332 91244 533384
rect 66076 531972 66128 532024
rect 77944 531972 77996 532024
rect 15844 530544 15896 530596
rect 91100 530544 91152 530596
rect 3516 514768 3568 514820
rect 14464 514768 14516 514820
rect 102784 512592 102836 512644
rect 122932 512592 122984 512644
rect 44088 511232 44140 511284
rect 580172 511232 580224 511284
rect 3332 502052 3384 502104
rect 7564 502052 7616 502104
rect 4068 475328 4120 475380
rect 5448 475328 5500 475380
rect 11704 475328 11756 475380
rect 54852 468460 54904 468512
rect 77300 468460 77352 468512
rect 52276 465672 52328 465724
rect 95884 465672 95936 465724
rect 59084 464312 59136 464364
rect 80060 464312 80112 464364
rect 50804 462952 50856 463004
rect 75920 462952 75972 463004
rect 94504 462952 94556 463004
rect 125692 462952 125744 463004
rect 2780 462544 2832 462596
rect 4804 462544 4856 462596
rect 52276 461592 52328 461644
rect 78680 461592 78732 461644
rect 63316 460912 63368 460964
rect 86960 460912 87012 460964
rect 64696 460164 64748 460216
rect 78680 460164 78732 460216
rect 64696 458872 64748 458924
rect 70492 458872 70544 458924
rect 59176 458804 59228 458856
rect 85580 458804 85632 458856
rect 77300 458192 77352 458244
rect 77944 458192 77996 458244
rect 124864 458192 124916 458244
rect 61752 457512 61804 457564
rect 73160 457512 73212 457564
rect 50896 457444 50948 457496
rect 83464 457444 83516 457496
rect 105636 457444 105688 457496
rect 123024 457444 123076 457496
rect 98552 456764 98604 456816
rect 98736 456764 98788 456816
rect 151084 456764 151136 456816
rect 61936 456016 61988 456068
rect 91100 456016 91152 456068
rect 101496 456016 101548 456068
rect 123208 456016 123260 456068
rect 112444 455404 112496 455456
rect 152464 455404 152516 455456
rect 55036 454724 55088 454776
rect 72056 454724 72108 454776
rect 35808 454656 35860 454708
rect 71044 454656 71096 454708
rect 91100 454044 91152 454096
rect 158720 454044 158772 454096
rect 67732 453976 67784 454028
rect 68284 453976 68336 454028
rect 49608 453296 49660 453348
rect 68744 453296 68796 453348
rect 91744 453296 91796 453348
rect 121644 453296 121696 453348
rect 68284 452684 68336 452736
rect 82084 452684 82136 452736
rect 72056 452616 72108 452668
rect 127624 452616 127676 452668
rect 61844 451936 61896 451988
rect 72424 451936 72476 451988
rect 3424 451868 3476 451920
rect 120816 451868 120868 451920
rect 14464 451188 14516 451240
rect 112444 451188 112496 451240
rect 116584 449964 116636 450016
rect 161572 449964 161624 450016
rect 71044 449896 71096 449948
rect 73252 449896 73304 449948
rect 144184 449896 144236 449948
rect 64604 449216 64656 449268
rect 74632 449216 74684 449268
rect 48136 449148 48188 449200
rect 80060 449148 80112 449200
rect 169024 449148 169076 449200
rect 169668 449148 169720 449200
rect 582472 449148 582524 449200
rect 3148 448536 3200 448588
rect 14464 448536 14516 448588
rect 80060 448536 80112 448588
rect 80888 448536 80940 448588
rect 169024 448536 169076 448588
rect 4804 447788 4856 447840
rect 68468 447788 68520 447840
rect 115204 447788 115256 447840
rect 124312 447788 124364 447840
rect 68468 447176 68520 447228
rect 68652 447176 68704 447228
rect 103520 447176 103572 447228
rect 49608 447108 49660 447160
rect 74724 447108 74776 447160
rect 95884 447108 95936 447160
rect 171140 447108 171192 447160
rect 78680 446904 78732 446956
rect 79140 446904 79192 446956
rect 41328 445816 41380 445868
rect 79140 445816 79192 445868
rect 106924 445816 106976 445868
rect 124956 445816 125008 445868
rect 76564 445748 76616 445800
rect 155224 445748 155276 445800
rect 54944 444456 54996 444508
rect 92480 444456 92532 444508
rect 93078 444456 93130 444508
rect 101404 444456 101456 444508
rect 126244 444456 126296 444508
rect 4804 444388 4856 444440
rect 118700 444388 118752 444440
rect 124128 444320 124180 444372
rect 132500 444320 132552 444372
rect 133788 444320 133840 444372
rect 133788 443640 133840 443692
rect 165620 443640 165672 443692
rect 67272 442892 67324 442944
rect 67732 442892 67784 442944
rect 124128 441600 124180 441652
rect 133144 441600 133196 441652
rect 56508 440852 56560 440904
rect 68284 440852 68336 440904
rect 64788 439016 64840 439068
rect 66996 439016 67048 439068
rect 67272 439016 67324 439068
rect 124128 438880 124180 438932
rect 186964 438880 187016 438932
rect 124128 438132 124180 438184
rect 124312 438132 124364 438184
rect 157984 438132 158036 438184
rect 57704 437452 57756 437504
rect 60556 437452 60608 437504
rect 66812 437452 66864 437504
rect 53656 435344 53708 435396
rect 66812 435344 66864 435396
rect 124128 432556 124180 432608
rect 135168 432556 135220 432608
rect 582380 432556 582432 432608
rect 60648 432012 60700 432064
rect 66904 432012 66956 432064
rect 50988 431876 51040 431928
rect 66904 431876 66956 431928
rect 48136 430584 48188 430636
rect 50988 430584 51040 430636
rect 36728 429088 36780 429140
rect 37188 429088 37240 429140
rect 66812 429088 66864 429140
rect 22744 428408 22796 428460
rect 36728 428408 36780 428460
rect 44088 425688 44140 425740
rect 57888 425688 57940 425740
rect 57704 425076 57756 425128
rect 57888 425076 57940 425128
rect 66260 425076 66312 425128
rect 56416 424328 56468 424380
rect 66076 424328 66128 424380
rect 66260 424328 66312 424380
rect 3148 422900 3200 422952
rect 15844 422900 15896 422952
rect 123024 422288 123076 422340
rect 123484 422288 123536 422340
rect 172520 422288 172572 422340
rect 48228 421540 48280 421592
rect 61384 421540 61436 421592
rect 66260 421540 66312 421592
rect 121552 418072 121604 418124
rect 126980 418072 127032 418124
rect 58992 416780 59044 416832
rect 63316 416780 63368 416832
rect 66904 416780 66956 416832
rect 65524 415148 65576 415200
rect 66444 415148 66496 415200
rect 124128 415148 124180 415200
rect 125692 415148 125744 415200
rect 57888 414672 57940 414724
rect 65524 414672 65576 414724
rect 123116 413924 123168 413976
rect 128360 413924 128412 413976
rect 121644 409844 121696 409896
rect 129096 409844 129148 409896
rect 63408 408416 63460 408468
rect 65892 408416 65944 408468
rect 66536 408416 66588 408468
rect 124128 407736 124180 407788
rect 135904 407736 135956 407788
rect 122104 407056 122156 407108
rect 122932 407056 122984 407108
rect 57612 406512 57664 406564
rect 57796 406512 57848 406564
rect 123208 406104 123260 406156
rect 125048 406104 125100 406156
rect 62028 405764 62080 405816
rect 64788 405764 64840 405816
rect 66628 405764 66680 405816
rect 57980 403588 58032 403640
rect 66352 403588 66404 403640
rect 163504 403588 163556 403640
rect 582380 403588 582432 403640
rect 120632 402976 120684 403028
rect 163504 402976 163556 403028
rect 53656 402228 53708 402280
rect 57980 402228 58032 402280
rect 50896 401548 50948 401600
rect 57612 401548 57664 401600
rect 66812 401548 66864 401600
rect 124128 401480 124180 401532
rect 129740 401480 129792 401532
rect 129740 400188 129792 400240
rect 130384 400188 130436 400240
rect 60004 399440 60056 399492
rect 66352 399440 66404 399492
rect 123484 398828 123536 398880
rect 124956 398828 125008 398880
rect 2780 398692 2832 398744
rect 4804 398692 4856 398744
rect 43996 398080 44048 398132
rect 52368 398080 52420 398132
rect 60004 398080 60056 398132
rect 39948 396720 40000 396772
rect 66996 396720 67048 396772
rect 121460 396040 121512 396092
rect 180064 396040 180116 396092
rect 123668 395496 123720 395548
rect 125600 395496 125652 395548
rect 55128 393252 55180 393304
rect 66260 393252 66312 393304
rect 124956 391960 125008 392012
rect 172612 391960 172664 392012
rect 15844 391348 15896 391400
rect 124956 391348 125008 391400
rect 111708 389784 111760 389836
rect 121552 389784 121604 389836
rect 61752 389240 61804 389292
rect 77392 389240 77444 389292
rect 11704 389172 11756 389224
rect 111616 389172 111668 389224
rect 102600 389104 102652 389156
rect 105544 389104 105596 389156
rect 117872 389104 117924 389156
rect 134524 389104 134576 389156
rect 169760 389172 169812 389224
rect 64696 388424 64748 388476
rect 71780 388424 71832 388476
rect 93400 388424 93452 388476
rect 100024 388424 100076 388476
rect 101404 388424 101456 388476
rect 120172 388424 120224 388476
rect 93768 388356 93820 388408
rect 94228 388356 94280 388408
rect 71780 387812 71832 387864
rect 73160 387812 73212 387864
rect 111616 387812 111668 387864
rect 112444 387812 112496 387864
rect 45468 387744 45520 387796
rect 76564 387744 76616 387796
rect 3424 387064 3476 387116
rect 89720 387064 89772 387116
rect 104072 387064 104124 387116
rect 135076 387064 135128 387116
rect 136640 387064 136692 387116
rect 61844 386316 61896 386368
rect 74632 386316 74684 386368
rect 77208 385636 77260 385688
rect 113180 385636 113232 385688
rect 65984 384956 66036 385008
rect 85580 384956 85632 385008
rect 86224 384956 86276 385008
rect 15844 384276 15896 384328
rect 123116 384276 123168 384328
rect 110236 382916 110288 382968
rect 177488 382916 177540 382968
rect 7564 382236 7616 382288
rect 118700 382236 118752 382288
rect 119436 382236 119488 382288
rect 4804 381488 4856 381540
rect 105636 381488 105688 381540
rect 175280 381488 175332 381540
rect 50804 380808 50856 380860
rect 81440 380808 81492 380860
rect 81440 379584 81492 379636
rect 82084 379584 82136 379636
rect 72424 379516 72476 379568
rect 73068 379516 73120 379568
rect 188344 379516 188396 379568
rect 64788 378836 64840 378888
rect 108304 378836 108356 378888
rect 99288 378768 99340 378820
rect 165712 378768 165764 378820
rect 52276 378088 52328 378140
rect 86960 378088 87012 378140
rect 53564 376728 53616 376780
rect 53748 376728 53800 376780
rect 185584 376728 185636 376780
rect 67732 374620 67784 374672
rect 124956 374620 125008 374672
rect 86224 374008 86276 374060
rect 211804 374008 211856 374060
rect 60648 373260 60700 373312
rect 164884 373260 164936 373312
rect 122104 372580 122156 372632
rect 122748 372580 122800 372632
rect 204904 372580 204956 372632
rect 70308 371832 70360 371884
rect 167000 371832 167052 371884
rect 125048 371220 125100 371272
rect 125508 371220 125560 371272
rect 258080 371220 258132 371272
rect 139308 369928 139360 369980
rect 242164 369928 242216 369980
rect 125600 369860 125652 369912
rect 126244 369860 126296 369912
rect 231124 369860 231176 369912
rect 142804 369112 142856 369164
rect 174636 369112 174688 369164
rect 121368 368500 121420 368552
rect 182824 368500 182876 368552
rect 119436 367752 119488 367804
rect 171232 367752 171284 367804
rect 137928 367072 137980 367124
rect 327080 367072 327132 367124
rect 81348 366324 81400 366376
rect 96436 366324 96488 366376
rect 124864 365780 124916 365832
rect 214564 365780 214616 365832
rect 104900 365712 104952 365764
rect 224224 365712 224276 365764
rect 81440 365644 81492 365696
rect 82084 365644 82136 365696
rect 143448 364420 143500 364472
rect 238024 364420 238076 364472
rect 81440 364352 81492 364404
rect 238116 364352 238168 364404
rect 131120 362992 131172 363044
rect 214656 362992 214708 363044
rect 90364 362924 90416 362976
rect 188436 362924 188488 362976
rect 137284 362652 137336 362704
rect 137836 362652 137888 362704
rect 63224 362176 63276 362228
rect 87052 362176 87104 362228
rect 87972 362176 88024 362228
rect 137836 361632 137888 361684
rect 164240 361632 164292 361684
rect 87972 361564 88024 361616
rect 240232 361564 240284 361616
rect 50804 361496 50856 361548
rect 54852 361496 54904 361548
rect 82820 361496 82872 361548
rect 92296 360816 92348 360868
rect 118700 360816 118752 360868
rect 124956 360272 125008 360324
rect 178684 360272 178736 360324
rect 99288 360204 99340 360256
rect 226984 360204 227036 360256
rect 66076 359456 66128 359508
rect 127716 359456 127768 359508
rect 128360 358844 128412 358896
rect 181536 358844 181588 358896
rect 136640 358776 136692 358828
rect 238760 358776 238812 358828
rect 3516 358572 3568 358624
rect 7564 358572 7616 358624
rect 93768 358028 93820 358080
rect 131120 358028 131172 358080
rect 118700 357416 118752 357468
rect 225604 357416 225656 357468
rect 64788 356668 64840 356720
rect 111800 356668 111852 356720
rect 70400 356600 70452 356652
rect 71688 356600 71740 356652
rect 141424 356124 141476 356176
rect 231216 356124 231268 356176
rect 71688 356056 71740 356108
rect 255412 356056 255464 356108
rect 155224 355988 155276 356040
rect 155960 355988 156012 356040
rect 97816 355308 97868 355360
rect 155316 355308 155368 355360
rect 120080 354696 120132 354748
rect 203524 354696 203576 354748
rect 122656 353948 122708 354000
rect 127624 353948 127676 354000
rect 60556 353336 60608 353388
rect 162124 353336 162176 353388
rect 132408 353268 132460 353320
rect 320180 353268 320232 353320
rect 54852 352520 54904 352572
rect 86960 352520 87012 352572
rect 104808 352520 104860 352572
rect 120724 352520 120776 352572
rect 89076 351976 89128 352028
rect 92664 351976 92716 352028
rect 85488 351908 85540 351960
rect 90364 351908 90416 351960
rect 125508 351976 125560 352028
rect 125692 351976 125744 352028
rect 144184 351976 144236 352028
rect 146300 351976 146352 352028
rect 195244 351976 195296 352028
rect 251272 351908 251324 351960
rect 88984 351840 89036 351892
rect 129648 351840 129700 351892
rect 118792 350548 118844 350600
rect 119344 350548 119396 350600
rect 249892 350548 249944 350600
rect 79968 349800 80020 349852
rect 111340 349800 111392 349852
rect 112444 349800 112496 349852
rect 156052 349800 156104 349852
rect 133880 349120 133932 349172
rect 236644 349120 236696 349172
rect 83464 348372 83516 348424
rect 109684 348372 109736 348424
rect 121644 347828 121696 347880
rect 122748 347828 122800 347880
rect 196624 347828 196676 347880
rect 77208 347760 77260 347812
rect 204352 347760 204404 347812
rect 79324 347692 79376 347744
rect 121644 347692 121696 347744
rect 204168 347692 204220 347744
rect 582380 347692 582432 347744
rect 152464 347080 152516 347132
rect 161664 347080 161716 347132
rect 85580 346944 85632 346996
rect 86316 346944 86368 346996
rect 203064 347012 203116 347064
rect 204168 347012 204220 347064
rect 2780 346264 2832 346316
rect 4804 346264 4856 346316
rect 115204 345108 115256 345160
rect 229192 345108 229244 345160
rect 91008 345040 91060 345092
rect 210424 345040 210476 345092
rect 87972 343680 88024 343732
rect 216036 343680 216088 343732
rect 73804 343612 73856 343664
rect 209136 343612 209188 343664
rect 62028 342320 62080 342372
rect 163688 342320 163740 342372
rect 93676 342252 93728 342304
rect 252652 342252 252704 342304
rect 130016 340960 130068 341012
rect 166264 340960 166316 341012
rect 102784 340892 102836 340944
rect 258172 340892 258224 340944
rect 78496 340144 78548 340196
rect 93124 340144 93176 340196
rect 114468 339532 114520 339584
rect 169024 339532 169076 339584
rect 64696 339464 64748 339516
rect 122196 339464 122248 339516
rect 132776 339464 132828 339516
rect 259460 339464 259512 339516
rect 79876 338716 79928 338768
rect 89076 338716 89128 338768
rect 67732 338512 67784 338564
rect 72424 338512 72476 338564
rect 148416 338172 148468 338224
rect 155224 338172 155276 338224
rect 106464 338104 106516 338156
rect 184296 338104 184348 338156
rect 115940 336812 115992 336864
rect 247040 336812 247092 336864
rect 67272 336744 67324 336796
rect 206376 336744 206428 336796
rect 61844 335384 61896 335436
rect 115296 335384 115348 335436
rect 127072 335384 127124 335436
rect 182916 335384 182968 335436
rect 73160 335316 73212 335368
rect 192484 335316 192536 335368
rect 76472 334636 76524 334688
rect 87052 334636 87104 334688
rect 3424 334568 3476 334620
rect 11704 334568 11756 334620
rect 67824 334568 67876 334620
rect 115204 334568 115256 334620
rect 141332 334024 141384 334076
rect 171784 334024 171836 334076
rect 101496 333956 101548 334008
rect 159548 333956 159600 334008
rect 66168 333344 66220 333396
rect 74540 333344 74592 333396
rect 75736 333208 75788 333260
rect 101404 333208 101456 333260
rect 97264 332664 97316 332716
rect 170404 332664 170456 332716
rect 115664 332596 115716 332648
rect 198096 332596 198148 332648
rect 60464 331848 60516 331900
rect 122104 331848 122156 331900
rect 133788 331304 133840 331356
rect 195428 331304 195480 331356
rect 72240 331236 72292 331288
rect 215944 331236 215996 331288
rect 59268 331168 59320 331220
rect 99380 331168 99432 331220
rect 80704 331100 80756 331152
rect 81348 331100 81400 331152
rect 82728 331100 82780 331152
rect 83464 331100 83516 331152
rect 85580 331100 85632 331152
rect 86592 331100 86644 331152
rect 114376 331100 114428 331152
rect 114744 331100 114796 331152
rect 126980 331100 127032 331152
rect 127900 331100 127952 331152
rect 137836 331100 137888 331152
rect 139400 331100 139452 331152
rect 70676 330760 70728 330812
rect 73804 330760 73856 330812
rect 122104 330556 122156 330608
rect 137284 330556 137336 330608
rect 17224 330488 17276 330540
rect 59268 330488 59320 330540
rect 96436 330488 96488 330540
rect 124864 330488 124916 330540
rect 178776 330488 178828 330540
rect 228364 330488 228416 330540
rect 98552 330352 98604 330404
rect 99288 330352 99340 330404
rect 77944 330216 77996 330268
rect 78588 330216 78640 330268
rect 79416 330216 79468 330268
rect 79968 330216 80020 330268
rect 117780 330216 117832 330268
rect 118608 330216 118660 330268
rect 110604 330080 110656 330132
rect 111708 330080 111760 330132
rect 92848 330012 92900 330064
rect 93768 330012 93820 330064
rect 74172 329944 74224 329996
rect 76564 329944 76616 329996
rect 95792 329944 95844 329996
rect 96528 329944 96580 329996
rect 113640 329944 113692 329996
rect 114468 329944 114520 329996
rect 147588 329944 147640 329996
rect 177304 329944 177356 329996
rect 132684 329876 132736 329928
rect 44088 329808 44140 329860
rect 69112 329808 69164 329860
rect 99380 329808 99432 329860
rect 100116 329808 100168 329860
rect 104164 329808 104216 329860
rect 105544 329808 105596 329860
rect 108580 329808 108632 329860
rect 108948 329808 109000 329860
rect 131488 329808 131540 329860
rect 132408 329808 132460 329860
rect 134156 329808 134208 329860
rect 135168 329808 135220 329860
rect 135260 329808 135312 329860
rect 135812 329808 135864 329860
rect 136916 329876 136968 329928
rect 137928 329876 137980 329928
rect 143540 329876 143592 329928
rect 140688 329808 140740 329860
rect 141424 329808 141476 329860
rect 153292 329808 153344 329860
rect 159364 329808 159416 329860
rect 122196 329740 122248 329792
rect 133788 329740 133840 329792
rect 166908 329128 166960 329180
rect 179420 329128 179472 329180
rect 188528 329128 188580 329180
rect 211896 329128 211948 329180
rect 241244 329128 241296 329180
rect 306380 329128 306432 329180
rect 36544 329060 36596 329112
rect 49608 329060 49660 329112
rect 135260 329060 135312 329112
rect 150348 329060 150400 329112
rect 248604 329060 248656 329112
rect 144828 328448 144880 328500
rect 158168 328448 158220 328500
rect 115296 328380 115348 328432
rect 141976 328380 142028 328432
rect 67364 327768 67416 327820
rect 91744 327768 91796 327820
rect 65892 327700 65944 327752
rect 133880 327700 133932 327752
rect 179420 327700 179472 327752
rect 192852 327700 192904 327752
rect 148600 327224 148652 327276
rect 152924 327224 152976 327276
rect 152096 327156 152148 327208
rect 160836 327156 160888 327208
rect 135536 327088 135588 327140
rect 249800 327088 249852 327140
rect 55956 327020 56008 327072
rect 56508 327020 56560 327072
rect 93860 327020 93912 327072
rect 143540 327020 143592 327072
rect 154856 327020 154908 327072
rect 69940 326952 69992 327004
rect 71044 326952 71096 327004
rect 152924 326884 152976 326936
rect 154304 326884 154356 326936
rect 155224 326884 155276 326936
rect 20 326340 72 326392
rect 55956 326340 56008 326392
rect 159640 326408 159692 326460
rect 199384 326408 199436 326460
rect 196716 326340 196768 326392
rect 203524 326340 203576 326392
rect 228456 326340 228508 326392
rect 156052 326000 156104 326052
rect 159456 326000 159508 326052
rect 156144 324980 156196 325032
rect 255504 324980 255556 325032
rect 181628 324912 181680 324964
rect 313924 324912 313976 324964
rect 59268 324300 59320 324352
rect 66812 324300 66864 324352
rect 159548 323620 159600 323672
rect 220820 323620 220872 323672
rect 160928 323552 160980 323604
rect 349160 323552 349212 323604
rect 61936 322940 61988 322992
rect 66812 322940 66864 322992
rect 156052 322940 156104 322992
rect 161020 322940 161072 322992
rect 230480 322464 230532 322516
rect 236736 322464 236788 322516
rect 185768 322260 185820 322312
rect 202880 322260 202932 322312
rect 166264 322192 166316 322244
rect 232504 322192 232556 322244
rect 156052 321580 156104 321632
rect 166448 321580 166500 321632
rect 193864 320900 193916 320952
rect 235264 320900 235316 320952
rect 156972 320832 157024 320884
rect 233884 320832 233936 320884
rect 157248 319948 157300 320000
rect 161572 319948 161624 320000
rect 162216 319948 162268 320000
rect 4068 319404 4120 319456
rect 15844 319404 15896 319456
rect 171784 319404 171836 319456
rect 248512 319404 248564 319456
rect 56508 318792 56560 318844
rect 66260 318792 66312 318844
rect 157248 318792 157300 318844
rect 178868 318792 178920 318844
rect 215852 318724 215904 318776
rect 216036 318724 216088 318776
rect 166356 318112 166408 318164
rect 202788 318112 202840 318164
rect 11704 318044 11756 318096
rect 46848 318044 46900 318096
rect 184204 318044 184256 318096
rect 227076 318044 227128 318096
rect 60648 317500 60700 317552
rect 66260 317500 66312 317552
rect 46848 317432 46900 317484
rect 66352 317432 66404 317484
rect 215852 317432 215904 317484
rect 300952 317432 301004 317484
rect 157248 316684 157300 316736
rect 189816 316684 189868 316736
rect 156696 316004 156748 316056
rect 254032 316004 254084 316056
rect 61844 315936 61896 315988
rect 66996 315936 67048 315988
rect 157248 315936 157300 315988
rect 167000 315936 167052 315988
rect 236736 315324 236788 315376
rect 242900 315324 242952 315376
rect 167000 315256 167052 315308
rect 178776 315256 178828 315308
rect 178868 315256 178920 315308
rect 245752 315256 245804 315308
rect 35256 314644 35308 314696
rect 66444 314644 66496 314696
rect 61844 314168 61896 314220
rect 66260 314168 66312 314220
rect 195428 313896 195480 313948
rect 225052 313896 225104 313948
rect 60556 313216 60608 313268
rect 66260 313216 66312 313268
rect 52276 312536 52328 312588
rect 61108 312536 61160 312588
rect 157156 312536 157208 312588
rect 244280 312536 244332 312588
rect 157248 311856 157300 311908
rect 193864 311856 193916 311908
rect 207572 311856 207624 311908
rect 282184 311856 282236 311908
rect 62028 311788 62080 311840
rect 66812 311788 66864 311840
rect 181536 311176 181588 311228
rect 230480 311176 230532 311228
rect 161020 311108 161072 311160
rect 210516 311108 210568 311160
rect 218704 311108 218756 311160
rect 309140 311108 309192 311160
rect 157248 310496 157300 310548
rect 166356 310496 166408 310548
rect 201684 310360 201736 310412
rect 202144 310360 202196 310412
rect 160836 309748 160888 309800
rect 244556 309748 244608 309800
rect 67088 309408 67140 309460
rect 67456 309408 67508 309460
rect 53564 309136 53616 309188
rect 66628 309136 66680 309188
rect 157156 309136 157208 309188
rect 177580 309136 177632 309188
rect 201684 309136 201736 309188
rect 580264 309136 580316 309188
rect 157248 309068 157300 309120
rect 172520 309068 172572 309120
rect 173808 309068 173860 309120
rect 214656 309068 214708 309120
rect 215208 309068 215260 309120
rect 231216 309068 231268 309120
rect 236736 309068 236788 309120
rect 49608 308388 49660 308440
rect 67088 308388 67140 308440
rect 173808 308388 173860 308440
rect 187056 308388 187108 308440
rect 18604 307776 18656 307828
rect 49608 307776 49660 307828
rect 215208 307776 215260 307828
rect 273904 307776 273956 307828
rect 65892 307708 65944 307760
rect 67088 307708 67140 307760
rect 39304 307028 39356 307080
rect 67180 307028 67232 307080
rect 164976 306892 165028 306944
rect 171784 306892 171836 306944
rect 232504 306416 232556 306468
rect 271144 306416 271196 306468
rect 173164 306348 173216 306400
rect 247316 306348 247368 306400
rect 3424 306280 3476 306332
rect 36544 306280 36596 306332
rect 157248 306280 157300 306332
rect 160100 306280 160152 306332
rect 233976 305804 234028 305856
rect 234528 305804 234580 305856
rect 170404 305600 170456 305652
rect 192668 305600 192720 305652
rect 191104 305260 191156 305312
rect 191656 305260 191708 305312
rect 157248 305192 157300 305244
rect 162124 305192 162176 305244
rect 234528 305056 234580 305108
rect 287336 305056 287388 305108
rect 191656 304988 191708 305040
rect 261576 304988 261628 305040
rect 160100 304240 160152 304292
rect 181628 304240 181680 304292
rect 222844 304240 222896 304292
rect 232504 304240 232556 304292
rect 238668 304240 238720 304292
rect 299572 304240 299624 304292
rect 156052 303628 156104 303680
rect 204996 303628 205048 303680
rect 206376 303628 206428 303680
rect 207020 303628 207072 303680
rect 256700 303628 256752 303680
rect 163596 302880 163648 302932
rect 176108 302880 176160 302932
rect 222936 302268 222988 302320
rect 223488 302268 223540 302320
rect 261484 302268 261536 302320
rect 157248 302200 157300 302252
rect 165528 302200 165580 302252
rect 167644 302200 167696 302252
rect 255596 302200 255648 302252
rect 64696 302132 64748 302184
rect 66812 302132 66864 302184
rect 199384 302132 199436 302184
rect 200580 302132 200632 302184
rect 170496 300908 170548 300960
rect 241428 300908 241480 300960
rect 200120 300840 200172 300892
rect 200580 300840 200632 300892
rect 269948 300840 270000 300892
rect 64604 300772 64656 300824
rect 66812 300772 66864 300824
rect 162216 300092 162268 300144
rect 225972 300092 226024 300144
rect 184204 299548 184256 299600
rect 253204 299548 253256 299600
rect 58900 299480 58952 299532
rect 66444 299480 66496 299532
rect 227076 299480 227128 299532
rect 228916 299480 228968 299532
rect 303620 299480 303672 299532
rect 157248 299140 157300 299192
rect 164148 299140 164200 299192
rect 155224 298800 155276 298852
rect 173348 298800 173400 298852
rect 165528 298732 165580 298784
rect 246396 298732 246448 298784
rect 200212 298120 200264 298172
rect 202880 298120 202932 298172
rect 209044 298120 209096 298172
rect 209412 298120 209464 298172
rect 265624 298120 265676 298172
rect 246304 297440 246356 297492
rect 254124 297440 254176 297492
rect 202880 297372 202932 297424
rect 295340 297372 295392 297424
rect 164976 297304 165028 297356
rect 165712 297304 165764 297356
rect 64696 296692 64748 296744
rect 66628 296692 66680 296744
rect 191104 296692 191156 296744
rect 245108 296692 245160 296744
rect 53748 296624 53800 296676
rect 66444 296624 66496 296676
rect 155224 296012 155276 296064
rect 175280 296012 175332 296064
rect 240784 296012 240836 296064
rect 156420 295944 156472 295996
rect 244464 295944 244516 295996
rect 245108 295944 245160 295996
rect 259552 295944 259604 295996
rect 156328 295264 156380 295316
rect 172704 295264 172756 295316
rect 173808 295264 173860 295316
rect 173808 294652 173860 294704
rect 197360 294652 197412 294704
rect 193864 294584 193916 294636
rect 245844 294584 245896 294636
rect 61752 294040 61804 294092
rect 66812 294040 66864 294092
rect 15844 293972 15896 294024
rect 67548 293972 67600 294024
rect 200028 293972 200080 294024
rect 222200 293972 222252 294024
rect 227812 293972 227864 294024
rect 228456 293972 228508 294024
rect 278044 293972 278096 294024
rect 59176 293904 59228 293956
rect 66812 293904 66864 293956
rect 238116 293904 238168 293956
rect 240508 293904 240560 293956
rect 204996 293224 205048 293276
rect 236000 293224 236052 293276
rect 2780 292816 2832 292868
rect 4804 292816 4856 292868
rect 156512 292612 156564 292664
rect 166264 292612 166316 292664
rect 157248 292544 157300 292596
rect 220176 292544 220228 292596
rect 231124 292544 231176 292596
rect 233148 292544 233200 292596
rect 583392 292544 583444 292596
rect 14464 292476 14516 292528
rect 60464 292476 60516 292528
rect 66904 292476 66956 292528
rect 197360 291796 197412 291848
rect 209044 291796 209096 291848
rect 222476 291660 222528 291712
rect 223028 291660 223080 291712
rect 223028 291252 223080 291304
rect 253940 291252 253992 291304
rect 156052 291184 156104 291236
rect 193864 291184 193916 291236
rect 204996 291184 205048 291236
rect 218612 291184 218664 291236
rect 236092 291184 236144 291236
rect 236644 291184 236696 291236
rect 306564 291184 306616 291236
rect 63316 289892 63368 289944
rect 66812 289892 66864 289944
rect 199476 289892 199528 289944
rect 256884 289892 256936 289944
rect 157248 289824 157300 289876
rect 247408 289824 247460 289876
rect 238024 289076 238076 289128
rect 242348 289076 242400 289128
rect 157248 288464 157300 288516
rect 224500 288464 224552 288516
rect 242348 288464 242400 288516
rect 280160 288464 280212 288516
rect 171232 288396 171284 288448
rect 244372 288396 244424 288448
rect 180340 287104 180392 287156
rect 223580 287104 223632 287156
rect 230756 287104 230808 287156
rect 52184 287036 52236 287088
rect 66628 287036 66680 287088
rect 157248 287036 157300 287088
rect 231308 287036 231360 287088
rect 233884 287104 233936 287156
rect 244188 287104 244240 287156
rect 255320 287036 255372 287088
rect 224224 286356 224276 286408
rect 229284 286356 229336 286408
rect 230112 286356 230164 286408
rect 163596 286288 163648 286340
rect 191196 286288 191248 286340
rect 210424 286220 210476 286272
rect 211436 286220 211488 286272
rect 220084 285880 220136 285932
rect 198832 285744 198884 285796
rect 205548 285744 205600 285796
rect 55128 285676 55180 285728
rect 66812 285676 66864 285728
rect 199384 285676 199436 285728
rect 204628 285676 204680 285728
rect 204904 285676 204956 285728
rect 208124 285676 208176 285728
rect 211804 285676 211856 285728
rect 213828 285676 213880 285728
rect 220728 285676 220780 285728
rect 222108 285676 222160 285728
rect 237564 285812 237616 285864
rect 238668 285812 238720 285864
rect 230112 285744 230164 285796
rect 246120 285744 246172 285796
rect 269764 285676 269816 285728
rect 200120 285268 200172 285320
rect 200948 285268 201000 285320
rect 222200 285268 222252 285320
rect 222660 285268 222712 285320
rect 57796 284928 57848 284980
rect 65524 284928 65576 284980
rect 159548 284384 159600 284436
rect 216772 284384 216824 284436
rect 230480 284384 230532 284436
rect 231676 284384 231728 284436
rect 281908 284384 281960 284436
rect 156420 284316 156472 284368
rect 243912 284316 243964 284368
rect 191196 283908 191248 283960
rect 201408 283908 201460 283960
rect 244188 283840 244240 283892
rect 282920 283840 282972 283892
rect 162124 283568 162176 283620
rect 188988 283568 189040 283620
rect 157248 283160 157300 283212
rect 162768 283160 162820 283212
rect 246304 283160 246356 283212
rect 247040 283160 247092 283212
rect 250076 283160 250128 283212
rect 245936 282820 245988 282872
rect 254124 282820 254176 282872
rect 582748 282820 582800 282872
rect 162768 282140 162820 282192
rect 184848 282140 184900 282192
rect 185032 282140 185084 282192
rect 197084 282140 197136 282192
rect 60556 281528 60608 281580
rect 66812 281528 66864 281580
rect 184848 281528 184900 281580
rect 197360 281528 197412 281580
rect 157248 281460 157300 281512
rect 184204 281460 184256 281512
rect 181628 281392 181680 281444
rect 197360 281392 197412 281444
rect 156880 280780 156932 280832
rect 171232 280780 171284 280832
rect 245936 280780 245988 280832
rect 248604 280780 248656 280832
rect 311992 280780 312044 280832
rect 63224 280168 63276 280220
rect 66812 280168 66864 280220
rect 245476 280168 245528 280220
rect 273996 280168 274048 280220
rect 195428 279692 195480 279744
rect 198740 279692 198792 279744
rect 158168 279624 158220 279676
rect 162216 279624 162268 279676
rect 157248 279488 157300 279540
rect 158720 279488 158772 279540
rect 171876 279420 171928 279472
rect 245936 279420 245988 279472
rect 251272 279420 251324 279472
rect 245660 278944 245712 278996
rect 247316 278944 247368 278996
rect 192576 278808 192628 278860
rect 197360 278808 197412 278860
rect 11704 278740 11756 278792
rect 59084 278740 59136 278792
rect 67180 278740 67232 278792
rect 251272 278740 251324 278792
rect 583208 278740 583260 278792
rect 191656 278672 191708 278724
rect 197360 278672 197412 278724
rect 157064 278060 157116 278112
rect 170588 278060 170640 278112
rect 180248 278060 180300 278112
rect 198832 278060 198884 278112
rect 245936 278060 245988 278112
rect 249800 278060 249852 278112
rect 158168 277992 158220 278044
rect 185032 277992 185084 278044
rect 246028 277992 246080 278044
rect 249984 277992 250036 278044
rect 583300 277992 583352 278044
rect 57704 277380 57756 277432
rect 66444 277380 66496 277432
rect 157340 276700 157392 276752
rect 197360 276700 197412 276752
rect 199384 276632 199436 276684
rect 245752 276632 245804 276684
rect 278136 276632 278188 276684
rect 155316 276564 155368 276616
rect 53472 276020 53524 276072
rect 66812 276020 66864 276072
rect 245936 275952 245988 276004
rect 254032 275952 254084 276004
rect 582656 275952 582708 276004
rect 157248 275272 157300 275324
rect 173256 275272 173308 275324
rect 160928 274728 160980 274780
rect 197360 274728 197412 274780
rect 56416 274660 56468 274712
rect 66812 274660 66864 274712
rect 157248 274660 157300 274712
rect 161020 274660 161072 274712
rect 156512 274592 156564 274644
rect 191104 274592 191156 274644
rect 196716 274524 196768 274576
rect 200028 274524 200080 274576
rect 182916 273912 182968 273964
rect 195520 273912 195572 273964
rect 62028 273232 62080 273284
rect 66812 273232 66864 273284
rect 245660 273232 245712 273284
rect 254032 273232 254084 273284
rect 176568 273164 176620 273216
rect 197360 273164 197412 273216
rect 185584 273096 185636 273148
rect 197452 273096 197504 273148
rect 260104 272484 260156 272536
rect 302240 272484 302292 272536
rect 63132 271872 63184 271924
rect 66812 271872 66864 271924
rect 245844 271872 245896 271924
rect 251272 271872 251324 271924
rect 259460 271872 259512 271924
rect 156972 271124 157024 271176
rect 191380 271124 191432 271176
rect 48228 270512 48280 270564
rect 66812 270512 66864 270564
rect 166448 270512 166500 270564
rect 197452 270512 197504 270564
rect 245844 270512 245896 270564
rect 252836 270512 252888 270564
rect 164240 270444 164292 270496
rect 197360 270444 197412 270496
rect 256792 270444 256844 270496
rect 583024 270444 583076 270496
rect 163688 270240 163740 270292
rect 164240 270240 164292 270292
rect 246304 269832 246356 269884
rect 247040 269832 247092 269884
rect 252652 269832 252704 269884
rect 4068 269764 4120 269816
rect 21456 269764 21508 269816
rect 245844 269764 245896 269816
rect 256792 269764 256844 269816
rect 181628 269560 181680 269612
rect 186320 269560 186372 269612
rect 64512 269084 64564 269136
rect 66812 269084 66864 269136
rect 157248 269084 157300 269136
rect 178960 269084 179012 269136
rect 21088 269016 21140 269068
rect 22744 269016 22796 269068
rect 67364 269016 67416 269068
rect 67640 269016 67692 269068
rect 156420 269016 156472 269068
rect 180340 269016 180392 269068
rect 245752 269016 245804 269068
rect 255412 269016 255464 269068
rect 178776 268948 178828 269000
rect 197360 268948 197412 269000
rect 55036 268336 55088 268388
rect 66996 268336 67048 268388
rect 180064 268336 180116 268388
rect 197360 268336 197412 268388
rect 255412 268336 255464 268388
rect 582656 268336 582708 268388
rect 195244 267112 195296 267164
rect 197452 267112 197504 267164
rect 3424 266976 3476 267028
rect 21364 266976 21416 267028
rect 245844 266976 245896 267028
rect 288532 266976 288584 267028
rect 64788 266500 64840 266552
rect 66168 266500 66220 266552
rect 66628 266500 66680 266552
rect 173532 266432 173584 266484
rect 197360 266432 197412 266484
rect 157248 266364 157300 266416
rect 184204 266364 184256 266416
rect 245936 266364 245988 266416
rect 263600 266364 263652 266416
rect 245936 265616 245988 265668
rect 251364 265616 251416 265668
rect 263692 265616 263744 265668
rect 583024 265616 583076 265668
rect 41144 264936 41196 264988
rect 66812 264936 66864 264988
rect 157248 264936 157300 264988
rect 171968 264936 172020 264988
rect 186136 264936 186188 264988
rect 197360 264936 197412 264988
rect 188344 264868 188396 264920
rect 197452 264868 197504 264920
rect 41328 264188 41380 264240
rect 58992 264188 59044 264240
rect 66812 264188 66864 264240
rect 166356 264188 166408 264240
rect 187240 264188 187292 264240
rect 246488 264188 246540 264240
rect 299664 264188 299716 264240
rect 245844 263984 245896 264036
rect 248420 263984 248472 264036
rect 60464 263576 60516 263628
rect 66720 263576 66772 263628
rect 195244 263576 195296 263628
rect 197360 263576 197412 263628
rect 52368 262828 52420 262880
rect 66812 262828 66864 262880
rect 251364 262828 251416 262880
rect 259460 262828 259512 262880
rect 156420 262284 156472 262336
rect 170404 262284 170456 262336
rect 159640 262216 159692 262268
rect 195244 262216 195296 262268
rect 164240 262148 164292 262200
rect 169760 262148 169812 262200
rect 161020 261536 161072 261588
rect 177580 261536 177632 261588
rect 186964 261536 187016 261588
rect 197360 261536 197412 261588
rect 246396 261536 246448 261588
rect 247408 261536 247460 261588
rect 248420 261536 248472 261588
rect 21456 261468 21508 261520
rect 63500 261468 63552 261520
rect 173348 261468 173400 261520
rect 199476 261468 199528 261520
rect 265716 261468 265768 261520
rect 580356 261468 580408 261520
rect 63500 260924 63552 260976
rect 64788 260924 64840 260976
rect 66812 260924 66864 260976
rect 157248 260856 157300 260908
rect 164240 260856 164292 260908
rect 156972 260788 157024 260840
rect 177488 260788 177540 260840
rect 245752 260720 245804 260772
rect 251456 260720 251508 260772
rect 156328 260108 156380 260160
rect 179052 260108 179104 260160
rect 253204 259496 253256 259548
rect 276664 259496 276716 259548
rect 178960 259428 179012 259480
rect 182180 259428 182232 259480
rect 193956 259428 194008 259480
rect 197360 259428 197412 259480
rect 244464 259428 244516 259480
rect 291200 259428 291252 259480
rect 169116 259360 169168 259412
rect 197452 259360 197504 259412
rect 245936 259360 245988 259412
rect 253204 259360 253256 259412
rect 264244 259360 264296 259412
rect 579804 259360 579856 259412
rect 184296 259292 184348 259344
rect 184756 259292 184808 259344
rect 184756 258680 184808 258732
rect 197360 258680 197412 258732
rect 53748 258068 53800 258120
rect 66260 258068 66312 258120
rect 245844 258068 245896 258120
rect 279424 258068 279476 258120
rect 245660 258000 245712 258052
rect 255596 258000 255648 258052
rect 156880 257932 156932 257984
rect 159548 257932 159600 257984
rect 157248 257320 157300 257372
rect 192576 257320 192628 257372
rect 255596 257320 255648 257372
rect 271236 257320 271288 257372
rect 162768 256708 162820 256760
rect 177948 256708 178000 256760
rect 197452 256708 197504 256760
rect 189816 256640 189868 256692
rect 197360 256640 197412 256692
rect 245936 256572 245988 256624
rect 259552 256572 259604 256624
rect 260748 256572 260800 256624
rect 178684 256164 178736 256216
rect 182916 256164 182968 256216
rect 155224 255960 155276 256012
rect 186964 255960 187016 256012
rect 260748 255960 260800 256012
rect 296720 255960 296772 256012
rect 64604 255280 64656 255332
rect 66812 255280 66864 255332
rect 191104 255280 191156 255332
rect 195428 255280 195480 255332
rect 3424 255212 3476 255264
rect 18604 255212 18656 255264
rect 245844 255212 245896 255264
rect 255504 255212 255556 255264
rect 245936 255144 245988 255196
rect 249800 255144 249852 255196
rect 157248 254600 157300 254652
rect 161664 254600 161716 254652
rect 162676 254600 162728 254652
rect 156512 254532 156564 254584
rect 173808 254532 173860 254584
rect 187700 254532 187752 254584
rect 188804 254532 188856 254584
rect 198004 254532 198056 254584
rect 56324 253920 56376 253972
rect 66812 253920 66864 253972
rect 162124 253920 162176 253972
rect 163688 253920 163740 253972
rect 165068 253920 165120 253972
rect 187700 253920 187752 253972
rect 193036 253920 193088 253972
rect 197360 253920 197412 253972
rect 54944 253852 54996 253904
rect 57152 253852 57204 253904
rect 245936 253852 245988 253904
rect 256884 253852 256936 253904
rect 157248 253580 157300 253632
rect 162768 253580 162820 253632
rect 54944 253172 54996 253224
rect 66904 253172 66956 253224
rect 160744 253172 160796 253224
rect 168380 253172 168432 253224
rect 256884 253172 256936 253224
rect 294052 253172 294104 253224
rect 187608 252628 187660 252680
rect 197360 252628 197412 252680
rect 57152 252560 57204 252612
rect 57612 252560 57664 252612
rect 66812 252560 66864 252612
rect 168380 252560 168432 252612
rect 169576 252560 169628 252612
rect 197452 252560 197504 252612
rect 245844 252492 245896 252544
rect 262220 252492 262272 252544
rect 262680 252492 262732 252544
rect 245936 252288 245988 252340
rect 248696 252288 248748 252340
rect 173808 251812 173860 251864
rect 187700 251812 187752 251864
rect 262680 251812 262732 251864
rect 583576 251812 583628 251864
rect 157248 251268 157300 251320
rect 169760 251268 169812 251320
rect 157156 251200 157208 251252
rect 180064 251200 180116 251252
rect 187700 251200 187752 251252
rect 188896 251200 188948 251252
rect 197360 251200 197412 251252
rect 245660 250520 245712 250572
rect 269856 250520 269908 250572
rect 170588 250452 170640 250504
rect 180340 250452 180392 250504
rect 185676 250452 185728 250504
rect 197084 250452 197136 250504
rect 265624 250452 265676 250504
rect 289820 250452 289872 250504
rect 60372 249772 60424 249824
rect 66444 249772 66496 249824
rect 157248 249772 157300 249824
rect 186964 249772 187016 249824
rect 191196 249772 191248 249824
rect 197360 249772 197412 249824
rect 192668 249704 192720 249756
rect 195888 249704 195940 249756
rect 191380 249636 191432 249688
rect 193128 249636 193180 249688
rect 197360 249636 197412 249688
rect 245936 249636 245988 249688
rect 249892 249636 249944 249688
rect 156972 249364 157024 249416
rect 159640 249364 159692 249416
rect 169024 249024 169076 249076
rect 191288 249024 191340 249076
rect 195888 248684 195940 248736
rect 197360 248684 197412 248736
rect 156512 248412 156564 248464
rect 172520 248412 172572 248464
rect 156236 247664 156288 247716
rect 164976 247664 165028 247716
rect 185860 247664 185912 247716
rect 199568 247664 199620 247716
rect 245936 247664 245988 247716
rect 582840 247664 582892 247716
rect 50988 247052 51040 247104
rect 66812 247052 66864 247104
rect 164148 247052 164200 247104
rect 185860 247052 185912 247104
rect 186228 247052 186280 247104
rect 187148 247052 187200 247104
rect 197360 247052 197412 247104
rect 171968 246304 172020 246356
rect 189816 246304 189868 246356
rect 157248 246032 157300 246084
rect 160836 246032 160888 246084
rect 246396 245692 246448 245744
rect 247224 245692 247276 245744
rect 158260 245624 158312 245676
rect 191748 245624 191800 245676
rect 197360 245624 197412 245676
rect 245844 245624 245896 245676
rect 248604 245624 248656 245676
rect 298192 245624 298244 245676
rect 53656 244876 53708 244928
rect 66076 244876 66128 244928
rect 66628 244876 66680 244928
rect 245936 244400 245988 244452
rect 248696 244400 248748 244452
rect 157984 244332 158036 244384
rect 193404 244332 193456 244384
rect 155684 244264 155736 244316
rect 198832 244264 198884 244316
rect 192484 244128 192536 244180
rect 197176 244128 197228 244180
rect 197452 244128 197504 244180
rect 193404 243584 193456 243636
rect 197360 243584 197412 243636
rect 154948 243516 155000 243568
rect 164240 243516 164292 243568
rect 164976 243516 165028 243568
rect 172520 243516 172572 243568
rect 194048 243516 194100 243568
rect 63408 242904 63460 242956
rect 66812 242904 66864 242956
rect 156052 242904 156104 242956
rect 192668 242904 192720 242956
rect 244464 242904 244516 242956
rect 244648 242904 244700 242956
rect 265624 242904 265676 242956
rect 64512 242156 64564 242208
rect 82820 242020 82872 242072
rect 152464 242020 152516 242072
rect 164148 242224 164200 242276
rect 269948 242224 270000 242276
rect 285680 242224 285732 242276
rect 168380 242156 168432 242208
rect 169668 242156 169720 242208
rect 197360 242156 197412 242208
rect 245108 242156 245160 242208
rect 252744 242156 252796 242208
rect 261576 242156 261628 242208
rect 278228 242156 278280 242208
rect 154120 242020 154172 242072
rect 165068 242020 165120 242072
rect 70400 241816 70452 241868
rect 71044 241816 71096 241868
rect 149152 241544 149204 241596
rect 154028 241544 154080 241596
rect 163688 241476 163740 241528
rect 191656 241476 191708 241528
rect 195336 241476 195388 241528
rect 197544 241476 197596 241528
rect 245936 241476 245988 241528
rect 255504 241476 255556 241528
rect 141470 241408 141522 241460
rect 149060 241408 149112 241460
rect 193864 241408 193916 241460
rect 197360 241408 197412 241460
rect 3424 241068 3476 241120
rect 7564 241068 7616 241120
rect 115848 240796 115900 240848
rect 155684 240796 155736 240848
rect 65984 240728 66036 240780
rect 76656 240728 76708 240780
rect 82820 240728 82872 240780
rect 128820 240728 128872 240780
rect 149520 240728 149572 240780
rect 199568 240728 199620 240780
rect 198740 240320 198792 240372
rect 200120 240252 200172 240304
rect 67824 240116 67876 240168
rect 76564 240116 76616 240168
rect 104900 240116 104952 240168
rect 105452 240116 105504 240168
rect 198648 240116 198700 240168
rect 200120 240116 200172 240168
rect 200304 240116 200356 240168
rect 202144 240116 202196 240168
rect 242256 240116 242308 240168
rect 244096 240116 244148 240168
rect 67548 240048 67600 240100
rect 69756 240048 69808 240100
rect 70308 240048 70360 240100
rect 115848 240048 115900 240100
rect 117228 240048 117280 240100
rect 224316 240048 224368 240100
rect 240876 240048 240928 240100
rect 243912 240048 243964 240100
rect 79048 239980 79100 240032
rect 79876 239980 79928 240032
rect 80520 239980 80572 240032
rect 81348 239980 81400 240032
rect 81532 239980 81584 240032
rect 82728 239980 82780 240032
rect 86040 239980 86092 240032
rect 86868 239980 86920 240032
rect 90456 239980 90508 240032
rect 90916 239980 90968 240032
rect 121736 239980 121788 240032
rect 122748 239980 122800 240032
rect 127440 239980 127492 240032
rect 128268 239980 128320 240032
rect 131856 239980 131908 240032
rect 132316 239980 132368 240032
rect 128912 239912 128964 239964
rect 129648 239912 129700 239964
rect 126152 239844 126204 239896
rect 228732 239980 228784 240032
rect 240048 239980 240100 240032
rect 252836 240048 252888 240100
rect 138112 239912 138164 239964
rect 138940 239912 138992 239964
rect 142252 239912 142304 239964
rect 143356 239912 143408 239964
rect 145288 239912 145340 239964
rect 146024 239912 146076 239964
rect 106832 239776 106884 239828
rect 107568 239776 107620 239828
rect 148232 239776 148284 239828
rect 148968 239776 149020 239828
rect 101128 239640 101180 239692
rect 102048 239640 102100 239692
rect 120172 239640 120224 239692
rect 121368 239640 121420 239692
rect 88984 239504 89036 239556
rect 89536 239504 89588 239556
rect 99380 239504 99432 239556
rect 100668 239504 100720 239556
rect 107752 239504 107804 239556
rect 108396 239504 108448 239556
rect 109592 239504 109644 239556
rect 110236 239504 110288 239556
rect 111064 239504 111116 239556
rect 111616 239504 111668 239556
rect 71688 239368 71740 239420
rect 79324 239368 79376 239420
rect 124680 239368 124732 239420
rect 125416 239368 125468 239420
rect 97632 239300 97684 239352
rect 104164 239300 104216 239352
rect 115296 239232 115348 239284
rect 115848 239232 115900 239284
rect 130384 239232 130436 239284
rect 130936 239232 130988 239284
rect 133144 239164 133196 239216
rect 133696 239164 133748 239216
rect 134616 239164 134668 239216
rect 135168 239164 135220 239216
rect 141056 239096 141108 239148
rect 142068 239096 142120 239148
rect 144000 239096 144052 239148
rect 144736 239096 144788 239148
rect 149060 239096 149112 239148
rect 149612 239096 149664 239148
rect 153936 239096 153988 239148
rect 154488 239096 154540 239148
rect 226892 238756 226944 238808
rect 238944 238756 238996 238808
rect 240048 238756 240100 238808
rect 219440 238688 219492 238740
rect 222844 238688 222896 238740
rect 242164 238688 242216 238740
rect 248512 238688 248564 238740
rect 107660 238620 107712 238672
rect 219900 238620 219952 238672
rect 60372 238076 60424 238128
rect 73804 238076 73856 238128
rect 224316 238076 224368 238128
rect 236644 238076 236696 238128
rect 67916 238008 67968 238060
rect 108304 238008 108356 238060
rect 215300 238008 215352 238060
rect 244464 238008 244516 238060
rect 199476 237804 199528 237856
rect 199936 237804 199988 237856
rect 201040 237804 201092 237856
rect 230572 237804 230624 237856
rect 231768 237804 231820 237856
rect 84200 237668 84252 237720
rect 93124 237668 93176 237720
rect 200120 237396 200172 237448
rect 201592 237396 201644 237448
rect 206836 237396 206888 237448
rect 207664 237396 207716 237448
rect 207940 237396 207992 237448
rect 209044 237396 209096 237448
rect 211252 237396 211304 237448
rect 211804 237396 211856 237448
rect 223028 237396 223080 237448
rect 223764 237396 223816 237448
rect 4804 237328 4856 237380
rect 53840 237328 53892 237380
rect 103520 237328 103572 237380
rect 137100 237328 137152 237380
rect 138020 237328 138072 237380
rect 164884 237328 164936 237380
rect 216036 237328 216088 237380
rect 265716 237328 265768 237380
rect 118700 237260 118752 237312
rect 152464 237260 152516 237312
rect 196900 237260 196952 237312
rect 208860 237260 208912 237312
rect 186964 237192 187016 237244
rect 215300 237192 215352 237244
rect 53840 236648 53892 236700
rect 54852 236648 54904 236700
rect 86224 236648 86276 236700
rect 91100 236648 91152 236700
rect 104256 236648 104308 236700
rect 152464 236648 152516 236700
rect 161480 236648 161532 236700
rect 162768 236648 162820 236700
rect 176016 236648 176068 236700
rect 185584 236648 185636 236700
rect 195888 236444 195940 236496
rect 196808 236444 196860 236496
rect 214656 236104 214708 236156
rect 216036 236104 216088 236156
rect 226984 236036 227036 236088
rect 229652 236036 229704 236088
rect 128820 235900 128872 235952
rect 181628 235900 181680 235952
rect 189908 235900 189960 235952
rect 204444 235900 204496 235952
rect 235356 235900 235408 235952
rect 252928 235900 252980 235952
rect 103704 235288 103756 235340
rect 119436 235288 119488 235340
rect 115940 235220 115992 235272
rect 137284 235220 137336 235272
rect 243636 235220 243688 235272
rect 284300 235220 284352 235272
rect 194692 234676 194744 234728
rect 211068 234676 211120 234728
rect 231124 234676 231176 234728
rect 232044 234676 232096 234728
rect 208400 234608 208452 234660
rect 240324 234608 240376 234660
rect 240784 234608 240836 234660
rect 252928 234608 252980 234660
rect 582840 234608 582892 234660
rect 21364 234540 21416 234592
rect 92480 234540 92532 234592
rect 122932 234540 122984 234592
rect 145932 234540 145984 234592
rect 146024 234540 146076 234592
rect 161020 234540 161072 234592
rect 177580 234540 177632 234592
rect 249892 234540 249944 234592
rect 133604 234472 133656 234524
rect 184388 234472 184440 234524
rect 188804 234472 188856 234524
rect 192484 234472 192536 234524
rect 192668 234472 192720 234524
rect 240968 234472 241020 234524
rect 241244 234472 241296 234524
rect 63224 233860 63276 233912
rect 75184 233860 75236 233912
rect 92480 233860 92532 233912
rect 111064 233860 111116 233912
rect 57704 233180 57756 233232
rect 124312 233180 124364 233232
rect 126704 233180 126756 233232
rect 173348 233180 173400 233232
rect 173532 233180 173584 233232
rect 182916 233180 182968 233232
rect 225236 233180 225288 233232
rect 155500 233112 155552 233164
rect 158260 233112 158312 233164
rect 194048 233112 194100 233164
rect 219532 233112 219584 233164
rect 107752 232500 107804 232552
rect 129004 232500 129056 232552
rect 138112 232500 138164 232552
rect 153108 232500 153160 232552
rect 155316 232500 155368 232552
rect 157340 232500 157392 232552
rect 173808 232500 173860 232552
rect 225604 231820 225656 231872
rect 226156 231820 226208 231872
rect 292580 231820 292632 231872
rect 54944 231752 54996 231804
rect 126244 231752 126296 231804
rect 148876 231752 148928 231804
rect 166448 231752 166500 231804
rect 180340 231752 180392 231804
rect 223028 231752 223080 231804
rect 147588 231684 147640 231736
rect 158168 231684 158220 231736
rect 199568 231684 199620 231736
rect 208400 231684 208452 231736
rect 226708 231140 226760 231192
rect 295432 231140 295484 231192
rect 77392 231072 77444 231124
rect 148508 231072 148560 231124
rect 158260 231072 158312 231124
rect 167644 231072 167696 231124
rect 228732 231072 228784 231124
rect 305184 231072 305236 231124
rect 63132 230392 63184 230444
rect 187700 230460 187752 230512
rect 187240 230392 187292 230444
rect 207664 230392 207716 230444
rect 142068 230324 142120 230376
rect 234068 230324 234120 230376
rect 213184 229712 213236 229764
rect 231952 229712 232004 229764
rect 287152 229712 287204 229764
rect 64788 229032 64840 229084
rect 170496 229032 170548 229084
rect 202144 229032 202196 229084
rect 252744 229032 252796 229084
rect 123024 228964 123076 229016
rect 199384 228964 199436 229016
rect 173256 228896 173308 228948
rect 220452 228896 220504 228948
rect 252744 228352 252796 228404
rect 313372 228352 313424 228404
rect 220084 227740 220136 227792
rect 220452 227740 220504 227792
rect 224224 227740 224276 227792
rect 115756 227672 115808 227724
rect 130384 227672 130436 227724
rect 227260 227740 227312 227792
rect 227812 227740 227864 227792
rect 284392 227740 284444 227792
rect 229744 227672 229796 227724
rect 135168 227060 135220 227112
rect 146760 227060 146812 227112
rect 148508 227060 148560 227112
rect 215944 227060 215996 227112
rect 217140 227060 217192 227112
rect 226340 227060 226392 227112
rect 56324 226992 56376 227044
rect 115204 226992 115256 227044
rect 119436 226992 119488 227044
rect 194968 226992 195020 227044
rect 214104 226992 214156 227044
rect 225604 226992 225656 227044
rect 282184 226992 282236 227044
rect 292672 226992 292724 227044
rect 86224 226244 86276 226296
rect 137376 226244 137428 226296
rect 144736 226244 144788 226296
rect 236828 226312 236880 226364
rect 313280 226312 313332 226364
rect 57796 225564 57848 225616
rect 142896 225564 142948 225616
rect 143356 225564 143408 225616
rect 230388 225564 230440 225616
rect 231124 225564 231176 225616
rect 238300 225564 238352 225616
rect 245844 225564 245896 225616
rect 76656 224884 76708 224936
rect 244280 224884 244332 224936
rect 132316 224204 132368 224256
rect 164884 224204 164936 224256
rect 193036 223592 193088 223644
rect 582472 223592 582524 223644
rect 160008 223524 160060 223576
rect 160928 223524 160980 223576
rect 188068 223524 188120 223576
rect 188804 223524 188856 223576
rect 191104 223524 191156 223576
rect 194968 223524 195020 223576
rect 217508 223524 217560 223576
rect 136548 222912 136600 222964
rect 160008 222912 160060 222964
rect 162216 222912 162268 222964
rect 199476 222912 199528 222964
rect 86960 222844 87012 222896
rect 188068 222844 188120 222896
rect 204996 222844 205048 222896
rect 582748 222844 582800 222896
rect 187700 222096 187752 222148
rect 193036 222096 193088 222148
rect 50528 222028 50580 222080
rect 50804 222028 50856 222080
rect 93860 222028 93912 222080
rect 99472 222028 99524 222080
rect 211252 222028 211304 222080
rect 211804 222028 211856 222080
rect 57612 221960 57664 222012
rect 188436 221960 188488 222012
rect 215944 221484 215996 221536
rect 246304 221484 246356 221536
rect 4804 221416 4856 221468
rect 50528 221416 50580 221468
rect 197084 221416 197136 221468
rect 255412 221416 255464 221468
rect 580908 220940 580960 220992
rect 583208 220940 583260 220992
rect 144828 220736 144880 220788
rect 235264 220736 235316 220788
rect 193036 220668 193088 220720
rect 193956 220668 194008 220720
rect 104992 220056 105044 220108
rect 193036 220056 193088 220108
rect 201500 220056 201552 220108
rect 301044 220056 301096 220108
rect 155408 219376 155460 219428
rect 242900 219376 242952 219428
rect 304264 219376 304316 219428
rect 580172 219376 580224 219428
rect 137928 219308 137980 219360
rect 213184 219308 213236 219360
rect 242900 218764 242952 218816
rect 243912 218764 243964 218816
rect 52184 218696 52236 218748
rect 143356 218696 143408 218748
rect 67732 217948 67784 218000
rect 137468 217948 137520 218000
rect 130936 217880 130988 217932
rect 181536 217880 181588 217932
rect 189080 217336 189132 217388
rect 231860 217336 231912 217388
rect 142896 217268 142948 217320
rect 218060 217268 218112 217320
rect 218980 217268 219032 217320
rect 219440 217268 219492 217320
rect 220268 217268 220320 217320
rect 291384 217268 291436 217320
rect 81624 216588 81676 216640
rect 191288 216588 191340 216640
rect 180064 216520 180116 216572
rect 255504 216520 255556 216572
rect 100668 215908 100720 215960
rect 173164 215908 173216 215960
rect 193956 215908 194008 215960
rect 207388 215908 207440 215960
rect 298744 215908 298796 215960
rect 309324 215908 309376 215960
rect 255504 215296 255556 215348
rect 255964 215296 256016 215348
rect 3332 215228 3384 215280
rect 40684 215228 40736 215280
rect 199384 214616 199436 214668
rect 230572 214616 230624 214668
rect 61752 214548 61804 214600
rect 115296 214548 115348 214600
rect 126888 214548 126940 214600
rect 197360 214548 197412 214600
rect 203340 214548 203392 214600
rect 211160 214548 211212 214600
rect 307944 214548 307996 214600
rect 167644 213936 167696 213988
rect 202972 213936 203024 213988
rect 203616 213936 203668 213988
rect 75184 213868 75236 213920
rect 195336 213868 195388 213920
rect 197360 213868 197412 213920
rect 227812 213868 227864 213920
rect 133880 213800 133932 213852
rect 244372 213800 244424 213852
rect 240968 213188 241020 213240
rect 285772 213188 285824 213240
rect 71044 212440 71096 212492
rect 233516 212440 233568 212492
rect 234436 212440 234488 212492
rect 146208 212372 146260 212424
rect 244556 212372 244608 212424
rect 69020 211080 69072 211132
rect 189080 211080 189132 211132
rect 162308 211012 162360 211064
rect 256792 211012 256844 211064
rect 197912 209788 197964 209840
rect 214472 209788 214524 209840
rect 239404 209788 239456 209840
rect 103428 209108 103480 209160
rect 133144 209108 133196 209160
rect 133696 209108 133748 209160
rect 193864 209108 193916 209160
rect 204904 209108 204956 209160
rect 302516 209108 302568 209160
rect 67640 209040 67692 209092
rect 205548 209040 205600 209092
rect 236644 209040 236696 209092
rect 298744 209040 298796 209092
rect 205548 208836 205600 208888
rect 206468 208836 206520 208888
rect 85580 208292 85632 208344
rect 197912 208292 197964 208344
rect 200028 207680 200080 207732
rect 230480 207680 230532 207732
rect 235264 207680 235316 207732
rect 294144 207680 294196 207732
rect 113088 207612 113140 207664
rect 236276 207612 236328 207664
rect 248696 207612 248748 207664
rect 93124 206932 93176 206984
rect 208308 206932 208360 206984
rect 110236 206864 110288 206916
rect 219440 206864 219492 206916
rect 220728 206864 220780 206916
rect 220728 206252 220780 206304
rect 280252 206252 280304 206304
rect 207848 206116 207900 206168
rect 208308 206116 208360 206168
rect 81348 205572 81400 205624
rect 157340 205572 157392 205624
rect 164884 205572 164936 205624
rect 240140 205572 240192 205624
rect 240876 205572 240928 205624
rect 95240 204892 95292 204944
rect 242992 204892 243044 204944
rect 70400 204212 70452 204264
rect 215484 204212 215536 204264
rect 74540 204144 74592 204196
rect 167644 204144 167696 204196
rect 215484 203600 215536 203652
rect 228548 203600 228600 203652
rect 262864 203600 262916 203652
rect 306656 203600 306708 203652
rect 173164 203532 173216 203584
rect 195428 203532 195480 203584
rect 225604 203532 225656 203584
rect 291292 203532 291344 203584
rect 3424 202784 3476 202836
rect 119436 202784 119488 202836
rect 121368 202784 121420 202836
rect 155224 202784 155276 202836
rect 171784 202172 171836 202224
rect 186964 202172 187016 202224
rect 193128 202172 193180 202224
rect 252652 202172 252704 202224
rect 125508 202104 125560 202156
rect 237380 202104 237432 202156
rect 247132 202104 247184 202156
rect 264244 202104 264296 202156
rect 310612 202104 310664 202156
rect 63316 201424 63368 201476
rect 214656 201424 214708 201476
rect 223028 200812 223080 200864
rect 229100 200812 229152 200864
rect 214932 200200 214984 200252
rect 225696 200200 225748 200252
rect 186136 200132 186188 200184
rect 247684 200132 247736 200184
rect 46848 200064 46900 200116
rect 217416 200064 217468 200116
rect 131028 199996 131080 200048
rect 187056 199996 187108 200048
rect 222108 198772 222160 198824
rect 238116 198772 238168 198824
rect 296904 198704 296956 198756
rect 110328 198636 110380 198688
rect 187608 198636 187660 198688
rect 192576 198636 192628 198688
rect 222108 198636 222160 198688
rect 58900 197956 58952 198008
rect 133788 197956 133840 198008
rect 202236 197956 202288 198008
rect 286324 197956 286376 198008
rect 133788 197276 133840 197328
rect 186136 197276 186188 197328
rect 207848 197276 207900 197328
rect 214932 197276 214984 197328
rect 195244 196664 195296 196716
rect 227076 196664 227128 196716
rect 228364 196664 228416 196716
rect 303804 196664 303856 196716
rect 89536 196596 89588 196648
rect 196900 196596 196952 196648
rect 214564 196596 214616 196648
rect 295616 196596 295668 196648
rect 56416 195916 56468 195968
rect 174636 195916 174688 195968
rect 79968 195848 80020 195900
rect 189264 195848 189316 195900
rect 189264 195304 189316 195356
rect 190368 195304 190420 195356
rect 228364 195304 228416 195356
rect 203616 195236 203668 195288
rect 279056 195236 279108 195288
rect 316684 195236 316736 195288
rect 325700 195236 325752 195288
rect 86868 194488 86920 194540
rect 168380 194488 168432 194540
rect 188896 193876 188948 193928
rect 251824 193876 251876 193928
rect 255964 193876 256016 193928
rect 268476 193876 268528 193928
rect 177948 193808 178000 193860
rect 302332 193808 302384 193860
rect 115204 193128 115256 193180
rect 198004 193128 198056 193180
rect 197268 192516 197320 192568
rect 228456 192516 228508 192568
rect 228640 192516 228692 192568
rect 235356 192516 235408 192568
rect 268384 192516 268436 192568
rect 296812 192516 296864 192568
rect 202788 192448 202840 192500
rect 305276 192448 305328 192500
rect 143448 191768 143500 191820
rect 209228 191768 209280 191820
rect 179328 191700 179380 191752
rect 180248 191700 180300 191752
rect 191288 191156 191340 191208
rect 233976 191156 234028 191208
rect 104900 191088 104952 191140
rect 179328 191088 179380 191140
rect 209044 191088 209096 191140
rect 281816 191088 281868 191140
rect 69664 190408 69716 190460
rect 193956 190408 194008 190460
rect 228548 189796 228600 189848
rect 244464 189796 244516 189848
rect 188988 189728 189040 189780
rect 231952 189728 232004 189780
rect 129648 189048 129700 189100
rect 166264 189048 166316 189100
rect 3516 188980 3568 189032
rect 35256 188980 35308 189032
rect 187056 188368 187108 188420
rect 221372 188368 221424 188420
rect 35164 188300 35216 188352
rect 162124 188300 162176 188352
rect 174636 188300 174688 188352
rect 288624 188300 288676 188352
rect 135168 187688 135220 187740
rect 163504 187688 163556 187740
rect 221372 187008 221424 187060
rect 232136 187008 232188 187060
rect 184848 186940 184900 186992
rect 247224 186940 247276 186992
rect 122748 186396 122800 186448
rect 174636 186396 174688 186448
rect 108948 186328 109000 186380
rect 193956 186328 194008 186380
rect 230388 185852 230440 185904
rect 231860 185852 231912 185904
rect 217968 185648 218020 185700
rect 229192 185648 229244 185700
rect 181536 185580 181588 185632
rect 240232 185580 240284 185632
rect 240784 185580 240836 185632
rect 296996 185580 297048 185632
rect 124128 184968 124180 185020
rect 164884 184968 164936 185020
rect 106188 184900 106240 184952
rect 182916 184900 182968 184952
rect 207664 184220 207716 184272
rect 238760 184220 238812 184272
rect 276664 184220 276716 184272
rect 292856 184220 292908 184272
rect 180156 184152 180208 184204
rect 192484 184152 192536 184204
rect 217324 184152 217376 184204
rect 284484 184152 284536 184204
rect 103428 183608 103480 183660
rect 169024 183608 169076 183660
rect 128268 183540 128320 183592
rect 214656 183540 214708 183592
rect 215208 182860 215260 182912
rect 234712 182860 234764 182912
rect 282276 182860 282328 182912
rect 294236 182860 294288 182912
rect 179328 182792 179380 182844
rect 226340 182792 226392 182844
rect 242256 182792 242308 182844
rect 253940 182792 253992 182844
rect 265624 182792 265676 182844
rect 281632 182792 281684 182844
rect 282184 182792 282236 182844
rect 309416 182792 309468 182844
rect 133144 182248 133196 182300
rect 164516 182248 164568 182300
rect 148232 182180 148284 182232
rect 214564 182180 214616 182232
rect 229744 182112 229796 182164
rect 230756 182112 230808 182164
rect 233976 181568 234028 181620
rect 245752 181568 245804 181620
rect 220084 181500 220136 181552
rect 234896 181500 234948 181552
rect 273904 181500 273956 181552
rect 295524 181500 295576 181552
rect 211804 181432 211856 181484
rect 226892 181432 226944 181484
rect 235448 181432 235500 181484
rect 248604 181432 248656 181484
rect 251824 181432 251876 181484
rect 298284 181432 298336 181484
rect 125968 180888 126020 180940
rect 170496 180888 170548 180940
rect 132408 180820 132460 180872
rect 203616 180820 203668 180872
rect 222936 180208 222988 180260
rect 240324 180208 240376 180260
rect 279424 180208 279476 180260
rect 290096 180208 290148 180260
rect 186228 180140 186280 180192
rect 223396 180140 223448 180192
rect 269856 180140 269908 180192
rect 291476 180140 291528 180192
rect 169576 180072 169628 180124
rect 226340 180072 226392 180124
rect 238116 180072 238168 180124
rect 278780 180072 278832 180124
rect 229284 179936 229336 179988
rect 237472 179936 237524 179988
rect 121000 179460 121052 179512
rect 167828 179460 167880 179512
rect 112260 179392 112312 179444
rect 171784 179392 171836 179444
rect 246304 179392 246356 179444
rect 247132 179392 247184 179444
rect 574744 179324 574796 179376
rect 580172 179324 580224 179376
rect 278780 179052 278832 179104
rect 280344 179052 280396 179104
rect 278228 178916 278280 178968
rect 278780 178916 278832 178968
rect 227076 178712 227128 178764
rect 234804 178712 234856 178764
rect 199936 178644 199988 178696
rect 245844 178644 245896 178696
rect 271236 178644 271288 178696
rect 285864 178644 285916 178696
rect 124496 178100 124548 178152
rect 187056 178100 187108 178152
rect 116952 178032 117004 178084
rect 196808 178032 196860 178084
rect 298744 178032 298796 178084
rect 299756 178032 299808 178084
rect 201132 177964 201184 178016
rect 227812 177964 227864 178016
rect 286324 177964 286376 178016
rect 287060 177964 287112 178016
rect 205548 177896 205600 177948
rect 223488 177896 223540 177948
rect 226892 177352 226944 177404
rect 238944 177352 238996 177404
rect 273996 177352 274048 177404
rect 284576 177352 284628 177404
rect 228456 177284 228508 177336
rect 233240 177284 233292 177336
rect 233884 177284 233936 177336
rect 251180 177284 251232 177336
rect 268476 177284 268528 177336
rect 283196 177284 283248 177336
rect 128176 176740 128228 176792
rect 166448 176740 166500 176792
rect 136088 176672 136140 176724
rect 158996 176672 159048 176724
rect 203524 176672 203576 176724
rect 213920 176604 213972 176656
rect 188804 176536 188856 176588
rect 228364 176536 228416 176588
rect 278136 176196 278188 176248
rect 285956 176196 286008 176248
rect 226340 175992 226392 176044
rect 233884 175992 233936 176044
rect 130752 175924 130804 175976
rect 165528 175924 165580 175976
rect 231768 175924 231820 175976
rect 245936 175924 245988 175976
rect 246396 175924 246448 175976
rect 253940 175924 253992 175976
rect 223672 175788 223724 175840
rect 163504 175176 163556 175228
rect 213920 175176 213972 175228
rect 243544 175312 243596 175364
rect 264980 175312 265032 175364
rect 253940 175244 253992 175296
rect 279332 175380 279384 175432
rect 164516 175108 164568 175160
rect 214012 175108 214064 175160
rect 231768 175176 231820 175228
rect 240140 175176 240192 175228
rect 230940 175108 230992 175160
rect 229744 174768 229796 174820
rect 232044 174768 232096 174820
rect 214104 174496 214156 174548
rect 229284 174496 229336 174548
rect 255964 173952 256016 174004
rect 264980 173952 265032 174004
rect 247776 173884 247828 173936
rect 265072 173884 265124 173936
rect 165528 173816 165580 173868
rect 214012 173816 214064 173868
rect 231584 173816 231636 173868
rect 247040 173816 247092 173868
rect 203616 173748 203668 173800
rect 213920 173748 213972 173800
rect 250536 172592 250588 172644
rect 264980 172592 265032 172644
rect 247684 172524 247736 172576
rect 265072 172524 265124 172576
rect 166264 172456 166316 172508
rect 213920 172456 213972 172508
rect 236368 172456 236420 172508
rect 238024 172456 238076 172508
rect 281540 172456 281592 172508
rect 291384 172456 291436 172508
rect 167644 172388 167696 172440
rect 215300 172388 215352 172440
rect 231124 172184 231176 172236
rect 233332 172184 233384 172236
rect 231768 171844 231820 171896
rect 237380 171844 237432 171896
rect 240876 171164 240928 171216
rect 264980 171164 265032 171216
rect 238116 171096 238168 171148
rect 265072 171096 265124 171148
rect 166448 171028 166500 171080
rect 214012 171028 214064 171080
rect 170496 170960 170548 171012
rect 213920 170960 213972 171012
rect 230664 170756 230716 170808
rect 232136 170756 232188 170808
rect 231216 170008 231268 170060
rect 233240 170008 233292 170060
rect 249248 169804 249300 169856
rect 264980 169804 265032 169856
rect 232136 169736 232188 169788
rect 236184 169736 236236 169788
rect 240968 169736 241020 169788
rect 265072 169736 265124 169788
rect 169300 169668 169352 169720
rect 214012 169668 214064 169720
rect 187056 169600 187108 169652
rect 213920 169600 213972 169652
rect 281540 169600 281592 169652
rect 287060 169600 287112 169652
rect 231676 169396 231728 169448
rect 234896 169396 234948 169448
rect 238392 168512 238444 168564
rect 238852 168512 238904 168564
rect 233976 168376 234028 168428
rect 264980 168376 265032 168428
rect 167828 168308 167880 168360
rect 214012 168308 214064 168360
rect 174636 168240 174688 168292
rect 213920 168240 213972 168292
rect 230940 168240 230992 168292
rect 233424 168240 233476 168292
rect 231676 167424 231728 167476
rect 236276 167424 236328 167476
rect 242164 167084 242216 167136
rect 264980 167084 265032 167136
rect 235264 167016 235316 167068
rect 265072 167016 265124 167068
rect 169116 166948 169168 167000
rect 213920 166948 213972 167000
rect 231308 166948 231360 167000
rect 234804 166948 234856 167000
rect 196808 166880 196860 166932
rect 214012 166880 214064 166932
rect 282828 166404 282880 166456
rect 288716 166404 288768 166456
rect 230572 166268 230624 166320
rect 230940 166268 230992 166320
rect 231676 166268 231728 166320
rect 232136 166268 232188 166320
rect 239680 165656 239732 165708
rect 264980 165656 265032 165708
rect 232780 165588 232832 165640
rect 265072 165588 265124 165640
rect 166356 165520 166408 165572
rect 214012 165520 214064 165572
rect 231124 165520 231176 165572
rect 234712 165520 234764 165572
rect 282828 165520 282880 165572
rect 302424 165520 302476 165572
rect 191288 165452 191340 165504
rect 213920 165452 213972 165504
rect 236920 164840 236972 164892
rect 265164 164840 265216 164892
rect 236644 164228 236696 164280
rect 264980 164228 265032 164280
rect 3240 164160 3292 164212
rect 15844 164160 15896 164212
rect 171784 164160 171836 164212
rect 214012 164160 214064 164212
rect 231584 164160 231636 164212
rect 249892 164160 249944 164212
rect 282828 164160 282880 164212
rect 299756 164160 299808 164212
rect 177488 164092 177540 164144
rect 213920 164092 213972 164144
rect 231492 163956 231544 164008
rect 236000 163956 236052 164008
rect 282828 163140 282880 163192
rect 288624 163140 288676 163192
rect 250628 162936 250680 162988
rect 264980 162936 265032 162988
rect 245200 162868 245252 162920
rect 265072 162868 265124 162920
rect 171968 162800 172020 162852
rect 213920 162800 213972 162852
rect 231768 162800 231820 162852
rect 247224 162800 247276 162852
rect 282736 162800 282788 162852
rect 306564 162800 306616 162852
rect 185676 162732 185728 162784
rect 214012 162732 214064 162784
rect 282828 162732 282880 162784
rect 301136 162732 301188 162784
rect 232596 162120 232648 162172
rect 241704 162120 241756 162172
rect 257344 161508 257396 161560
rect 264980 161508 265032 161560
rect 246488 161440 246540 161492
rect 265072 161440 265124 161492
rect 169208 161372 169260 161424
rect 214012 161372 214064 161424
rect 231768 161372 231820 161424
rect 240232 161372 240284 161424
rect 282736 161372 282788 161424
rect 299572 161372 299624 161424
rect 193956 161304 194008 161356
rect 213920 161304 213972 161356
rect 282828 161304 282880 161356
rect 296996 161304 297048 161356
rect 231308 160964 231360 161016
rect 233516 160964 233568 161016
rect 246396 160148 246448 160200
rect 264980 160148 265032 160200
rect 240784 160080 240836 160132
rect 265072 160080 265124 160132
rect 182916 160012 182968 160064
rect 213920 160012 213972 160064
rect 231768 160012 231820 160064
rect 251272 160012 251324 160064
rect 282460 160012 282512 160064
rect 302516 160012 302568 160064
rect 195520 159944 195572 159996
rect 214012 159944 214064 159996
rect 231676 159944 231728 159996
rect 244556 159944 244608 159996
rect 282552 159740 282604 159792
rect 285956 159740 286008 159792
rect 171876 159332 171928 159384
rect 188344 159332 188396 159384
rect 244924 159332 244976 159384
rect 265164 159332 265216 159384
rect 167736 158992 167788 159044
rect 169208 158992 169260 159044
rect 260196 158720 260248 158772
rect 264980 158720 265032 158772
rect 169024 158652 169076 158704
rect 213920 158652 213972 158704
rect 282092 158652 282144 158704
rect 292856 158652 292908 158704
rect 181536 158584 181588 158636
rect 214012 158584 214064 158636
rect 231492 158108 231544 158160
rect 233884 158108 233936 158160
rect 233884 157972 233936 158024
rect 242256 157972 242308 158024
rect 253296 157972 253348 158024
rect 265072 157972 265124 158024
rect 282276 157972 282328 158024
rect 298376 157972 298428 158024
rect 251916 157360 251968 157412
rect 264980 157360 265032 157412
rect 166540 157292 166592 157344
rect 213920 157292 213972 157344
rect 231768 157292 231820 157344
rect 242992 157292 243044 157344
rect 180340 157224 180392 157276
rect 214012 157224 214064 157276
rect 231492 156612 231544 156664
rect 240324 156612 240376 156664
rect 250444 156000 250496 156052
rect 264980 156000 265032 156052
rect 241060 155932 241112 155984
rect 265072 155932 265124 155984
rect 178868 155864 178920 155916
rect 213920 155864 213972 155916
rect 282184 155864 282236 155916
rect 309232 155864 309284 155916
rect 230756 155796 230808 155848
rect 232504 155796 232556 155848
rect 282828 155796 282880 155848
rect 303804 155796 303856 155848
rect 231768 155388 231820 155440
rect 237472 155388 237524 155440
rect 239496 154640 239548 154692
rect 264980 154640 265032 154692
rect 238208 154572 238260 154624
rect 265164 154572 265216 154624
rect 231584 154504 231636 154556
rect 245844 154504 245896 154556
rect 282368 154504 282420 154556
rect 295616 154504 295668 154556
rect 282092 154436 282144 154488
rect 294236 154436 294288 154488
rect 231676 154300 231728 154352
rect 234068 154300 234120 154352
rect 234160 153824 234212 153876
rect 265624 153824 265676 153876
rect 264520 153416 264572 153468
rect 265808 153416 265860 153468
rect 203616 153212 203668 153264
rect 213920 153212 213972 153264
rect 211896 152056 211948 152108
rect 214012 152056 214064 152108
rect 238392 151852 238444 151904
rect 247868 151852 247920 151904
rect 264980 151852 265032 151904
rect 166264 151784 166316 151836
rect 213920 151784 213972 151836
rect 230756 151784 230808 151836
rect 238024 151784 238076 151836
rect 265072 151784 265124 151836
rect 231768 151716 231820 151768
rect 244464 151716 244516 151768
rect 282828 151716 282880 151768
rect 305184 151716 305236 151768
rect 184296 150492 184348 150544
rect 214012 150492 214064 150544
rect 264520 150492 264572 150544
rect 266268 150492 266320 150544
rect 169116 150424 169168 150476
rect 213920 150424 213972 150476
rect 242440 150424 242492 150476
rect 264980 150424 265032 150476
rect 169208 150356 169260 150408
rect 214012 150356 214064 150408
rect 231768 150356 231820 150408
rect 247132 150356 247184 150408
rect 2780 150288 2832 150340
rect 4804 150288 4856 150340
rect 231492 150288 231544 150340
rect 244280 150288 244332 150340
rect 203524 149676 203576 149728
rect 213920 149676 213972 149728
rect 252008 149676 252060 149728
rect 265072 149676 265124 149728
rect 245108 149064 245160 149116
rect 264980 149064 265032 149116
rect 231768 148996 231820 149048
rect 255320 148996 255372 149048
rect 282828 148928 282880 148980
rect 290096 148928 290148 148980
rect 281540 148860 281592 148912
rect 283196 148860 283248 148912
rect 231308 148316 231360 148368
rect 248420 148316 248472 148368
rect 263140 147704 263192 147756
rect 265716 147704 265768 147756
rect 166356 147636 166408 147688
rect 213920 147636 213972 147688
rect 253480 147636 253532 147688
rect 264980 147636 265032 147688
rect 282828 147568 282880 147620
rect 307944 147568 307996 147620
rect 231124 146956 231176 147008
rect 240968 146956 241020 147008
rect 232872 146888 232924 146940
rect 254676 146888 254728 146940
rect 256240 146888 256292 146940
rect 265164 146888 265216 146940
rect 259000 146820 259052 146872
rect 265256 146820 265308 146872
rect 249432 146616 249484 146668
rect 257344 146616 257396 146668
rect 185676 146276 185728 146328
rect 213920 146276 213972 146328
rect 230756 146140 230808 146192
rect 232596 146140 232648 146192
rect 170404 145528 170456 145580
rect 209044 145528 209096 145580
rect 234068 144984 234120 145036
rect 265072 144984 265124 145036
rect 203524 144916 203576 144968
rect 213920 144916 213972 144968
rect 232504 144916 232556 144968
rect 264980 144916 265032 144968
rect 282460 144848 282512 144900
rect 310612 144848 310664 144900
rect 281908 144780 281960 144832
rect 298284 144780 298336 144832
rect 230296 144168 230348 144220
rect 242900 144168 242952 144220
rect 243820 144168 243872 144220
rect 265164 144168 265216 144220
rect 204904 143624 204956 143676
rect 213920 143624 213972 143676
rect 177488 143556 177540 143608
rect 214012 143556 214064 143608
rect 240968 143556 241020 143608
rect 264980 143556 265032 143608
rect 231768 143488 231820 143540
rect 250076 143488 250128 143540
rect 282092 143488 282144 143540
rect 295340 143488 295392 143540
rect 185584 142808 185636 142860
rect 200764 142808 200816 142860
rect 230664 142808 230716 142860
rect 251180 142808 251232 142860
rect 260288 142196 260340 142248
rect 265072 142196 265124 142248
rect 207756 142128 207808 142180
rect 213920 142128 213972 142180
rect 254676 142128 254728 142180
rect 264980 142128 265032 142180
rect 281908 142060 281960 142112
rect 284576 142060 284628 142112
rect 186964 141448 187016 141500
rect 195244 141448 195296 141500
rect 231216 141448 231268 141500
rect 254584 141448 254636 141500
rect 192576 141380 192628 141432
rect 214012 141380 214064 141432
rect 230940 141380 230992 141432
rect 255964 141380 256016 141432
rect 282276 141312 282328 141364
rect 285864 141312 285916 141364
rect 261668 140836 261720 140888
rect 265164 140836 265216 140888
rect 256056 140768 256108 140820
rect 264980 140768 265032 140820
rect 231308 140700 231360 140752
rect 236092 140700 236144 140752
rect 282276 140700 282328 140752
rect 311992 140700 312044 140752
rect 281724 140632 281776 140684
rect 300952 140632 301004 140684
rect 234344 140020 234396 140072
rect 260196 140020 260248 140072
rect 210424 139476 210476 139528
rect 214012 139476 214064 139528
rect 260380 139476 260432 139528
rect 265900 139476 265952 139528
rect 206284 139408 206336 139460
rect 213920 139408 213972 139460
rect 256148 139408 256200 139460
rect 264980 139408 265032 139460
rect 231768 139340 231820 139392
rect 255412 139340 255464 139392
rect 282276 139340 282328 139392
rect 302240 139340 302292 139392
rect 282828 139272 282880 139324
rect 296904 139272 296956 139324
rect 173164 138660 173216 138712
rect 214472 138660 214524 138712
rect 250720 138660 250772 138712
rect 265624 138660 265676 138712
rect 211804 137980 211856 138032
rect 213920 137980 213972 138032
rect 257620 137980 257672 138032
rect 264980 137980 265032 138032
rect 3516 137912 3568 137964
rect 32404 137912 32456 137964
rect 231584 137912 231636 137964
rect 252652 137912 252704 137964
rect 281724 137912 281776 137964
rect 291476 137912 291528 137964
rect 231676 137572 231728 137624
rect 238300 137572 238352 137624
rect 167736 137232 167788 137284
rect 215944 137232 215996 137284
rect 178868 136620 178920 136672
rect 213920 136620 213972 136672
rect 254584 136620 254636 136672
rect 264980 136620 265032 136672
rect 231400 136552 231452 136604
rect 247776 136552 247828 136604
rect 281908 136484 281960 136536
rect 301044 136484 301096 136536
rect 231308 135940 231360 135992
rect 239680 135940 239732 135992
rect 177396 135872 177448 135924
rect 198188 135872 198240 135924
rect 239588 135872 239640 135924
rect 265256 135872 265308 135924
rect 207664 135328 207716 135380
rect 214012 135328 214064 135380
rect 202788 135260 202840 135312
rect 213920 135260 213972 135312
rect 258724 135260 258776 135312
rect 265072 135260 265124 135312
rect 231768 135192 231820 135244
rect 260104 135192 260156 135244
rect 282092 135192 282144 135244
rect 289820 135192 289872 135244
rect 231492 135124 231544 135176
rect 247684 135124 247736 135176
rect 169024 134580 169076 134632
rect 202788 134580 202840 134632
rect 177396 134512 177448 134564
rect 211896 134512 211948 134564
rect 209320 133900 209372 133952
rect 213920 133900 213972 133952
rect 257344 133900 257396 133952
rect 264980 133900 265032 133952
rect 282276 133832 282328 133884
rect 294144 133832 294196 133884
rect 282828 133764 282880 133816
rect 292672 133764 292724 133816
rect 230572 133560 230624 133612
rect 233976 133560 234028 133612
rect 231676 133220 231728 133272
rect 238116 133220 238168 133272
rect 247684 132540 247736 132592
rect 264980 132540 265032 132592
rect 206468 132472 206520 132524
rect 213920 132472 213972 132524
rect 233884 132472 233936 132524
rect 265072 132472 265124 132524
rect 231768 132404 231820 132456
rect 257436 132404 257488 132456
rect 282736 132404 282788 132456
rect 306656 132404 306708 132456
rect 282828 132336 282880 132388
rect 299664 132336 299716 132388
rect 181536 131724 181588 131776
rect 214656 131724 214708 131776
rect 232596 131180 232648 131232
rect 191288 131112 191340 131164
rect 213920 131112 213972 131164
rect 230940 131112 230992 131164
rect 232780 131112 232832 131164
rect 261576 131180 261628 131232
rect 265072 131180 265124 131232
rect 264980 131112 265032 131164
rect 231768 131044 231820 131096
rect 249248 131044 249300 131096
rect 282276 131044 282328 131096
rect 313372 131044 313424 131096
rect 281540 130568 281592 130620
rect 284484 130568 284536 130620
rect 202328 129820 202380 129872
rect 214012 129820 214064 129872
rect 171784 129752 171836 129804
rect 213920 129752 213972 129804
rect 235356 129752 235408 129804
rect 264980 129752 265032 129804
rect 231768 129684 231820 129736
rect 264244 129684 264296 129736
rect 282092 129684 282144 129736
rect 309416 129684 309468 129736
rect 230756 129548 230808 129600
rect 236920 129548 236972 129600
rect 209228 128392 209280 128444
rect 214012 128392 214064 128444
rect 178776 128324 178828 128376
rect 213920 128324 213972 128376
rect 237012 128324 237064 128376
rect 264980 128324 265032 128376
rect 231768 128256 231820 128308
rect 242164 128256 242216 128308
rect 282828 128256 282880 128308
rect 313280 128256 313332 128308
rect 282736 128188 282788 128240
rect 287244 128188 287296 128240
rect 231124 127712 231176 127764
rect 235264 127712 235316 127764
rect 250812 127576 250864 127628
rect 258724 127576 258776 127628
rect 185768 127032 185820 127084
rect 213920 127032 213972 127084
rect 173256 126964 173308 127016
rect 214012 126964 214064 127016
rect 246304 126964 246356 127016
rect 264980 126964 265032 127016
rect 231768 126896 231820 126948
rect 239404 126896 239456 126948
rect 282276 126896 282328 126948
rect 288532 126896 288584 126948
rect 249340 126284 249392 126336
rect 265900 126284 265952 126336
rect 231400 126216 231452 126268
rect 249432 126216 249484 126268
rect 196808 125672 196860 125724
rect 214012 125672 214064 125724
rect 169208 125604 169260 125656
rect 213920 125604 213972 125656
rect 258724 125604 258776 125656
rect 264980 125604 265032 125656
rect 230480 125536 230532 125588
rect 234160 125536 234212 125588
rect 282828 125536 282880 125588
rect 314660 125536 314712 125588
rect 282092 125468 282144 125520
rect 298192 125468 298244 125520
rect 186964 124856 187016 124908
rect 206284 124856 206336 124908
rect 230664 124856 230716 124908
rect 240784 124856 240836 124908
rect 176016 124176 176068 124228
rect 213920 124176 213972 124228
rect 235264 124176 235316 124228
rect 264980 124176 265032 124228
rect 231768 124108 231820 124160
rect 261760 124108 261812 124160
rect 282276 124108 282328 124160
rect 307760 124108 307812 124160
rect 231400 124040 231452 124092
rect 250628 124040 250680 124092
rect 282828 124040 282880 124092
rect 294052 124040 294104 124092
rect 210608 123088 210660 123140
rect 214012 123088 214064 123140
rect 262128 123020 262180 123072
rect 265072 123020 265124 123072
rect 174636 122816 174688 122868
rect 213920 122816 213972 122868
rect 257528 122816 257580 122868
rect 264980 122816 265032 122868
rect 231768 122748 231820 122800
rect 263048 122748 263100 122800
rect 282460 122748 282512 122800
rect 303620 122748 303672 122800
rect 231492 122680 231544 122732
rect 244924 122680 244976 122732
rect 282644 122068 282696 122120
rect 295524 122068 295576 122120
rect 199476 121524 199528 121576
rect 214012 121524 214064 121576
rect 178960 121456 179012 121508
rect 213920 121456 213972 121508
rect 252100 121456 252152 121508
rect 264980 121456 265032 121508
rect 231768 121388 231820 121440
rect 246488 121388 246540 121440
rect 282828 121388 282880 121440
rect 305276 121388 305328 121440
rect 169300 120708 169352 120760
rect 214840 120708 214892 120760
rect 191380 120096 191432 120148
rect 213920 120096 213972 120148
rect 231400 120096 231452 120148
rect 238024 120096 238076 120148
rect 240784 120096 240836 120148
rect 264980 120096 265032 120148
rect 231492 120028 231544 120080
rect 253296 120028 253348 120080
rect 282092 120028 282144 120080
rect 285772 120028 285824 120080
rect 282184 119348 282236 119400
rect 307852 119348 307904 119400
rect 206284 118736 206336 118788
rect 213920 118736 213972 118788
rect 181628 118668 181680 118720
rect 214012 118668 214064 118720
rect 230940 118668 230992 118720
rect 234344 118668 234396 118720
rect 231584 118600 231636 118652
rect 251916 118600 251968 118652
rect 281816 118396 281868 118448
rect 284392 118396 284444 118448
rect 264336 117988 264388 118040
rect 264612 117988 264664 118040
rect 230756 117920 230808 117972
rect 241060 117920 241112 117972
rect 207848 117376 207900 117428
rect 213920 117376 213972 117428
rect 253204 117376 253256 117428
rect 265072 117376 265124 117428
rect 170588 117308 170640 117360
rect 214012 117308 214064 117360
rect 242164 117308 242216 117360
rect 264980 117308 265032 117360
rect 231768 117240 231820 117292
rect 242256 117240 242308 117292
rect 282828 117240 282880 117292
rect 292764 117240 292816 117292
rect 231492 117172 231544 117224
rect 236828 117172 236880 117224
rect 282368 117104 282420 117156
rect 287152 117104 287204 117156
rect 206376 116016 206428 116068
rect 214012 116016 214064 116068
rect 263232 116016 263284 116068
rect 265072 116016 265124 116068
rect 189816 115948 189868 116000
rect 213920 115948 213972 116000
rect 253296 115948 253348 116000
rect 264980 115948 265032 116000
rect 203708 115880 203760 115932
rect 204996 115880 205048 115932
rect 231492 115880 231544 115932
rect 263140 115880 263192 115932
rect 282828 115880 282880 115932
rect 302332 115880 302384 115932
rect 230940 115812 230992 115864
rect 238208 115812 238260 115864
rect 282276 115336 282328 115388
rect 285680 115336 285732 115388
rect 195336 115200 195388 115252
rect 214932 115200 214984 115252
rect 205088 114520 205140 114572
rect 213920 114520 213972 114572
rect 242348 114520 242400 114572
rect 264980 114520 265032 114572
rect 231676 114452 231728 114504
rect 239496 114452 239548 114504
rect 230572 114112 230624 114164
rect 232688 114112 232740 114164
rect 188436 113228 188488 113280
rect 214012 113228 214064 113280
rect 249248 113228 249300 113280
rect 265072 113228 265124 113280
rect 176200 113160 176252 113212
rect 213920 113160 213972 113212
rect 234160 113160 234212 113212
rect 264980 113160 265032 113212
rect 231768 113092 231820 113144
rect 264520 113092 264572 113144
rect 282828 113092 282880 113144
rect 303712 113092 303764 113144
rect 231308 113024 231360 113076
rect 259000 113024 259052 113076
rect 282000 113024 282052 113076
rect 291200 113024 291252 113076
rect 184388 112412 184440 112464
rect 214840 112412 214892 112464
rect 187056 111800 187108 111852
rect 213920 111800 213972 111852
rect 260472 111800 260524 111852
rect 264980 111800 265032 111852
rect 168288 111732 168340 111784
rect 169116 111732 169168 111784
rect 231768 111732 231820 111784
rect 247868 111732 247920 111784
rect 282828 111732 282880 111784
rect 290004 111732 290056 111784
rect 231676 111664 231728 111716
rect 235448 111664 235500 111716
rect 209136 110508 209188 110560
rect 213920 110508 213972 110560
rect 255964 110508 256016 110560
rect 264980 110508 265032 110560
rect 170496 110440 170548 110492
rect 214012 110440 214064 110492
rect 244924 110440 244976 110492
rect 265072 110440 265124 110492
rect 167828 110372 167880 110424
rect 184296 110372 184348 110424
rect 231768 110372 231820 110424
rect 252008 110372 252060 110424
rect 282276 110372 282328 110424
rect 296812 110372 296864 110424
rect 231216 110304 231268 110356
rect 242440 110304 242492 110356
rect 282828 109760 282880 109812
rect 287336 109760 287388 109812
rect 200856 109080 200908 109132
rect 202328 109080 202380 109132
rect 173348 109012 173400 109064
rect 213920 109012 213972 109064
rect 257436 109012 257488 109064
rect 264980 109012 265032 109064
rect 231400 108944 231452 108996
rect 256240 108944 256292 108996
rect 231768 108876 231820 108928
rect 245108 108876 245160 108928
rect 281724 108876 281776 108928
rect 284300 108876 284352 108928
rect 282276 108264 282328 108316
rect 296720 108264 296772 108316
rect 210516 107720 210568 107772
rect 214012 107720 214064 107772
rect 259000 107720 259052 107772
rect 264980 107720 265032 107772
rect 202328 107652 202380 107704
rect 213920 107652 213972 107704
rect 250536 107652 250588 107704
rect 265072 107652 265124 107704
rect 231216 107584 231268 107636
rect 253480 107584 253532 107636
rect 231768 107516 231820 107568
rect 250720 107516 250772 107568
rect 184480 106360 184532 106412
rect 213920 106360 213972 106412
rect 253388 106360 253440 106412
rect 264980 106360 265032 106412
rect 167828 106292 167880 106344
rect 214012 106292 214064 106344
rect 251916 106292 251968 106344
rect 265072 106292 265124 106344
rect 231768 106224 231820 106276
rect 260380 106224 260432 106276
rect 282828 106224 282880 106276
rect 291292 106224 291344 106276
rect 166540 105544 166592 105596
rect 204904 105544 204956 105596
rect 230756 105544 230808 105596
rect 253940 105544 253992 105596
rect 204996 104932 205048 104984
rect 213920 104932 213972 104984
rect 258816 104932 258868 104984
rect 265072 104932 265124 104984
rect 174728 104864 174780 104916
rect 214012 104864 214064 104916
rect 260196 104864 260248 104916
rect 264980 104864 265032 104916
rect 231308 104796 231360 104848
rect 243820 104796 243872 104848
rect 254860 104796 254912 104848
rect 257620 104796 257672 104848
rect 282828 104796 282880 104848
rect 310520 104796 310572 104848
rect 282000 104728 282052 104780
rect 292580 104728 292632 104780
rect 231308 103912 231360 103964
rect 234068 103912 234120 103964
rect 191196 103504 191248 103556
rect 213920 103504 213972 103556
rect 233976 103504 234028 103556
rect 264980 103504 265032 103556
rect 282828 103436 282880 103488
rect 289912 103436 289964 103488
rect 231584 103368 231636 103420
rect 240968 103368 241020 103420
rect 282736 103096 282788 103148
rect 288440 103096 288492 103148
rect 230572 102824 230624 102876
rect 232504 102824 232556 102876
rect 173440 102756 173492 102808
rect 191380 102756 191432 102808
rect 192668 102212 192720 102264
rect 213920 102212 213972 102264
rect 171968 102144 172020 102196
rect 214012 102144 214064 102196
rect 250628 102144 250680 102196
rect 264980 102144 265032 102196
rect 231676 102076 231728 102128
rect 254676 102076 254728 102128
rect 282828 102076 282880 102128
rect 309324 102076 309376 102128
rect 231400 102008 231452 102060
rect 239588 102008 239640 102060
rect 260380 100784 260432 100836
rect 265072 100784 265124 100836
rect 177580 100716 177632 100768
rect 213920 100716 213972 100768
rect 246396 100716 246448 100768
rect 264980 100716 265032 100768
rect 231768 100648 231820 100700
rect 261668 100648 261720 100700
rect 281724 100648 281776 100700
rect 295432 100648 295484 100700
rect 231676 100580 231728 100632
rect 245016 100580 245068 100632
rect 167736 99968 167788 100020
rect 211804 99968 211856 100020
rect 211896 99424 211948 99476
rect 214012 99424 214064 99476
rect 169116 99356 169168 99408
rect 213920 99356 213972 99408
rect 245200 99356 245252 99408
rect 264980 99356 265032 99408
rect 231400 99288 231452 99340
rect 246580 99288 246632 99340
rect 231216 99220 231268 99272
rect 243544 99220 243596 99272
rect 253480 98336 253532 98388
rect 256148 98336 256200 98388
rect 211804 98064 211856 98116
rect 214012 98064 214064 98116
rect 167920 97996 167972 98048
rect 213920 97996 213972 98048
rect 256240 97996 256292 98048
rect 264980 97996 265032 98048
rect 3424 97928 3476 97980
rect 17224 97928 17276 97980
rect 169576 97928 169628 97980
rect 232780 97928 232832 97980
rect 231216 97860 231268 97912
rect 256056 97860 256108 97912
rect 184664 97248 184716 97300
rect 213276 97248 213328 97300
rect 263140 96704 263192 96756
rect 265072 96704 265124 96756
rect 229008 96636 229060 96688
rect 256148 96636 256200 96688
rect 264980 96636 265032 96688
rect 223672 96024 223724 96076
rect 164976 95956 165028 96008
rect 185676 95956 185728 96008
rect 165896 95888 165948 95940
rect 210608 95888 210660 95940
rect 244280 95616 244332 95668
rect 249800 95616 249852 95668
rect 230480 95480 230532 95532
rect 232504 95480 232556 95532
rect 225604 95276 225656 95328
rect 187976 95208 188028 95260
rect 213920 95208 213972 95260
rect 227076 95208 227128 95260
rect 229100 95208 229152 95260
rect 262680 95208 262732 95260
rect 213368 95140 213420 95192
rect 281540 95140 281592 95192
rect 67456 94528 67508 94580
rect 108304 94528 108356 94580
rect 64696 94460 64748 94512
rect 111064 94460 111116 94512
rect 222936 94460 222988 94512
rect 234252 94460 234304 94512
rect 125416 93916 125468 93968
rect 169208 93916 169260 93968
rect 110144 93848 110196 93900
rect 207848 93848 207900 93900
rect 249800 93780 249852 93832
rect 273996 93780 274048 93832
rect 261484 93712 261536 93764
rect 281724 93712 281776 93764
rect 162768 93168 162820 93220
rect 177396 93168 177448 93220
rect 179052 93168 179104 93220
rect 214564 93168 214616 93220
rect 108120 93100 108172 93152
rect 121460 93100 121512 93152
rect 121736 93100 121788 93152
rect 174636 93100 174688 93152
rect 209136 93100 209188 93152
rect 259000 93100 259052 93152
rect 105728 92488 105780 92540
rect 112444 92488 112496 92540
rect 222844 92488 222896 92540
rect 230020 92488 230072 92540
rect 136088 92420 136140 92472
rect 166356 92420 166408 92472
rect 152096 92352 152148 92404
rect 162768 92352 162820 92404
rect 166448 91808 166500 91860
rect 178868 91808 178920 91860
rect 208400 91808 208452 91860
rect 253480 91808 253532 91860
rect 67364 91740 67416 91792
rect 106924 91740 106976 91792
rect 164884 91740 164936 91792
rect 207664 91740 207716 91792
rect 214564 91740 214616 91792
rect 265808 91740 265860 91792
rect 115480 91128 115532 91180
rect 133144 91128 133196 91180
rect 100024 91060 100076 91112
rect 104256 91060 104308 91112
rect 118056 91060 118108 91112
rect 135904 91060 135956 91112
rect 113456 90992 113508 91044
rect 206284 90992 206336 91044
rect 111616 90924 111668 90976
rect 170588 90924 170640 90976
rect 176108 90380 176160 90432
rect 209320 90380 209372 90432
rect 218704 90380 218756 90432
rect 239680 90380 239732 90432
rect 66168 90312 66220 90364
rect 104164 90312 104216 90364
rect 207664 90312 207716 90364
rect 267280 90312 267332 90364
rect 115572 89632 115624 89684
rect 181628 89632 181680 89684
rect 121184 89564 121236 89616
rect 165896 89564 165948 89616
rect 221464 89020 221516 89072
rect 245108 89020 245160 89072
rect 67548 88952 67600 89004
rect 115204 88952 115256 89004
rect 213276 88952 213328 89004
rect 260472 88952 260524 89004
rect 203524 88340 203576 88392
rect 208400 88340 208452 88392
rect 119712 88272 119764 88324
rect 199476 88272 199528 88324
rect 206284 87660 206336 87712
rect 229836 87660 229888 87712
rect 165068 87592 165120 87644
rect 203616 87592 203668 87644
rect 214748 87592 214800 87644
rect 247960 87592 248012 87644
rect 93216 86912 93268 86964
rect 167828 86912 167880 86964
rect 151544 86844 151596 86896
rect 166264 86844 166316 86896
rect 220084 86300 220136 86352
rect 254860 86300 254912 86352
rect 184296 86232 184348 86284
rect 235540 86232 235592 86284
rect 3148 85484 3200 85536
rect 11704 85484 11756 85536
rect 105544 85484 105596 85536
rect 205088 85484 205140 85536
rect 126520 85416 126572 85468
rect 196808 85416 196860 85468
rect 215944 84872 215996 84924
rect 231308 84872 231360 84924
rect 226984 84804 227036 84856
rect 245200 84804 245252 84856
rect 96528 84124 96580 84176
rect 182916 84124 182968 84176
rect 97816 84056 97868 84108
rect 173348 84056 173400 84108
rect 195244 83512 195296 83564
rect 232872 83512 232924 83564
rect 178684 83444 178736 83496
rect 281540 83444 281592 83496
rect 100576 82764 100628 82816
rect 187056 82764 187108 82816
rect 107568 82696 107620 82748
rect 184388 82696 184440 82748
rect 95148 81336 95200 81388
rect 202328 81336 202380 81388
rect 129648 81268 129700 81320
rect 177488 81268 177540 81320
rect 133788 79976 133840 80028
rect 216036 79976 216088 80028
rect 117228 79908 117280 79960
rect 173440 79908 173492 79960
rect 118516 78616 118568 78668
rect 169208 78616 169260 78668
rect 151636 78548 151688 78600
rect 165068 78548 165120 78600
rect 174544 77936 174596 77988
rect 241520 77936 241572 77988
rect 91008 77188 91060 77240
rect 174728 77188 174780 77240
rect 126244 76508 126296 76560
rect 265716 76508 265768 76560
rect 104256 75828 104308 75880
rect 170496 75828 170548 75880
rect 119988 75148 120040 75200
rect 254768 75148 254820 75200
rect 124864 74468 124916 74520
rect 206468 74468 206520 74520
rect 114284 74400 114336 74452
rect 164884 74400 164936 74452
rect 117136 73108 117188 73160
rect 162124 73108 162176 73160
rect 151728 73040 151780 73092
rect 181536 73040 181588 73092
rect 3424 71680 3476 71732
rect 39304 71680 39356 71732
rect 64788 71680 64840 71732
rect 204996 71680 205048 71732
rect 119896 71612 119948 71664
rect 167736 71612 167788 71664
rect 102048 70320 102100 70372
rect 179052 70320 179104 70372
rect 131028 70252 131080 70304
rect 173164 70252 173216 70304
rect 122748 68960 122800 69012
rect 210424 68960 210476 69012
rect 130384 68280 130436 68332
rect 169760 68280 169812 68332
rect 110236 67532 110288 67584
rect 176108 67532 176160 67584
rect 133144 67464 133196 67516
rect 166448 67464 166500 67516
rect 104716 66172 104768 66224
rect 180156 66172 180208 66224
rect 124036 66104 124088 66156
rect 195336 66104 195388 66156
rect 103336 64812 103388 64864
rect 200856 64812 200908 64864
rect 122104 64744 122156 64796
rect 192668 64744 192720 64796
rect 228456 64132 228508 64184
rect 267740 64132 267792 64184
rect 111708 63452 111760 63504
rect 199384 63452 199436 63504
rect 93768 62772 93820 62824
rect 267096 62772 267148 62824
rect 121368 62024 121420 62076
rect 186964 62024 187016 62076
rect 77208 61344 77260 61396
rect 253388 61344 253440 61396
rect 107568 60052 107620 60104
rect 229744 60052 229796 60104
rect 79968 59984 80020 60036
rect 251916 59984 251968 60036
rect 3056 59304 3108 59356
rect 33784 59304 33836 59356
rect 112444 59304 112496 59356
rect 191288 59304 191340 59356
rect 86868 58624 86920 58676
rect 250444 58624 250496 58676
rect 99196 57876 99248 57928
rect 178776 57876 178828 57928
rect 100668 57196 100720 57248
rect 236736 57196 236788 57248
rect 115664 56516 115716 56568
rect 216128 56516 216180 56568
rect 91008 55836 91060 55888
rect 243728 55836 243780 55888
rect 110328 55156 110380 55208
rect 206376 55156 206428 55208
rect 97908 54476 97960 54528
rect 242256 54476 242308 54528
rect 85488 53728 85540 53780
rect 214656 53728 214708 53780
rect 102048 53048 102100 53100
rect 257436 53048 257488 53100
rect 86776 52368 86828 52420
rect 211804 52368 211856 52420
rect 124128 52300 124180 52352
rect 176016 52300 176068 52352
rect 95056 51008 95108 51060
rect 210516 51008 210568 51060
rect 111708 50328 111760 50380
rect 255964 50328 256016 50380
rect 70308 48968 70360 49020
rect 260196 48968 260248 49020
rect 115848 47608 115900 47660
rect 244924 47608 244976 47660
rect 31668 47540 31720 47592
rect 254584 47540 254636 47592
rect 98644 46248 98696 46300
rect 207664 46248 207716 46300
rect 22008 46180 22060 46232
rect 245016 46180 245068 46232
rect 3424 45500 3476 45552
rect 36544 45500 36596 45552
rect 66168 44888 66220 44940
rect 258816 44888 258868 44940
rect 50988 44820 51040 44872
rect 249800 44820 249852 44872
rect 124864 43460 124916 43512
rect 209228 43460 209280 43512
rect 217232 43460 217284 43512
rect 259460 43460 259512 43512
rect 34428 43392 34480 43444
rect 246396 43392 246448 43444
rect 122748 42100 122800 42152
rect 213276 42100 213328 42152
rect 45468 42032 45520 42084
rect 239496 42032 239548 42084
rect 85488 40740 85540 40792
rect 260104 40740 260156 40792
rect 46848 40672 46900 40724
rect 235356 40672 235408 40724
rect 99288 37952 99340 38004
rect 184296 37952 184348 38004
rect 49608 37884 49660 37936
rect 253296 37884 253348 37936
rect 200764 36592 200816 36644
rect 269120 36592 269172 36644
rect 56508 36524 56560 36576
rect 242164 36524 242216 36576
rect 4068 35232 4120 35284
rect 185584 35232 185636 35284
rect 53564 35164 53616 35216
rect 251824 35164 251876 35216
rect 61936 33804 61988 33856
rect 267188 33804 267240 33856
rect 53748 33736 53800 33788
rect 278780 33736 278832 33788
rect 3148 33056 3200 33108
rect 35164 33056 35216 33108
rect 124128 32444 124180 32496
rect 258724 32444 258776 32496
rect 44088 32376 44140 32428
rect 296720 32376 296772 32428
rect 54944 31084 54996 31136
rect 218704 31084 218756 31136
rect 37096 31016 37148 31068
rect 243636 31016 243688 31068
rect 59176 29656 59228 29708
rect 233976 29656 234028 29708
rect 62028 29588 62080 29640
rect 324412 29588 324464 29640
rect 84108 28296 84160 28348
rect 209136 28296 209188 28348
rect 1400 28228 1452 28280
rect 231216 28228 231268 28280
rect 90364 26868 90416 26920
rect 221464 26868 221516 26920
rect 113088 25508 113140 25560
rect 235264 25508 235316 25560
rect 111616 24080 111668 24132
rect 262864 24080 262916 24132
rect 123484 22788 123536 22840
rect 160744 22788 160796 22840
rect 39948 22720 40000 22772
rect 232688 22720 232740 22772
rect 188344 21428 188396 21480
rect 269120 21428 269172 21480
rect 92388 21360 92440 21412
rect 204904 21360 204956 21412
rect 3424 20612 3476 20664
rect 51724 20612 51776 20664
rect 48228 19932 48280 19984
rect 289820 19932 289872 19984
rect 103428 18640 103480 18692
rect 222936 18640 222988 18692
rect 55128 18572 55180 18624
rect 310520 18572 310572 18624
rect 209044 17280 209096 17332
rect 302240 17280 302292 17332
rect 81348 17212 81400 17264
rect 240784 17212 240836 17264
rect 181444 15920 181496 15972
rect 269764 15920 269816 15972
rect 110328 15852 110380 15904
rect 239404 15852 239456 15904
rect 135260 14696 135312 14748
rect 136456 14696 136508 14748
rect 121092 14492 121144 14544
rect 203524 14492 203576 14544
rect 12164 14424 12216 14476
rect 226984 14424 227036 14476
rect 118608 13132 118660 13184
rect 231124 13132 231176 13184
rect 60648 13064 60700 13116
rect 253204 13064 253256 13116
rect 198004 11772 198056 11824
rect 245200 11772 245252 11824
rect 96252 11704 96304 11756
rect 215944 11704 215996 11756
rect 259460 11704 259512 11756
rect 260656 11704 260708 11756
rect 307852 11704 307904 11756
rect 309048 11704 309100 11756
rect 332692 11704 332744 11756
rect 333888 11704 333940 11756
rect 114468 10344 114520 10396
rect 220084 10344 220136 10396
rect 9588 10276 9640 10328
rect 180064 10276 180116 10328
rect 184204 10276 184256 10328
rect 244096 10276 244148 10328
rect 77392 8984 77444 9036
rect 98644 8984 98696 9036
rect 177304 8984 177356 9036
rect 242900 8984 242952 9036
rect 97816 8916 97868 8968
rect 264244 8916 264296 8968
rect 224224 7556 224276 7608
rect 253480 7556 253532 7608
rect 71504 6196 71556 6248
rect 233884 6196 233936 6248
rect 47860 6128 47912 6180
rect 228364 6128 228416 6180
rect 238024 6128 238076 6180
rect 267740 6128 267792 6180
rect 340972 6128 341024 6180
rect 349160 6128 349212 6180
rect 304356 5516 304408 5568
rect 305092 5516 305144 5568
rect 95148 4836 95200 4888
rect 267004 4836 267056 4888
rect 20628 4768 20680 4820
rect 228456 4768 228508 4820
rect 318064 4768 318116 4820
rect 329196 4768 329248 4820
rect 232504 4156 232556 4208
rect 235816 4156 235868 4208
rect 296076 4088 296128 4140
rect 298100 4088 298152 4140
rect 304264 3952 304316 4004
rect 307944 3952 307996 4004
rect 11152 3544 11204 3596
rect 12256 3544 12308 3596
rect 35992 3544 36044 3596
rect 37096 3544 37148 3596
rect 44272 3544 44324 3596
rect 45376 3544 45428 3596
rect 64328 3544 64380 3596
rect 64788 3544 64840 3596
rect 69112 3544 69164 3596
rect 70216 3544 70268 3596
rect 119896 3544 119948 3596
rect 126244 3544 126296 3596
rect 2872 3476 2924 3528
rect 3976 3476 4028 3528
rect 8760 3476 8812 3528
rect 9588 3476 9640 3528
rect 9956 3476 10008 3528
rect 10968 3476 11020 3528
rect 17040 3476 17092 3528
rect 17868 3476 17920 3528
rect 18236 3476 18288 3528
rect 19248 3476 19300 3528
rect 19432 3476 19484 3528
rect 20536 3476 20588 3528
rect 24216 3476 24268 3528
rect 24768 3476 24820 3528
rect 25320 3476 25372 3528
rect 26148 3476 26200 3528
rect 27712 3476 27764 3528
rect 28816 3476 28868 3528
rect 32404 3476 32456 3528
rect 33048 3476 33100 3528
rect 33600 3476 33652 3528
rect 34428 3476 34480 3528
rect 34796 3476 34848 3528
rect 35808 3476 35860 3528
rect 40684 3476 40736 3528
rect 41236 3476 41288 3528
rect 43076 3476 43128 3528
rect 43996 3476 44048 3528
rect 48964 3476 49016 3528
rect 49608 3476 49660 3528
rect 50160 3476 50212 3528
rect 50896 3476 50948 3528
rect 52552 3476 52604 3528
rect 53564 3476 53616 3528
rect 56048 3476 56100 3528
rect 56508 3476 56560 3528
rect 57244 3476 57296 3528
rect 57888 3476 57940 3528
rect 58440 3476 58492 3528
rect 59176 3476 59228 3528
rect 59636 3476 59688 3528
rect 60648 3476 60700 3528
rect 63224 3476 63276 3528
rect 97816 3476 97868 3528
rect 98644 3476 98696 3528
rect 99288 3476 99340 3528
rect 99840 3476 99892 3528
rect 100668 3476 100720 3528
rect 101036 3476 101088 3528
rect 102048 3476 102100 3528
rect 105728 3476 105780 3528
rect 106188 3476 106240 3528
rect 106924 3476 106976 3528
rect 107568 3476 107620 3528
rect 108120 3476 108172 3528
rect 108948 3476 109000 3528
rect 109316 3476 109368 3528
rect 110328 3476 110380 3528
rect 110512 3476 110564 3528
rect 111524 3476 111576 3528
rect 114008 3476 114060 3528
rect 114468 3476 114520 3528
rect 115204 3476 115256 3528
rect 115848 3476 115900 3528
rect 116400 3476 116452 3528
rect 117044 3476 117096 3528
rect 117596 3476 117648 3528
rect 118608 3476 118660 3528
rect 118792 3476 118844 3528
rect 119988 3476 120040 3528
rect 123484 3476 123536 3528
rect 124128 3476 124180 3528
rect 129372 3476 129424 3528
rect 130384 3476 130436 3528
rect 202144 3476 202196 3528
rect 257068 3476 257120 3528
rect 313924 3476 313976 3528
rect 315028 3476 315080 3528
rect 316040 3476 316092 3528
rect 317328 3476 317380 3528
rect 324320 3476 324372 3528
rect 325608 3476 325660 3528
rect 336004 3476 336056 3528
rect 337476 3476 337528 3528
rect 340880 3476 340932 3528
rect 342168 3476 342220 3528
rect 350448 3476 350500 3528
rect 353300 3476 353352 3528
rect 582196 3476 582248 3528
rect 583484 3476 583536 3528
rect 6460 3408 6512 3460
rect 15844 3408 15896 3460
rect 26516 3408 26568 3460
rect 65524 3408 65576 3460
rect 66168 3408 66220 3460
rect 67916 3408 67968 3460
rect 68928 3408 68980 3460
rect 72608 3408 72660 3460
rect 73068 3408 73120 3460
rect 75000 3408 75052 3460
rect 75828 3408 75880 3460
rect 76196 3408 76248 3460
rect 77208 3408 77260 3460
rect 80888 3408 80940 3460
rect 81348 3408 81400 3460
rect 83280 3408 83332 3460
rect 84108 3408 84160 3460
rect 84476 3408 84528 3460
rect 85488 3408 85540 3460
rect 89168 3408 89220 3460
rect 89628 3408 89680 3460
rect 91560 3408 91612 3460
rect 92388 3408 92440 3460
rect 92756 3408 92808 3460
rect 93768 3408 93820 3460
rect 97448 3408 97500 3460
rect 97908 3408 97960 3460
rect 102232 3408 102284 3460
rect 123392 3408 123444 3460
rect 124680 3408 124732 3460
rect 214564 3408 214616 3460
rect 285404 3408 285456 3460
rect 306472 3408 306524 3460
rect 323584 3408 323636 3460
rect 332692 3408 332744 3460
rect 71044 3340 71096 3392
rect 78588 3340 78640 3392
rect 87604 3340 87656 3392
rect 122288 3272 122340 3324
rect 122748 3272 122800 3324
rect 346952 3272 347004 3324
rect 351920 3272 351972 3324
rect 280804 3136 280856 3188
rect 283104 3136 283156 3188
rect 269764 3068 269816 3120
rect 272432 3068 272484 3120
rect 347044 3068 347096 3120
rect 349252 3068 349304 3120
rect 90364 3000 90416 3052
rect 91008 3000 91060 3052
rect 581000 3000 581052 3052
rect 583392 3000 583444 3052
rect 93952 2932 94004 2984
rect 94964 2932 95016 2984
rect 51356 2116 51408 2168
rect 90272 2116 90324 2168
rect 198096 2116 198148 2168
rect 254676 2116 254728 2168
rect 7656 2048 7708 2100
rect 32312 2048 32364 2100
rect 87972 2048 88024 2100
rect 222844 2048 222896 2100
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 67640 703520 67692 703526
rect 72946 703520 73058 704960
rect 75828 703588 75880 703594
rect 75828 703530 75880 703536
rect 8128 702642 8156 703520
rect 8116 702636 8168 702642
rect 8116 702578 8168 702584
rect 24320 699718 24348 703520
rect 40512 700330 40540 703520
rect 67640 703462 67692 703468
rect 59268 703384 59320 703390
rect 59268 703326 59320 703332
rect 57888 702976 57940 702982
rect 57888 702918 57940 702924
rect 53748 702568 53800 702574
rect 53748 702510 53800 702516
rect 40500 700324 40552 700330
rect 40500 700266 40552 700272
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 25504 699712 25556 699718
rect 25504 699654 25556 699660
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 11704 683188 11756 683194
rect 11704 683130 11756 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3424 658144
rect 3476 658135 3478 658144
rect 7564 658164 7616 658170
rect 3424 658106 3476 658112
rect 7564 658106 7616 658112
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 2778 619168 2834 619177
rect 2778 619103 2780 619112
rect 2832 619103 2834 619112
rect 4804 619132 4856 619138
rect 2780 619074 2832 619080
rect 4804 619074 4856 619080
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3424 589960 3476 589966
rect 3424 589902 3476 589908
rect 3436 580009 3464 589902
rect 3422 580000 3478 580009
rect 3422 579935 3478 579944
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3330 553888 3386 553897
rect 3330 553823 3386 553832
rect 3344 553450 3372 553823
rect 3332 553444 3384 553450
rect 3332 553386 3384 553392
rect 3436 540258 3464 566879
rect 3424 540252 3476 540258
rect 3424 540194 3476 540200
rect 3424 538892 3476 538898
rect 3424 538834 3476 538840
rect 3436 527921 3464 538834
rect 4816 536110 4844 619074
rect 7576 592686 7604 658106
rect 7564 592680 7616 592686
rect 7564 592622 7616 592628
rect 11716 543046 11744 683130
rect 14464 670744 14516 670750
rect 14464 670686 14516 670692
rect 11704 543040 11756 543046
rect 11704 542982 11756 542988
rect 14476 541686 14504 670686
rect 17224 632120 17276 632126
rect 17224 632062 17276 632068
rect 17236 576162 17264 632062
rect 25516 596154 25544 699654
rect 25504 596148 25556 596154
rect 25504 596090 25556 596096
rect 52274 590744 52330 590753
rect 52274 590679 52330 590688
rect 50896 585200 50948 585206
rect 50896 585142 50948 585148
rect 48136 582412 48188 582418
rect 48136 582354 48188 582360
rect 17224 576156 17276 576162
rect 17224 576098 17276 576104
rect 34520 576156 34572 576162
rect 34520 576098 34572 576104
rect 34532 575550 34560 576098
rect 34520 575544 34572 575550
rect 34520 575486 34572 575492
rect 35808 575544 35860 575550
rect 35808 575486 35860 575492
rect 32404 553444 32456 553450
rect 32404 553386 32456 553392
rect 14464 541680 14516 541686
rect 14464 541622 14516 541628
rect 32416 538218 32444 553386
rect 32404 538212 32456 538218
rect 32404 538154 32456 538160
rect 4804 536104 4856 536110
rect 4804 536046 4856 536052
rect 7564 534744 7616 534750
rect 7564 534686 7616 534692
rect 5448 533384 5500 533390
rect 5448 533326 5500 533332
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3332 502104 3384 502110
rect 3332 502046 3384 502052
rect 3344 501809 3372 502046
rect 3330 501800 3386 501809
rect 3330 501735 3386 501744
rect 2778 462632 2834 462641
rect 2778 462567 2780 462576
rect 2832 462567 2834 462576
rect 2780 462538 2832 462544
rect 3436 451926 3464 527847
rect 3514 514856 3570 514865
rect 3514 514791 3516 514800
rect 3568 514791 3570 514800
rect 3516 514762 3568 514768
rect 4066 475688 4122 475697
rect 4066 475623 4122 475632
rect 4080 475386 4108 475623
rect 5460 475386 5488 533326
rect 7576 502110 7604 534686
rect 15844 530596 15896 530602
rect 15844 530538 15896 530544
rect 14464 514820 14516 514826
rect 14464 514762 14516 514768
rect 7564 502104 7616 502110
rect 7564 502046 7616 502052
rect 4068 475380 4120 475386
rect 4068 475322 4120 475328
rect 5448 475380 5500 475386
rect 5448 475322 5500 475328
rect 11704 475380 11756 475386
rect 11704 475322 11756 475328
rect 4804 462596 4856 462602
rect 4804 462538 4856 462544
rect 3424 451920 3476 451926
rect 3424 451862 3476 451868
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 4816 447846 4844 462538
rect 4804 447840 4856 447846
rect 4804 447782 4856 447788
rect 4804 444440 4856 444446
rect 4804 444382 4856 444388
rect 3146 423600 3202 423609
rect 3146 423535 3202 423544
rect 3160 422958 3188 423535
rect 3148 422952 3200 422958
rect 3148 422894 3200 422900
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 2780 398744 2832 398750
rect 2780 398686 2832 398692
rect 2792 397497 2820 398686
rect 2778 397488 2834 397497
rect 2778 397423 2834 397432
rect 3436 388793 3464 410479
rect 4816 398750 4844 444382
rect 4804 398744 4856 398750
rect 4804 398686 4856 398692
rect 11716 389230 11744 475322
rect 14476 451246 14504 514762
rect 14464 451240 14516 451246
rect 14464 451182 14516 451188
rect 14464 448588 14516 448594
rect 14464 448530 14516 448536
rect 11704 389224 11756 389230
rect 11704 389166 11756 389172
rect 3422 388784 3478 388793
rect 3422 388719 3478 388728
rect 3424 387116 3476 387122
rect 3424 387058 3476 387064
rect 3436 371385 3464 387058
rect 7564 382288 7616 382294
rect 7564 382230 7616 382236
rect 4804 381540 4856 381546
rect 4804 381482 4856 381488
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 2780 346316 2832 346322
rect 2780 346258 2832 346264
rect 2792 345409 2820 346258
rect 2778 345400 2834 345409
rect 2778 345335 2834 345344
rect 3436 334626 3464 371311
rect 3516 358624 3568 358630
rect 3516 358566 3568 358572
rect 3528 358465 3556 358566
rect 3514 358456 3570 358465
rect 3514 358391 3570 358400
rect 4816 346322 4844 381482
rect 7576 358630 7604 382230
rect 7564 358624 7616 358630
rect 7564 358566 7616 358572
rect 4804 346316 4856 346322
rect 4804 346258 4856 346264
rect 3424 334620 3476 334626
rect 3424 334562 3476 334568
rect 11704 334620 11756 334626
rect 11704 334562 11756 334568
rect 7562 328536 7618 328545
rect 7562 328471 7618 328480
rect 20 326392 72 326398
rect 20 326334 72 326340
rect 32 6769 60 326334
rect 4068 319456 4120 319462
rect 4068 319398 4120 319404
rect 4080 319297 4108 319398
rect 4066 319288 4122 319297
rect 4066 319223 4122 319232
rect 3424 306332 3476 306338
rect 3424 306274 3476 306280
rect 3436 306241 3464 306274
rect 3422 306232 3478 306241
rect 3422 306167 3478 306176
rect 2778 293176 2834 293185
rect 2778 293111 2834 293120
rect 2792 292874 2820 293111
rect 2780 292868 2832 292874
rect 2780 292810 2832 292816
rect 4080 269822 4108 319223
rect 4804 292868 4856 292874
rect 4804 292810 4856 292816
rect 4068 269816 4120 269822
rect 4068 269758 4120 269764
rect 3422 267200 3478 267209
rect 3422 267135 3478 267144
rect 3436 267034 3464 267135
rect 3424 267028 3476 267034
rect 3424 266970 3476 266976
rect 3424 255264 3476 255270
rect 3424 255206 3476 255212
rect 3436 254153 3464 255206
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3424 241120 3476 241126
rect 3422 241088 3424 241097
rect 3476 241088 3478 241097
rect 3422 241023 3478 241032
rect 4816 237386 4844 292810
rect 7576 241126 7604 328471
rect 11716 318102 11744 334562
rect 11704 318096 11756 318102
rect 11704 318038 11756 318044
rect 14476 292534 14504 448530
rect 15856 422958 15884 530538
rect 35820 454714 35848 575486
rect 41328 572756 41380 572762
rect 41328 572698 41380 572704
rect 37188 561740 37240 561746
rect 37188 561682 37240 561688
rect 35808 454708 35860 454714
rect 35808 454650 35860 454656
rect 37200 429146 37228 561682
rect 39948 543040 40000 543046
rect 39948 542982 40000 542988
rect 39960 542434 39988 542982
rect 39948 542428 40000 542434
rect 39948 542370 40000 542376
rect 36728 429140 36780 429146
rect 36728 429082 36780 429088
rect 37188 429140 37240 429146
rect 37188 429082 37240 429088
rect 36740 428466 36768 429082
rect 22744 428460 22796 428466
rect 22744 428402 22796 428408
rect 36728 428460 36780 428466
rect 36728 428402 36780 428408
rect 15844 422952 15896 422958
rect 15844 422894 15896 422900
rect 15856 391406 15884 422894
rect 15844 391400 15896 391406
rect 15844 391342 15896 391348
rect 15844 384328 15896 384334
rect 15844 384270 15896 384276
rect 15856 319462 15884 384270
rect 17224 330540 17276 330546
rect 17224 330482 17276 330488
rect 15844 319456 15896 319462
rect 15844 319398 15896 319404
rect 15844 294024 15896 294030
rect 15844 293966 15896 293972
rect 14464 292528 14516 292534
rect 14464 292470 14516 292476
rect 11704 278792 11756 278798
rect 11704 278734 11756 278740
rect 7564 241120 7616 241126
rect 7564 241062 7616 241068
rect 4804 237380 4856 237386
rect 4804 237322 4856 237328
rect 4804 221468 4856 221474
rect 4804 221410 4856 221416
rect 3332 215280 3384 215286
rect 3332 215222 3384 215228
rect 3344 214985 3372 215222
rect 3330 214976 3386 214985
rect 3330 214911 3386 214920
rect 3514 207632 3570 207641
rect 3514 207567 3570 207576
rect 3424 202836 3476 202842
rect 3424 202778 3476 202784
rect 3436 201929 3464 202778
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3528 200114 3556 207567
rect 3436 200086 3556 200114
rect 3240 164212 3292 164218
rect 3240 164154 3292 164160
rect 3252 162897 3280 164154
rect 3238 162888 3294 162897
rect 3238 162823 3294 162832
rect 2780 150340 2832 150346
rect 2780 150282 2832 150288
rect 2792 149841 2820 150282
rect 2778 149832 2834 149841
rect 2778 149767 2834 149776
rect 3436 110673 3464 200086
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3528 188873 3556 188974
rect 3514 188864 3570 188873
rect 3514 188799 3570 188808
rect 4816 150346 4844 221410
rect 4804 150340 4856 150346
rect 4804 150282 4856 150288
rect 3516 137964 3568 137970
rect 3516 137906 3568 137912
rect 3528 136785 3556 137906
rect 3514 136776 3570 136785
rect 3514 136711 3570 136720
rect 3422 110664 3478 110673
rect 3422 110599 3478 110608
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 11716 85542 11744 278734
rect 15856 164218 15884 293966
rect 15844 164212 15896 164218
rect 15844 164154 15896 164160
rect 17236 97986 17264 330482
rect 18604 307828 18656 307834
rect 18604 307770 18656 307776
rect 18616 255270 18644 307770
rect 21456 269816 21508 269822
rect 21456 269758 21508 269764
rect 21088 269068 21140 269074
rect 21088 269010 21140 269016
rect 21100 267734 21128 269010
rect 21100 267706 21404 267734
rect 21376 267034 21404 267706
rect 21364 267028 21416 267034
rect 21364 266970 21416 266976
rect 18604 255264 18656 255270
rect 18604 255206 18656 255212
rect 21376 234598 21404 266970
rect 21468 261526 21496 269758
rect 22756 269074 22784 428402
rect 39960 396778 39988 542370
rect 41340 449177 41368 572698
rect 44088 560312 44140 560318
rect 44088 560254 44140 560260
rect 44100 511290 44128 560254
rect 45468 536104 45520 536110
rect 45468 536046 45520 536052
rect 44088 511284 44140 511290
rect 44088 511226 44140 511232
rect 41326 449168 41382 449177
rect 41326 449103 41382 449112
rect 41328 445868 41380 445874
rect 41328 445810 41380 445816
rect 39948 396772 40000 396778
rect 39948 396714 40000 396720
rect 36544 329112 36596 329118
rect 36544 329054 36596 329060
rect 32402 328672 32458 328681
rect 32402 328607 32458 328616
rect 22744 269068 22796 269074
rect 22744 269010 22796 269016
rect 21456 261520 21508 261526
rect 21456 261462 21508 261468
rect 21364 234592 21416 234598
rect 21364 234534 21416 234540
rect 32416 137970 32444 328607
rect 33782 327448 33838 327457
rect 33782 327383 33838 327392
rect 32404 137964 32456 137970
rect 32404 137906 32456 137912
rect 17224 97980 17276 97986
rect 17224 97922 17276 97928
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 11704 85536 11756 85542
rect 11704 85478 11756 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 30286 83464 30342 83473
rect 30286 83399 30342 83408
rect 12346 80744 12402 80753
rect 12346 80679 12402 80688
rect 5446 79520 5502 79529
rect 5446 79455 5502 79464
rect 3424 71732 3476 71738
rect 3424 71674 3476 71680
rect 3436 71641 3464 71674
rect 3422 71632 3478 71641
rect 3422 71567 3478 71576
rect 3056 59356 3108 59362
rect 3056 59298 3108 59304
rect 3068 58585 3096 59298
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 3424 45552 3476 45558
rect 3422 45520 3424 45529
rect 3476 45520 3478 45529
rect 3422 45455 3478 45464
rect 4068 35284 4120 35290
rect 4068 35226 4120 35232
rect 3148 33108 3200 33114
rect 3148 33050 3200 33056
rect 3160 32473 3188 33050
rect 3146 32464 3202 32473
rect 3146 32399 3202 32408
rect 1400 28280 1452 28286
rect 1400 28222 1452 28228
rect 110 24168 166 24177
rect 110 24103 166 24112
rect 18 6760 74 6769
rect 18 6695 74 6704
rect 124 490 152 24103
rect 1412 16574 1440 28222
rect 3974 25528 4030 25537
rect 3974 25463 4030 25472
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 1412 16546 1716 16574
rect 400 598 612 626
rect 400 490 428 598
rect 124 462 428 490
rect 584 480 612 598
rect 1688 480 1716 16546
rect 3988 3534 4016 25463
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 2884 480 2912 3470
rect 4080 480 4108 35226
rect 5460 6914 5488 79455
rect 10966 51776 11022 51785
rect 10966 51711 11022 51720
rect 9588 10328 9640 10334
rect 9588 10270 9640 10276
rect 5276 6886 5488 6914
rect 5276 480 5304 6886
rect 9600 3534 9628 10270
rect 10980 3534 11008 51711
rect 12164 14476 12216 14482
rect 12164 14418 12216 14424
rect 11152 3596 11204 3602
rect 11152 3538 11204 3544
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9956 3528 10008 3534
rect 9956 3470 10008 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6472 480 6500 3402
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 7668 480 7696 2042
rect 8772 480 8800 3470
rect 9968 480 9996 3470
rect 11164 480 11192 3538
rect 12176 3482 12204 14418
rect 12360 6914 12388 80679
rect 15842 79384 15898 79393
rect 15842 79319 15898 79328
rect 13726 77888 13782 77897
rect 13726 77823 13782 77832
rect 13740 6914 13768 77823
rect 15106 66872 15162 66881
rect 15106 66807 15162 66816
rect 15120 6914 15148 66807
rect 12268 6886 12388 6914
rect 13556 6886 13768 6914
rect 14752 6886 15148 6914
rect 12268 3602 12296 6886
rect 12256 3596 12308 3602
rect 12256 3538 12308 3544
rect 12176 3454 12388 3482
rect 12360 480 12388 3454
rect 13556 480 13584 6886
rect 14752 480 14780 6886
rect 15856 3466 15884 79319
rect 19246 75168 19302 75177
rect 19246 75103 19302 75112
rect 17866 55856 17922 55865
rect 17866 55791 17922 55800
rect 17880 3534 17908 55791
rect 19260 3534 19288 75103
rect 23386 73808 23442 73817
rect 23386 73743 23442 73752
rect 20534 59936 20590 59945
rect 20534 59871 20590 59880
rect 20548 3534 20576 59871
rect 22008 46232 22060 46238
rect 22008 46174 22060 46180
rect 22020 6914 22048 46174
rect 23400 6914 23428 73743
rect 26146 68232 26202 68241
rect 26146 68167 26202 68176
rect 24766 39264 24822 39273
rect 24766 39199 24822 39208
rect 21836 6886 22048 6914
rect 23032 6886 23428 6914
rect 20628 4820 20680 4826
rect 20628 4762 20680 4768
rect 17040 3528 17092 3534
rect 17040 3470 17092 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 18236 3528 18288 3534
rect 18236 3470 18288 3476
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 20536 3528 20588 3534
rect 20536 3470 20588 3476
rect 15844 3460 15896 3466
rect 15844 3402 15896 3408
rect 15934 3360 15990 3369
rect 15934 3295 15990 3304
rect 15948 480 15976 3295
rect 17052 480 17080 3470
rect 18248 480 18276 3470
rect 19444 480 19472 3470
rect 20640 480 20668 4762
rect 21836 480 21864 6886
rect 23032 480 23060 6886
rect 24780 3534 24808 39199
rect 26160 3534 26188 68167
rect 28906 26888 28962 26897
rect 28906 26823 28962 26832
rect 28814 21312 28870 21321
rect 28814 21247 28870 21256
rect 28828 3534 28856 21247
rect 24216 3528 24268 3534
rect 24216 3470 24268 3476
rect 24768 3528 24820 3534
rect 24768 3470 24820 3476
rect 25320 3528 25372 3534
rect 25320 3470 25372 3476
rect 26148 3528 26200 3534
rect 26148 3470 26200 3476
rect 27712 3528 27764 3534
rect 27712 3470 27764 3476
rect 28816 3528 28868 3534
rect 28816 3470 28868 3476
rect 24228 480 24256 3470
rect 25332 480 25360 3470
rect 26516 3460 26568 3466
rect 26516 3402 26568 3408
rect 26528 480 26556 3402
rect 27724 480 27752 3470
rect 28920 480 28948 26823
rect 30300 6914 30328 83399
rect 33046 62792 33102 62801
rect 33046 62727 33102 62736
rect 32402 58712 32458 58721
rect 32402 58647 32458 58656
rect 31668 47592 31720 47598
rect 31668 47534 31720 47540
rect 31680 6914 31708 47534
rect 32416 6914 32444 58647
rect 30116 6886 30328 6914
rect 31312 6886 31708 6914
rect 32324 6886 32444 6914
rect 30116 480 30144 6886
rect 31312 480 31340 6886
rect 32324 2106 32352 6886
rect 33060 3534 33088 62727
rect 33796 59362 33824 327383
rect 35256 314696 35308 314702
rect 35256 314638 35308 314644
rect 35268 189038 35296 314638
rect 36556 306338 36584 329054
rect 40682 327312 40738 327321
rect 40682 327247 40738 327256
rect 39304 307080 39356 307086
rect 39304 307022 39356 307028
rect 36544 306332 36596 306338
rect 36544 306274 36596 306280
rect 36542 223000 36598 223009
rect 36542 222935 36598 222944
rect 35256 189032 35308 189038
rect 35256 188974 35308 188980
rect 35164 188352 35216 188358
rect 35164 188294 35216 188300
rect 33784 59356 33836 59362
rect 33784 59298 33836 59304
rect 34428 43444 34480 43450
rect 34428 43386 34480 43392
rect 34440 3534 34468 43386
rect 35176 33114 35204 188294
rect 35806 69592 35862 69601
rect 35806 69527 35862 69536
rect 35164 33108 35216 33114
rect 35164 33050 35216 33056
rect 35820 3534 35848 69527
rect 36556 45558 36584 222935
rect 39316 71738 39344 307022
rect 40696 215286 40724 327247
rect 41144 264988 41196 264994
rect 41144 264930 41196 264936
rect 40684 215280 40736 215286
rect 40684 215222 40736 215228
rect 41156 72457 41184 264930
rect 41340 264246 41368 445810
rect 44100 425746 44128 511226
rect 44088 425740 44140 425746
rect 44088 425682 44140 425688
rect 43996 398132 44048 398138
rect 43996 398074 44048 398080
rect 41328 264240 41380 264246
rect 41328 264182 41380 264188
rect 44008 240145 44036 398074
rect 45480 387802 45508 536046
rect 48148 449206 48176 582354
rect 49608 571396 49660 571402
rect 49608 571338 49660 571344
rect 48228 557592 48280 557598
rect 48228 557534 48280 557540
rect 48136 449200 48188 449206
rect 48136 449142 48188 449148
rect 48136 430636 48188 430642
rect 48136 430578 48188 430584
rect 45468 387796 45520 387802
rect 45468 387738 45520 387744
rect 44088 329860 44140 329866
rect 44088 329802 44140 329808
rect 43994 240136 44050 240145
rect 43994 240071 44050 240080
rect 41234 82104 41290 82113
rect 41234 82039 41290 82048
rect 41142 72448 41198 72457
rect 41142 72383 41198 72392
rect 39304 71732 39356 71738
rect 39304 71674 39356 71680
rect 38566 50280 38622 50289
rect 38566 50215 38622 50224
rect 37186 48920 37242 48929
rect 37186 48855 37242 48864
rect 36544 45552 36596 45558
rect 36544 45494 36596 45500
rect 37096 31068 37148 31074
rect 37096 31010 37148 31016
rect 37108 16574 37136 31010
rect 37016 16546 37136 16574
rect 35992 3596 36044 3602
rect 35992 3538 36044 3544
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 33048 3528 33100 3534
rect 33048 3470 33100 3476
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 34796 3528 34848 3534
rect 34796 3470 34848 3476
rect 35808 3528 35860 3534
rect 35808 3470 35860 3476
rect 32312 2100 32364 2106
rect 32312 2042 32364 2048
rect 32416 480 32444 3470
rect 33612 480 33640 3470
rect 34808 480 34836 3470
rect 36004 480 36032 3538
rect 37016 3482 37044 16546
rect 37200 6914 37228 48855
rect 38580 6914 38608 50215
rect 39948 22772 40000 22778
rect 39948 22714 40000 22720
rect 39960 6914 39988 22714
rect 37108 6886 37228 6914
rect 38396 6886 38608 6914
rect 39592 6886 39988 6914
rect 37108 3602 37136 6886
rect 37096 3596 37148 3602
rect 37096 3538 37148 3544
rect 37016 3454 37228 3482
rect 37200 480 37228 3454
rect 38396 480 38424 6886
rect 39592 480 39620 6886
rect 41248 3534 41276 82039
rect 43994 76528 44050 76537
rect 43994 76463 44050 76472
rect 41878 7712 41934 7721
rect 41878 7647 41934 7656
rect 40684 3528 40736 3534
rect 40684 3470 40736 3476
rect 41236 3528 41288 3534
rect 41236 3470 41288 3476
rect 40696 480 40724 3470
rect 41892 480 41920 7647
rect 44008 3534 44036 76463
rect 44100 32434 44128 329802
rect 46848 318096 46900 318102
rect 46848 318038 46900 318044
rect 46860 317490 46888 318038
rect 46848 317484 46900 317490
rect 46848 317426 46900 317432
rect 46860 200122 46888 317426
rect 48148 235793 48176 430578
rect 48240 421598 48268 557534
rect 49620 453354 49648 571338
rect 50804 463004 50856 463010
rect 50804 462946 50856 462952
rect 49608 453348 49660 453354
rect 49608 453290 49660 453296
rect 49608 447160 49660 447166
rect 49608 447102 49660 447108
rect 48228 421592 48280 421598
rect 48228 421534 48280 421540
rect 49620 329118 49648 447102
rect 50816 380866 50844 462946
rect 50908 457502 50936 585142
rect 50988 564392 51040 564398
rect 50988 564334 51040 564340
rect 50896 457496 50948 457502
rect 50896 457438 50948 457444
rect 51000 431934 51028 564334
rect 52288 465730 52316 590679
rect 53656 566500 53708 566506
rect 53656 566442 53708 566448
rect 52368 545080 52420 545086
rect 52368 545022 52420 545028
rect 52276 465724 52328 465730
rect 52276 465666 52328 465672
rect 52276 461644 52328 461650
rect 52276 461586 52328 461592
rect 50988 431928 51040 431934
rect 50988 431870 51040 431876
rect 51000 430642 51028 431870
rect 50988 430636 51040 430642
rect 50988 430578 51040 430584
rect 50896 401600 50948 401606
rect 50896 401542 50948 401548
rect 50804 380860 50856 380866
rect 50804 380802 50856 380808
rect 50804 361548 50856 361554
rect 50804 361490 50856 361496
rect 49608 329112 49660 329118
rect 49608 329054 49660 329060
rect 49608 308440 49660 308446
rect 49608 308382 49660 308388
rect 49620 307834 49648 308382
rect 49608 307828 49660 307834
rect 49608 307770 49660 307776
rect 48228 270564 48280 270570
rect 48228 270506 48280 270512
rect 48134 235784 48190 235793
rect 48134 235719 48190 235728
rect 46848 200116 46900 200122
rect 46848 200058 46900 200064
rect 45468 42084 45520 42090
rect 45468 42026 45520 42032
rect 44088 32428 44140 32434
rect 44088 32370 44140 32376
rect 45282 15872 45338 15881
rect 45282 15807 45338 15816
rect 44272 3596 44324 3602
rect 44272 3538 44324 3544
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 43996 3528 44048 3534
rect 43996 3470 44048 3476
rect 43088 480 43116 3470
rect 44284 480 44312 3538
rect 45296 3482 45324 15807
rect 45480 6914 45508 42026
rect 46848 40724 46900 40730
rect 46848 40666 46900 40672
rect 46860 6914 46888 40666
rect 48240 19990 48268 270506
rect 49620 231849 49648 307770
rect 49606 231840 49662 231849
rect 49606 231775 49662 231784
rect 50816 222086 50844 361490
rect 50908 240009 50936 401542
rect 52288 378146 52316 461586
rect 52380 398138 52408 545022
rect 53668 435402 53696 566442
rect 53760 564398 53788 702510
rect 55036 574796 55088 574802
rect 55036 574738 55088 574744
rect 53748 564392 53800 564398
rect 53748 564334 53800 564340
rect 53748 547188 53800 547194
rect 53748 547130 53800 547136
rect 53656 435396 53708 435402
rect 53656 435338 53708 435344
rect 53668 431954 53696 435338
rect 53576 431926 53696 431954
rect 52368 398132 52420 398138
rect 52368 398074 52420 398080
rect 52366 385656 52422 385665
rect 52366 385591 52422 385600
rect 52276 378140 52328 378146
rect 52276 378082 52328 378088
rect 52276 312588 52328 312594
rect 52276 312530 52328 312536
rect 52184 287088 52236 287094
rect 52184 287030 52236 287036
rect 50988 247104 51040 247110
rect 50988 247046 51040 247052
rect 50894 240000 50950 240009
rect 50894 239935 50950 239944
rect 50528 222080 50580 222086
rect 50528 222022 50580 222028
rect 50804 222080 50856 222086
rect 50804 222022 50856 222028
rect 50540 221474 50568 222022
rect 50528 221468 50580 221474
rect 50528 221410 50580 221416
rect 50894 72584 50950 72593
rect 50894 72519 50950 72528
rect 49608 37936 49660 37942
rect 49608 37878 49660 37884
rect 48228 19984 48280 19990
rect 48228 19926 48280 19932
rect 45388 6886 45508 6914
rect 46676 6886 46888 6914
rect 45388 3602 45416 6886
rect 45376 3596 45428 3602
rect 45376 3538 45428 3544
rect 45296 3454 45508 3482
rect 45480 480 45508 3454
rect 46676 480 46704 6886
rect 47860 6180 47912 6186
rect 47860 6122 47912 6128
rect 47872 480 47900 6122
rect 49620 3534 49648 37878
rect 50908 3534 50936 72519
rect 51000 44878 51028 247046
rect 51722 224224 51778 224233
rect 51722 224159 51778 224168
rect 50988 44872 51040 44878
rect 50988 44814 51040 44820
rect 51736 20670 51764 224159
rect 52196 218754 52224 287030
rect 52288 226273 52316 312530
rect 52380 262886 52408 385591
rect 53576 376786 53604 431926
rect 53760 402974 53788 547130
rect 54852 468512 54904 468518
rect 54852 468454 54904 468460
rect 53668 402946 53788 402974
rect 53668 402286 53696 402946
rect 53656 402280 53708 402286
rect 53656 402222 53708 402228
rect 53564 376780 53616 376786
rect 53564 376722 53616 376728
rect 53564 309188 53616 309194
rect 53564 309130 53616 309136
rect 53472 276072 53524 276078
rect 53472 276014 53524 276020
rect 52368 262880 52420 262886
rect 52368 262822 52420 262828
rect 52274 226264 52330 226273
rect 52274 226199 52330 226208
rect 52184 218748 52236 218754
rect 52184 218690 52236 218696
rect 52380 202881 52408 262822
rect 53484 213897 53512 276014
rect 53470 213888 53526 213897
rect 53470 213823 53526 213832
rect 53576 206961 53604 309130
rect 53668 244934 53696 402222
rect 53748 376780 53800 376786
rect 53748 376722 53800 376728
rect 53760 296682 53788 376722
rect 54864 361554 54892 468454
rect 55048 454782 55076 574738
rect 57704 567248 57756 567254
rect 57704 567190 57756 567196
rect 56508 558952 56560 558958
rect 56508 558894 56560 558900
rect 55128 539640 55180 539646
rect 55128 539582 55180 539588
rect 55036 454776 55088 454782
rect 55036 454718 55088 454724
rect 54944 444508 54996 444514
rect 54944 444450 54996 444456
rect 54852 361548 54904 361554
rect 54852 361490 54904 361496
rect 54852 352572 54904 352578
rect 54852 352514 54904 352520
rect 53748 296676 53800 296682
rect 53748 296618 53800 296624
rect 53748 258120 53800 258126
rect 53748 258062 53800 258068
rect 53656 244928 53708 244934
rect 53656 244870 53708 244876
rect 53562 206952 53618 206961
rect 53562 206887 53618 206896
rect 52366 202872 52422 202881
rect 52366 202807 52422 202816
rect 53654 54496 53710 54505
rect 53654 54431 53710 54440
rect 53564 35216 53616 35222
rect 53564 35158 53616 35164
rect 51724 20664 51776 20670
rect 51724 20606 51776 20612
rect 53576 3534 53604 35158
rect 53668 16574 53696 54431
rect 53760 33794 53788 258062
rect 53840 237380 53892 237386
rect 53840 237322 53892 237328
rect 53852 236706 53880 237322
rect 54864 236706 54892 352514
rect 54956 253910 54984 444450
rect 55140 393310 55168 539582
rect 56520 538214 56548 558894
rect 56428 538186 56548 538214
rect 56428 534070 56456 538186
rect 56416 534064 56468 534070
rect 56416 534006 56468 534012
rect 56428 424386 56456 534006
rect 56508 440904 56560 440910
rect 56508 440846 56560 440852
rect 56416 424380 56468 424386
rect 56416 424322 56468 424328
rect 55128 393304 55180 393310
rect 55128 393246 55180 393252
rect 56520 327078 56548 440846
rect 57716 437510 57744 567190
rect 57796 545760 57848 545766
rect 57796 545702 57848 545708
rect 57704 437504 57756 437510
rect 57704 437446 57756 437452
rect 57704 425128 57756 425134
rect 57704 425070 57756 425076
rect 57612 406564 57664 406570
rect 57612 406506 57664 406512
rect 57624 401606 57652 406506
rect 57612 401600 57664 401606
rect 57612 401542 57664 401548
rect 57716 366353 57744 425070
rect 57808 406570 57836 545702
rect 57900 545086 57928 702918
rect 59176 586560 59228 586566
rect 59176 586502 59228 586508
rect 58992 554804 59044 554810
rect 58992 554746 59044 554752
rect 57888 545080 57940 545086
rect 57888 545022 57940 545028
rect 57888 425740 57940 425746
rect 57888 425682 57940 425688
rect 57900 425134 57928 425682
rect 57888 425128 57940 425134
rect 57888 425070 57940 425076
rect 59004 416838 59032 554746
rect 59084 464364 59136 464370
rect 59084 464306 59136 464312
rect 58992 416832 59044 416838
rect 58992 416774 59044 416780
rect 57888 414724 57940 414730
rect 57888 414666 57940 414672
rect 57796 406564 57848 406570
rect 57796 406506 57848 406512
rect 57702 366344 57758 366353
rect 57702 366279 57758 366288
rect 55956 327072 56008 327078
rect 55956 327014 56008 327020
rect 56508 327072 56560 327078
rect 56508 327014 56560 327020
rect 55968 326398 55996 327014
rect 55956 326392 56008 326398
rect 55956 326334 56008 326340
rect 56508 318844 56560 318850
rect 56508 318786 56560 318792
rect 55128 285728 55180 285734
rect 55128 285670 55180 285676
rect 55036 268388 55088 268394
rect 55036 268330 55088 268336
rect 54944 253904 54996 253910
rect 54944 253846 54996 253852
rect 54944 253224 54996 253230
rect 54944 253166 54996 253172
rect 53840 236700 53892 236706
rect 53840 236642 53892 236648
rect 54852 236700 54904 236706
rect 54852 236642 54904 236648
rect 54956 231810 54984 253166
rect 54944 231804 54996 231810
rect 54944 231746 54996 231752
rect 53748 33788 53800 33794
rect 53748 33730 53800 33736
rect 54944 31136 54996 31142
rect 54944 31078 54996 31084
rect 53668 16546 53788 16574
rect 48964 3528 49016 3534
rect 48964 3470 49016 3476
rect 49608 3528 49660 3534
rect 49608 3470 49660 3476
rect 50160 3528 50212 3534
rect 50160 3470 50212 3476
rect 50896 3528 50948 3534
rect 50896 3470 50948 3476
rect 52552 3528 52604 3534
rect 52552 3470 52604 3476
rect 53564 3528 53616 3534
rect 53564 3470 53616 3476
rect 48976 480 49004 3470
rect 50172 480 50200 3470
rect 51356 2168 51408 2174
rect 51356 2110 51408 2116
rect 51368 480 51396 2110
rect 52564 480 52592 3470
rect 53760 480 53788 16546
rect 54956 480 54984 31078
rect 55048 17241 55076 268330
rect 55140 18630 55168 285670
rect 56416 274712 56468 274718
rect 56416 274654 56468 274660
rect 56324 253972 56376 253978
rect 56324 253914 56376 253920
rect 56336 227050 56364 253914
rect 56324 227044 56376 227050
rect 56324 226986 56376 226992
rect 56428 195974 56456 274654
rect 56416 195968 56468 195974
rect 56416 195910 56468 195916
rect 56520 69737 56548 318786
rect 57796 284980 57848 284986
rect 57796 284922 57848 284928
rect 57704 277432 57756 277438
rect 57704 277374 57756 277380
rect 57152 253904 57204 253910
rect 57152 253846 57204 253852
rect 57164 252618 57192 253846
rect 57152 252612 57204 252618
rect 57152 252554 57204 252560
rect 57612 252612 57664 252618
rect 57612 252554 57664 252560
rect 57624 222018 57652 252554
rect 57716 233238 57744 277374
rect 57704 233232 57756 233238
rect 57704 233174 57756 233180
rect 57808 225622 57836 284922
rect 57900 241505 57928 414666
rect 57980 403640 58032 403646
rect 57980 403582 58032 403588
rect 57992 402286 58020 403582
rect 57980 402280 58032 402286
rect 57980 402222 58032 402228
rect 59096 388929 59124 464306
rect 59188 458862 59216 586502
rect 59280 554742 59308 703326
rect 61844 703180 61896 703186
rect 61844 703122 61896 703128
rect 60648 564460 60700 564466
rect 60648 564402 60700 564408
rect 59268 554736 59320 554742
rect 59268 554678 59320 554684
rect 59176 458856 59228 458862
rect 59176 458798 59228 458804
rect 59174 445904 59230 445913
rect 59174 445839 59230 445848
rect 59082 388920 59138 388929
rect 59082 388855 59138 388864
rect 59188 351937 59216 445839
rect 60556 437504 60608 437510
rect 60556 437446 60608 437452
rect 59266 411360 59322 411369
rect 59266 411295 59322 411304
rect 59174 351928 59230 351937
rect 59174 351863 59230 351872
rect 58900 299532 58952 299538
rect 58900 299474 58952 299480
rect 57886 241496 57942 241505
rect 57886 241431 57942 241440
rect 57796 225616 57848 225622
rect 57796 225558 57848 225564
rect 57612 222012 57664 222018
rect 57612 221954 57664 221960
rect 58912 198014 58940 299474
rect 59188 293962 59216 351863
rect 59280 331226 59308 411295
rect 60004 399492 60056 399498
rect 60004 399434 60056 399440
rect 60016 398138 60044 399434
rect 60004 398132 60056 398138
rect 60004 398074 60056 398080
rect 60568 353977 60596 437446
rect 60660 432070 60688 564402
rect 61856 547806 61884 703122
rect 66168 702500 66220 702506
rect 66168 702442 66220 702448
rect 61936 590708 61988 590714
rect 61936 590650 61988 590656
rect 61844 547800 61896 547806
rect 61844 547742 61896 547748
rect 61856 547194 61884 547742
rect 61844 547188 61896 547194
rect 61844 547130 61896 547136
rect 61752 457564 61804 457570
rect 61752 457506 61804 457512
rect 60648 432064 60700 432070
rect 60648 432006 60700 432012
rect 60660 373318 60688 432006
rect 61384 421592 61436 421598
rect 61384 421534 61436 421540
rect 60648 373312 60700 373318
rect 60648 373254 60700 373260
rect 60554 353968 60610 353977
rect 60554 353903 60610 353912
rect 60556 353388 60608 353394
rect 60556 353330 60608 353336
rect 60464 331900 60516 331906
rect 60464 331842 60516 331848
rect 59268 331220 59320 331226
rect 59268 331162 59320 331168
rect 59280 330546 59308 331162
rect 59268 330540 59320 330546
rect 59268 330482 59320 330488
rect 59268 324352 59320 324358
rect 59268 324294 59320 324300
rect 59176 293956 59228 293962
rect 59176 293898 59228 293904
rect 59084 278792 59136 278798
rect 59084 278734 59136 278740
rect 58992 264240 59044 264246
rect 58992 264182 59044 264188
rect 59004 237969 59032 264182
rect 58990 237960 59046 237969
rect 58990 237895 59046 237904
rect 59096 220833 59124 278734
rect 59082 220824 59138 220833
rect 59082 220759 59138 220768
rect 58900 198008 58952 198014
rect 58900 197950 58952 197956
rect 56506 69728 56562 69737
rect 56506 69663 56562 69672
rect 57886 53136 57942 53145
rect 57886 53071 57942 53080
rect 56508 36576 56560 36582
rect 56508 36518 56560 36524
rect 55128 18624 55180 18630
rect 55128 18566 55180 18572
rect 55034 17232 55090 17241
rect 55034 17167 55090 17176
rect 56520 3534 56548 36518
rect 57900 3534 57928 53071
rect 59176 29708 59228 29714
rect 59176 29650 59228 29656
rect 59188 3534 59216 29650
rect 59280 22681 59308 324294
rect 60476 292534 60504 331842
rect 60568 313274 60596 353330
rect 60648 317552 60700 317558
rect 60648 317494 60700 317500
rect 60556 313268 60608 313274
rect 60556 313210 60608 313216
rect 60464 292528 60516 292534
rect 60464 292470 60516 292476
rect 60556 281580 60608 281586
rect 60556 281522 60608 281528
rect 60464 263628 60516 263634
rect 60464 263570 60516 263576
rect 60372 249824 60424 249830
rect 60372 249766 60424 249772
rect 60384 238134 60412 249766
rect 60372 238128 60424 238134
rect 60372 238070 60424 238076
rect 60476 223553 60504 263570
rect 60568 237153 60596 281522
rect 60554 237144 60610 237153
rect 60554 237079 60610 237088
rect 60462 223544 60518 223553
rect 60462 223479 60518 223488
rect 60660 71097 60688 317494
rect 61396 313177 61424 421534
rect 61764 389298 61792 457506
rect 61948 456074 61976 590650
rect 63316 587920 63368 587926
rect 63316 587862 63368 587868
rect 62028 547936 62080 547942
rect 62028 547878 62080 547884
rect 61936 456068 61988 456074
rect 61936 456010 61988 456016
rect 61844 451988 61896 451994
rect 61844 451930 61896 451936
rect 61752 389292 61804 389298
rect 61752 389234 61804 389240
rect 61856 386374 61884 451930
rect 62040 405822 62068 547878
rect 63328 460970 63356 587862
rect 64696 581052 64748 581058
rect 64696 580994 64748 581000
rect 63408 549296 63460 549302
rect 63408 549238 63460 549244
rect 63316 460964 63368 460970
rect 63316 460906 63368 460912
rect 63328 451274 63356 460906
rect 63236 451246 63356 451274
rect 62028 405816 62080 405822
rect 62028 405758 62080 405764
rect 61844 386368 61896 386374
rect 61844 386310 61896 386316
rect 63236 362234 63264 451246
rect 63316 416832 63368 416838
rect 63316 416774 63368 416780
rect 63224 362228 63276 362234
rect 63224 362170 63276 362176
rect 62028 342372 62080 342378
rect 62028 342314 62080 342320
rect 61844 335436 61896 335442
rect 61844 335378 61896 335384
rect 61856 315994 61884 335378
rect 61936 322992 61988 322998
rect 61936 322934 61988 322940
rect 61844 315988 61896 315994
rect 61844 315930 61896 315936
rect 61844 314220 61896 314226
rect 61844 314162 61896 314168
rect 61106 313168 61162 313177
rect 61106 313103 61162 313112
rect 61382 313168 61438 313177
rect 61382 313103 61438 313112
rect 61120 312594 61148 313103
rect 61108 312588 61160 312594
rect 61108 312530 61160 312536
rect 61752 294092 61804 294098
rect 61752 294034 61804 294040
rect 61764 214606 61792 294034
rect 61856 233209 61884 314162
rect 61842 233200 61898 233209
rect 61842 233135 61898 233144
rect 61752 214600 61804 214606
rect 61752 214542 61804 214548
rect 61948 199345 61976 322934
rect 62040 311846 62068 342314
rect 62028 311840 62080 311846
rect 62028 311782 62080 311788
rect 63328 289950 63356 416774
rect 63420 408474 63448 549238
rect 64708 460222 64736 580994
rect 66074 579728 66130 579737
rect 66074 579663 66130 579672
rect 64788 568608 64840 568614
rect 64788 568550 64840 568556
rect 64696 460216 64748 460222
rect 64696 460158 64748 460164
rect 64696 458924 64748 458930
rect 64696 458866 64748 458872
rect 64604 449268 64656 449274
rect 64604 449210 64656 449216
rect 63408 408468 63460 408474
rect 63408 408410 63460 408416
rect 64616 387705 64644 449210
rect 64708 388482 64736 458866
rect 64800 439074 64828 568550
rect 65524 554736 65576 554742
rect 65524 554678 65576 554684
rect 64788 439068 64840 439074
rect 64788 439010 64840 439016
rect 65536 415206 65564 554678
rect 66088 532030 66116 579663
rect 66180 546417 66208 702442
rect 67456 599616 67508 599622
rect 67456 599558 67508 599564
rect 66810 588296 66866 588305
rect 66810 588231 66866 588240
rect 66824 587926 66852 588231
rect 66812 587920 66864 587926
rect 66812 587862 66864 587868
rect 66260 586560 66312 586566
rect 66258 586528 66260 586537
rect 66312 586528 66314 586537
rect 66258 586463 66314 586472
rect 66810 582448 66866 582457
rect 66810 582383 66812 582392
rect 66864 582383 66866 582392
rect 66812 582354 66864 582360
rect 66994 581088 67050 581097
rect 66994 581023 66996 581032
rect 67048 581023 67050 581032
rect 66996 580994 67048 581000
rect 66902 575648 66958 575657
rect 66902 575583 66958 575592
rect 66916 575550 66944 575583
rect 66904 575544 66956 575550
rect 66904 575486 66956 575492
rect 67468 575385 67496 599558
rect 67548 596828 67600 596834
rect 67548 596770 67600 596776
rect 67454 575376 67510 575385
rect 67454 575311 67510 575320
rect 67468 574802 67496 575311
rect 67456 574796 67508 574802
rect 67456 574738 67508 574744
rect 66442 573200 66498 573209
rect 66442 573135 66498 573144
rect 66456 572762 66484 573135
rect 66444 572756 66496 572762
rect 66444 572698 66496 572704
rect 66442 571840 66498 571849
rect 66442 571775 66498 571784
rect 66456 571402 66484 571775
rect 66444 571396 66496 571402
rect 66444 571338 66496 571344
rect 67270 570208 67326 570217
rect 67270 570143 67326 570152
rect 66810 568848 66866 568857
rect 66810 568783 66866 568792
rect 66824 568614 66852 568783
rect 66812 568608 66864 568614
rect 66812 568550 66864 568556
rect 66902 567488 66958 567497
rect 66902 567423 66958 567432
rect 66916 567254 66944 567423
rect 66904 567248 66956 567254
rect 66904 567190 66956 567196
rect 66626 564632 66682 564641
rect 66626 564567 66682 564576
rect 66640 564466 66668 564567
rect 66628 564460 66680 564466
rect 66628 564402 66680 564408
rect 66444 564392 66496 564398
rect 66444 564334 66496 564340
rect 66456 564097 66484 564334
rect 66442 564088 66498 564097
rect 66442 564023 66498 564032
rect 66442 562048 66498 562057
rect 66442 561983 66498 561992
rect 66456 561746 66484 561983
rect 66444 561740 66496 561746
rect 66444 561682 66496 561688
rect 66626 560416 66682 560425
rect 66626 560351 66682 560360
rect 66640 560318 66668 560351
rect 66628 560312 66680 560318
rect 66628 560254 66680 560260
rect 66626 559056 66682 559065
rect 66626 558991 66682 559000
rect 66640 558958 66668 558991
rect 66628 558952 66680 558958
rect 66628 558894 66680 558900
rect 66350 555248 66406 555257
rect 66350 555183 66406 555192
rect 66364 554810 66392 555183
rect 66352 554804 66404 554810
rect 66352 554746 66404 554752
rect 66260 554736 66312 554742
rect 66258 554704 66260 554713
rect 66312 554704 66314 554713
rect 66258 554639 66314 554648
rect 66534 549672 66590 549681
rect 66534 549607 66590 549616
rect 66548 549302 66576 549607
rect 66536 549296 66588 549302
rect 66536 549238 66588 549244
rect 66534 548312 66590 548321
rect 66534 548247 66590 548256
rect 66548 547942 66576 548247
rect 66536 547936 66588 547942
rect 66536 547878 66588 547884
rect 66812 547800 66864 547806
rect 66812 547742 66864 547748
rect 66824 547641 66852 547742
rect 66810 547632 66866 547641
rect 66810 547567 66866 547576
rect 66166 546408 66222 546417
rect 66166 546343 66222 546352
rect 66180 545766 66208 546343
rect 66168 545760 66220 545766
rect 66168 545702 66220 545708
rect 66812 545080 66864 545086
rect 66812 545022 66864 545028
rect 66824 544921 66852 545022
rect 66810 544912 66866 544921
rect 66810 544847 66866 544856
rect 66810 542736 66866 542745
rect 66810 542671 66866 542680
rect 66824 542434 66852 542671
rect 66812 542428 66864 542434
rect 66812 542370 66864 542376
rect 67086 541784 67142 541793
rect 67086 541719 67142 541728
rect 67100 541686 67128 541719
rect 67088 541680 67140 541686
rect 67088 541622 67140 541628
rect 67100 539510 67128 541622
rect 67088 539504 67140 539510
rect 67088 539446 67140 539452
rect 66168 536172 66220 536178
rect 66168 536114 66220 536120
rect 66076 532024 66128 532030
rect 66076 531966 66128 531972
rect 65982 447808 66038 447817
rect 65982 447743 66038 447752
rect 65524 415200 65576 415206
rect 65524 415142 65576 415148
rect 65536 414730 65564 415142
rect 65524 414724 65576 414730
rect 65524 414666 65576 414672
rect 65892 408468 65944 408474
rect 65892 408410 65944 408416
rect 64788 405816 64840 405822
rect 64788 405758 64840 405764
rect 64696 388476 64748 388482
rect 64696 388418 64748 388424
rect 64602 387696 64658 387705
rect 64602 387631 64658 387640
rect 64800 378894 64828 405758
rect 65904 390969 65932 408410
rect 65890 390960 65946 390969
rect 65890 390895 65946 390904
rect 65996 385014 66024 447743
rect 66076 424380 66128 424386
rect 66076 424322 66128 424328
rect 65984 385008 66036 385014
rect 65984 384950 66036 384956
rect 64788 378888 64840 378894
rect 64788 378830 64840 378836
rect 66088 359514 66116 424322
rect 66180 389201 66208 536114
rect 67284 442950 67312 570143
rect 67560 566817 67588 596770
rect 67546 566808 67602 566817
rect 67546 566743 67602 566752
rect 67560 566506 67588 566743
rect 67548 566500 67600 566506
rect 67548 566442 67600 566448
rect 67652 558929 67680 703462
rect 71044 702840 71096 702846
rect 71044 702782 71096 702788
rect 69020 592680 69072 592686
rect 69020 592622 69072 592628
rect 67730 589928 67786 589937
rect 67730 589863 67786 589872
rect 67744 585857 67772 589863
rect 69032 588962 69060 592622
rect 71056 592034 71084 702782
rect 72988 699553 73016 703520
rect 73068 703316 73120 703322
rect 73068 703258 73120 703264
rect 72974 699544 73030 699553
rect 72974 699479 73030 699488
rect 70872 592006 71084 592034
rect 73080 592034 73108 703258
rect 75736 592136 75788 592142
rect 75736 592078 75788 592084
rect 73080 592006 73200 592034
rect 70872 590714 70900 592006
rect 72422 590880 72478 590889
rect 72422 590815 72478 590824
rect 70860 590708 70912 590714
rect 70860 590650 70912 590656
rect 71688 590708 71740 590714
rect 71688 590650 71740 590656
rect 70308 589416 70360 589422
rect 70308 589358 70360 589364
rect 70320 589098 70348 589358
rect 70104 589070 70348 589098
rect 70872 589098 70900 590650
rect 71700 589966 71728 590650
rect 71688 589960 71740 589966
rect 71688 589902 71740 589908
rect 72436 589098 72464 590815
rect 73172 590073 73200 592006
rect 73618 590744 73674 590753
rect 75748 590714 75776 592078
rect 73618 590679 73674 590688
rect 75000 590708 75052 590714
rect 73158 590064 73214 590073
rect 73158 589999 73214 590008
rect 73172 589098 73200 589999
rect 70872 589070 71208 589098
rect 72128 589070 72464 589098
rect 73048 589070 73200 589098
rect 73632 589098 73660 590679
rect 75000 590650 75052 590656
rect 75736 590708 75788 590714
rect 75736 590650 75788 590656
rect 73632 589070 73968 589098
rect 75012 588962 75040 590650
rect 75840 589404 75868 703530
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 89180 700398 89208 703520
rect 93768 703452 93820 703458
rect 93768 703394 93820 703400
rect 89812 702636 89864 702642
rect 89812 702578 89864 702584
rect 83464 700392 83516 700398
rect 83464 700334 83516 700340
rect 89168 700392 89220 700398
rect 89168 700334 89220 700340
rect 79968 597576 80020 597582
rect 79968 597518 80020 597524
rect 79980 596154 80008 597518
rect 83476 596174 83504 700334
rect 89076 700324 89128 700330
rect 89076 700266 89128 700272
rect 87604 605872 87656 605878
rect 87604 605814 87656 605820
rect 79968 596148 80020 596154
rect 83476 596146 83780 596174
rect 79968 596090 80020 596096
rect 77024 594856 77076 594862
rect 77024 594798 77076 594804
rect 75794 589376 75868 589404
rect 75794 588962 75822 589376
rect 77036 589098 77064 594798
rect 77942 592104 77998 592113
rect 77942 592039 77998 592048
rect 79784 592068 79836 592074
rect 77956 589098 77984 592039
rect 79784 592010 79836 592016
rect 78404 590844 78456 590850
rect 78404 590786 78456 590792
rect 76728 589070 77064 589098
rect 77648 589070 77984 589098
rect 69032 588934 69520 588962
rect 74888 588934 75040 588962
rect 75656 588948 75822 588962
rect 75656 588934 75808 588948
rect 69492 588674 69520 588934
rect 75656 588849 75684 588934
rect 75642 588840 75698 588849
rect 78416 588826 78444 590786
rect 79796 589098 79824 592010
rect 79980 591954 80008 596090
rect 83464 593428 83516 593434
rect 83464 593370 83516 593376
rect 79980 591926 80100 591954
rect 79488 589070 79824 589098
rect 80072 589098 80100 591926
rect 82542 591016 82598 591025
rect 82542 590951 82598 590960
rect 81348 589484 81400 589490
rect 81348 589426 81400 589432
rect 81360 589274 81388 589426
rect 81314 589246 81388 589274
rect 80072 589070 80408 589098
rect 81314 589084 81342 589246
rect 82556 589098 82584 590951
rect 83476 589098 83504 593370
rect 83752 591977 83780 596146
rect 87616 594590 87644 605814
rect 87604 594584 87656 594590
rect 87604 594526 87656 594532
rect 83738 591968 83794 591977
rect 83738 591903 83794 591912
rect 86866 590880 86922 590889
rect 86866 590815 86922 590824
rect 84106 590744 84162 590753
rect 84106 590679 84162 590688
rect 84120 589404 84148 590679
rect 82248 589070 82584 589098
rect 83168 589070 83504 589098
rect 84074 589376 84148 589404
rect 84074 589084 84102 589376
rect 86880 589274 86908 590815
rect 86834 589246 86908 589274
rect 86834 589084 86862 589246
rect 78416 588798 78568 588826
rect 75642 588775 75698 588784
rect 84382 588704 84438 588713
rect 69480 588668 69532 588674
rect 87878 588704 87934 588713
rect 87768 588662 87878 588690
rect 84382 588639 84438 588648
rect 87878 588639 87934 588648
rect 88984 588668 89036 588674
rect 69480 588610 69532 588616
rect 84396 588470 84424 588639
rect 88984 588610 89036 588616
rect 85580 588600 85632 588606
rect 85008 588548 85580 588554
rect 85008 588542 85632 588548
rect 85008 588526 85620 588542
rect 85928 588526 86264 588554
rect 86236 588470 86264 588526
rect 84384 588464 84436 588470
rect 84384 588406 84436 588412
rect 86224 588464 86276 588470
rect 88890 588432 88946 588441
rect 86224 588406 86276 588412
rect 88688 588390 88890 588418
rect 88890 588367 88946 588376
rect 67730 585848 67786 585857
rect 67730 585783 67786 585792
rect 67744 585206 67772 585783
rect 67732 585200 67784 585206
rect 67732 585142 67784 585148
rect 67730 583808 67786 583817
rect 67730 583743 67786 583752
rect 67638 558920 67694 558929
rect 67638 558855 67694 558864
rect 67652 557598 67680 558855
rect 67640 557592 67692 557598
rect 67640 557534 67692 557540
rect 67362 556336 67418 556345
rect 67362 556271 67418 556280
rect 67272 442944 67324 442950
rect 67272 442886 67324 442892
rect 66994 439920 67050 439929
rect 66994 439855 67050 439864
rect 67008 439074 67036 439855
rect 66996 439068 67048 439074
rect 66996 439010 67048 439016
rect 67272 439068 67324 439074
rect 67272 439010 67324 439016
rect 66810 437744 66866 437753
rect 66810 437679 66866 437688
rect 66824 437510 66852 437679
rect 66812 437504 66864 437510
rect 66812 437446 66864 437452
rect 66812 435396 66864 435402
rect 66812 435338 66864 435344
rect 66824 435305 66852 435338
rect 66810 435296 66866 435305
rect 66810 435231 66866 435240
rect 66902 433120 66958 433129
rect 66902 433055 66958 433064
rect 66916 432070 66944 433055
rect 66904 432064 66956 432070
rect 66904 432006 66956 432012
rect 66904 431928 66956 431934
rect 66904 431870 66956 431876
rect 66916 430953 66944 431870
rect 66902 430944 66958 430953
rect 66902 430879 66958 430888
rect 66812 429140 66864 429146
rect 66812 429082 66864 429088
rect 66824 428505 66852 429082
rect 66810 428496 66866 428505
rect 66810 428431 66866 428440
rect 66258 426320 66314 426329
rect 66258 426255 66314 426264
rect 66272 425134 66300 426255
rect 66260 425128 66312 425134
rect 66260 425070 66312 425076
rect 66260 424380 66312 424386
rect 66260 424322 66312 424328
rect 66272 424153 66300 424322
rect 66258 424144 66314 424153
rect 66258 424079 66314 424088
rect 66258 421968 66314 421977
rect 66258 421903 66314 421912
rect 66272 421598 66300 421903
rect 66260 421592 66312 421598
rect 66260 421534 66312 421540
rect 66902 417344 66958 417353
rect 66902 417279 66958 417288
rect 66916 416838 66944 417279
rect 66904 416832 66956 416838
rect 66904 416774 66956 416780
rect 66444 415200 66496 415206
rect 66442 415168 66444 415177
rect 66496 415168 66498 415177
rect 66442 415103 66498 415112
rect 66536 408468 66588 408474
rect 66536 408410 66588 408416
rect 66548 408377 66576 408410
rect 66534 408368 66590 408377
rect 66534 408303 66590 408312
rect 66626 406192 66682 406201
rect 66626 406127 66682 406136
rect 66640 405822 66668 406127
rect 66628 405816 66680 405822
rect 66628 405758 66680 405764
rect 66350 403744 66406 403753
rect 66350 403679 66406 403688
rect 66364 403646 66392 403679
rect 66352 403640 66404 403646
rect 66352 403582 66404 403588
rect 66812 401600 66864 401606
rect 66810 401568 66812 401577
rect 66864 401568 66866 401577
rect 66810 401503 66866 401512
rect 66352 399492 66404 399498
rect 66352 399434 66404 399440
rect 66364 399401 66392 399434
rect 66350 399392 66406 399401
rect 66350 399327 66406 399336
rect 66994 396944 67050 396953
rect 66994 396879 67050 396888
rect 67008 396778 67036 396879
rect 66996 396772 67048 396778
rect 66996 396714 67048 396720
rect 66260 393304 66312 393310
rect 66260 393246 66312 393252
rect 66272 392601 66300 393246
rect 66258 392592 66314 392601
rect 66258 392527 66314 392536
rect 66166 389192 66222 389201
rect 66166 389127 66222 389136
rect 66076 359508 66128 359514
rect 66076 359450 66128 359456
rect 64788 356720 64840 356726
rect 64788 356662 64840 356668
rect 64696 339516 64748 339522
rect 64696 339458 64748 339464
rect 64602 332888 64658 332897
rect 64602 332823 64658 332832
rect 64616 300830 64644 332823
rect 64708 302190 64736 339458
rect 64696 302184 64748 302190
rect 64696 302126 64748 302132
rect 64604 300824 64656 300830
rect 64604 300766 64656 300772
rect 64696 296744 64748 296750
rect 64696 296686 64748 296692
rect 63316 289944 63368 289950
rect 63316 289886 63368 289892
rect 63224 280220 63276 280226
rect 63224 280162 63276 280168
rect 62028 273284 62080 273290
rect 62028 273226 62080 273232
rect 61934 199336 61990 199345
rect 61934 199271 61990 199280
rect 60646 71088 60702 71097
rect 60646 71023 60702 71032
rect 61936 33856 61988 33862
rect 61936 33798 61988 33804
rect 59266 22672 59322 22681
rect 59266 22607 59322 22616
rect 61948 16574 61976 33798
rect 62040 29646 62068 273226
rect 63132 271924 63184 271930
rect 63132 271866 63184 271872
rect 63144 230450 63172 271866
rect 63236 233918 63264 280162
rect 63224 233912 63276 233918
rect 63224 233854 63276 233860
rect 63132 230444 63184 230450
rect 63132 230386 63184 230392
rect 63328 201482 63356 289886
rect 64512 269136 64564 269142
rect 64512 269078 64564 269084
rect 63500 261520 63552 261526
rect 63500 261462 63552 261468
rect 63512 260982 63540 261462
rect 63500 260976 63552 260982
rect 63500 260918 63552 260924
rect 63408 242956 63460 242962
rect 63408 242898 63460 242904
rect 63316 201476 63368 201482
rect 63316 201418 63368 201424
rect 63420 65521 63448 242898
rect 64524 242214 64552 269078
rect 64604 255332 64656 255338
rect 64604 255274 64656 255280
rect 64512 242208 64564 242214
rect 64512 242150 64564 242156
rect 64616 224913 64644 255274
rect 64602 224904 64658 224913
rect 64602 224839 64658 224848
rect 64708 217297 64736 296686
rect 64800 266558 64828 356662
rect 65982 346352 66038 346361
rect 65982 346287 66038 346296
rect 65892 327752 65944 327758
rect 65892 327694 65944 327700
rect 65904 307766 65932 327694
rect 65996 320249 66024 346287
rect 67284 345014 67312 439010
rect 67376 419529 67404 556271
rect 67454 552256 67510 552265
rect 67454 552191 67510 552200
rect 67362 419520 67418 419529
rect 67362 419455 67418 419464
rect 67468 412729 67496 552191
rect 67548 540932 67600 540938
rect 67548 540874 67600 540880
rect 67560 539646 67588 540874
rect 67548 539640 67600 539646
rect 67548 539582 67600 539588
rect 67548 539504 67600 539510
rect 67548 539446 67600 539452
rect 67454 412720 67510 412729
rect 67454 412655 67510 412664
rect 67362 396944 67418 396953
rect 67362 396879 67418 396888
rect 67376 347721 67404 396879
rect 67362 347712 67418 347721
rect 67362 347647 67418 347656
rect 67192 344986 67312 345014
rect 67192 341193 67220 344986
rect 67178 341184 67234 341193
rect 67178 341119 67234 341128
rect 66074 336968 66130 336977
rect 66074 336903 66130 336912
rect 65982 320240 66038 320249
rect 65982 320175 66038 320184
rect 65892 307760 65944 307766
rect 65892 307702 65944 307708
rect 65522 304736 65578 304745
rect 65522 304671 65578 304680
rect 65536 284986 65564 304671
rect 66088 302569 66116 336903
rect 66168 333396 66220 333402
rect 66168 333338 66220 333344
rect 66074 302560 66130 302569
rect 66074 302495 66130 302504
rect 65524 284980 65576 284986
rect 65524 284922 65576 284928
rect 66180 276185 66208 333338
rect 67192 328409 67220 341119
rect 67272 336796 67324 336802
rect 67272 336738 67324 336744
rect 67178 328400 67234 328409
rect 67178 328335 67234 328344
rect 66810 324864 66866 324873
rect 66810 324799 66866 324808
rect 66824 324358 66852 324799
rect 66812 324352 66864 324358
rect 66812 324294 66864 324300
rect 66810 323776 66866 323785
rect 66810 323711 66866 323720
rect 66824 322998 66852 323711
rect 66812 322992 66864 322998
rect 66812 322934 66864 322940
rect 67284 322697 67312 336738
rect 67364 327820 67416 327826
rect 67364 327762 67416 327768
rect 67270 322688 67326 322697
rect 67270 322623 67326 322632
rect 66258 319424 66314 319433
rect 66258 319359 66314 319368
rect 66272 318850 66300 319359
rect 66260 318844 66312 318850
rect 67376 318794 67404 327762
rect 66260 318786 66312 318792
rect 67284 318766 67404 318794
rect 66350 318336 66406 318345
rect 66350 318271 66406 318280
rect 66260 317552 66312 317558
rect 66258 317520 66260 317529
rect 66312 317520 66314 317529
rect 66364 317490 66392 318271
rect 66258 317455 66314 317464
rect 66352 317484 66404 317490
rect 66352 317426 66404 317432
rect 66996 315988 67048 315994
rect 66996 315930 67048 315936
rect 66442 315344 66498 315353
rect 66442 315279 66498 315288
rect 66456 314702 66484 315279
rect 66444 314696 66496 314702
rect 66444 314638 66496 314644
rect 66258 314256 66314 314265
rect 66258 314191 66260 314200
rect 66312 314191 66314 314200
rect 66260 314162 66312 314168
rect 66260 313268 66312 313274
rect 66260 313210 66312 313216
rect 66272 312089 66300 313210
rect 66258 312080 66314 312089
rect 66258 312015 66314 312024
rect 66812 311840 66864 311846
rect 66812 311782 66864 311788
rect 66824 311001 66852 311782
rect 66810 310992 66866 311001
rect 66810 310927 66866 310936
rect 66626 309904 66682 309913
rect 66626 309839 66682 309848
rect 66640 309194 66668 309839
rect 66628 309188 66680 309194
rect 66628 309130 66680 309136
rect 66812 302184 66864 302190
rect 66812 302126 66864 302132
rect 66824 301481 66852 302126
rect 66810 301472 66866 301481
rect 66810 301407 66866 301416
rect 66812 300824 66864 300830
rect 66812 300766 66864 300772
rect 66442 300656 66498 300665
rect 66442 300591 66498 300600
rect 66456 299538 66484 300591
rect 66824 299577 66852 300766
rect 66810 299568 66866 299577
rect 66444 299532 66496 299538
rect 66810 299503 66866 299512
rect 66444 299474 66496 299480
rect 66626 297392 66682 297401
rect 66626 297327 66682 297336
rect 66640 296750 66668 297327
rect 66628 296744 66680 296750
rect 67008 296714 67036 315930
rect 67088 309460 67140 309466
rect 67088 309402 67140 309408
rect 67100 309097 67128 309402
rect 67284 309134 67312 318766
rect 67468 309466 67496 412655
rect 67560 394777 67588 539446
rect 67744 454034 67772 583743
rect 67822 577008 67878 577017
rect 67822 576943 67878 576952
rect 67836 538966 67864 576943
rect 68652 540932 68704 540938
rect 68652 540874 68704 540880
rect 68664 540841 68692 540874
rect 68650 540832 68706 540841
rect 68650 540767 68706 540776
rect 69848 539640 69900 539646
rect 69848 539582 69900 539588
rect 69860 539458 69888 539582
rect 69736 539444 69888 539458
rect 69722 539430 69888 539444
rect 68480 539158 68816 539186
rect 67824 538960 67876 538966
rect 67824 538902 67876 538908
rect 68480 535537 68508 539158
rect 69722 539050 69750 539430
rect 70656 539158 70716 539186
rect 69676 539022 69750 539050
rect 69676 535537 69704 539022
rect 70688 538218 70716 539158
rect 71240 539158 71576 539186
rect 72436 539158 72496 539186
rect 73172 539158 73416 539186
rect 74000 539158 74336 539186
rect 74644 539158 75256 539186
rect 76024 539158 76176 539186
rect 76760 539158 77096 539186
rect 77312 539158 78016 539186
rect 78784 539158 78936 539186
rect 79520 539158 79856 539186
rect 80776 539158 80836 539186
rect 70676 538212 70728 538218
rect 70676 538154 70728 538160
rect 70688 535537 70716 538154
rect 68466 535528 68522 535537
rect 68466 535463 68522 535472
rect 69662 535528 69718 535537
rect 69662 535463 69718 535472
rect 70674 535528 70730 535537
rect 70674 535463 70730 535472
rect 71240 528554 71268 539158
rect 72436 537538 72464 539158
rect 72424 537532 72476 537538
rect 72424 537474 72476 537480
rect 70504 528526 71268 528554
rect 70504 458930 70532 528526
rect 70492 458924 70544 458930
rect 70492 458866 70544 458872
rect 72056 454776 72108 454782
rect 72056 454718 72108 454724
rect 71044 454708 71096 454714
rect 71044 454650 71096 454656
rect 67732 454028 67784 454034
rect 67732 453970 67784 453976
rect 68284 454028 68336 454034
rect 68284 453970 68336 453976
rect 68296 452742 68324 453970
rect 68744 453348 68796 453354
rect 68744 453290 68796 453296
rect 68284 452736 68336 452742
rect 68284 452678 68336 452684
rect 67732 442944 67784 442950
rect 67732 442886 67784 442892
rect 67744 442105 67772 442886
rect 67730 442096 67786 442105
rect 67730 442031 67786 442040
rect 67546 394768 67602 394777
rect 67546 394703 67602 394712
rect 67560 330177 67588 394703
rect 67638 380216 67694 380225
rect 67638 380151 67694 380160
rect 67546 330168 67602 330177
rect 67546 330103 67602 330112
rect 67456 309460 67508 309466
rect 67456 309402 67508 309408
rect 67284 309106 67404 309134
rect 67086 309088 67142 309097
rect 67086 309023 67142 309032
rect 67100 308446 67128 309023
rect 67088 308440 67140 308446
rect 67088 308382 67140 308388
rect 67178 308000 67234 308009
rect 67178 307935 67234 307944
rect 67088 307760 67140 307766
rect 67088 307702 67140 307708
rect 66628 296686 66680 296692
rect 66732 296686 67036 296714
rect 66444 296676 66496 296682
rect 66444 296618 66496 296624
rect 66456 296313 66484 296618
rect 66442 296304 66498 296313
rect 66442 296239 66498 296248
rect 66732 288969 66760 296686
rect 66810 294128 66866 294137
rect 66810 294063 66812 294072
rect 66864 294063 66866 294072
rect 66812 294034 66864 294040
rect 66812 293956 66864 293962
rect 66812 293898 66864 293904
rect 66824 291145 66852 293898
rect 66994 293040 67050 293049
rect 66994 292975 67050 292984
rect 66904 292528 66956 292534
rect 66904 292470 66956 292476
rect 66916 292233 66944 292470
rect 66902 292224 66958 292233
rect 66902 292159 66958 292168
rect 66810 291136 66866 291145
rect 66810 291071 66866 291080
rect 66810 290048 66866 290057
rect 66810 289983 66866 289992
rect 66824 289950 66852 289983
rect 66812 289944 66864 289950
rect 66812 289886 66864 289892
rect 66718 288960 66774 288969
rect 66718 288895 66774 288904
rect 66626 287872 66682 287881
rect 66626 287807 66682 287816
rect 66640 287094 66668 287807
rect 66628 287088 66680 287094
rect 67008 287054 67036 292975
rect 66628 287030 66680 287036
rect 66916 287026 67036 287054
rect 66810 286784 66866 286793
rect 66810 286719 66866 286728
rect 66824 285734 66852 286719
rect 66812 285728 66864 285734
rect 66812 285670 66864 285676
rect 66810 281616 66866 281625
rect 66810 281551 66812 281560
rect 66864 281551 66866 281560
rect 66812 281522 66864 281528
rect 66810 280528 66866 280537
rect 66810 280463 66866 280472
rect 66824 280226 66852 280463
rect 66812 280220 66864 280226
rect 66812 280162 66864 280168
rect 66442 278352 66498 278361
rect 66442 278287 66498 278296
rect 66456 277438 66484 278287
rect 66444 277432 66496 277438
rect 66444 277374 66496 277380
rect 66810 277264 66866 277273
rect 66810 277199 66866 277208
rect 66166 276176 66222 276185
rect 66166 276111 66222 276120
rect 66824 276078 66852 277199
rect 66812 276072 66864 276078
rect 66812 276014 66864 276020
rect 66810 275360 66866 275369
rect 66810 275295 66866 275304
rect 66824 274718 66852 275295
rect 66812 274712 66864 274718
rect 66812 274654 66864 274660
rect 66810 274272 66866 274281
rect 66810 274207 66866 274216
rect 66824 273290 66852 274207
rect 66812 273284 66864 273290
rect 66812 273226 66864 273232
rect 66810 273184 66866 273193
rect 66810 273119 66866 273128
rect 65890 272096 65946 272105
rect 65890 272031 65946 272040
rect 64788 266552 64840 266558
rect 64788 266494 64840 266500
rect 64788 260976 64840 260982
rect 64788 260918 64840 260924
rect 64800 229090 64828 260918
rect 65904 243409 65932 272031
rect 66824 271930 66852 273119
rect 66812 271924 66864 271930
rect 66812 271866 66864 271872
rect 66810 271008 66866 271017
rect 66810 270943 66866 270952
rect 66824 270570 66852 270943
rect 66812 270564 66864 270570
rect 66812 270506 66864 270512
rect 66810 269920 66866 269929
rect 66810 269855 66866 269864
rect 66824 269142 66852 269855
rect 66812 269136 66864 269142
rect 66812 269078 66864 269084
rect 66626 267744 66682 267753
rect 66626 267679 66682 267688
rect 66640 266558 66668 267679
rect 66168 266552 66220 266558
rect 66168 266494 66220 266500
rect 66628 266552 66680 266558
rect 66628 266494 66680 266500
rect 65982 257408 66038 257417
rect 65982 257343 66038 257352
rect 65890 243400 65946 243409
rect 65890 243335 65946 243344
rect 65996 240786 66024 257343
rect 66076 244928 66128 244934
rect 66076 244870 66128 244876
rect 65984 240780 66036 240786
rect 65984 240722 66036 240728
rect 66088 230489 66116 244870
rect 66180 235929 66208 266494
rect 66810 265840 66866 265849
rect 66810 265775 66866 265784
rect 66824 264994 66852 265775
rect 66812 264988 66864 264994
rect 66812 264930 66864 264936
rect 66718 264752 66774 264761
rect 66718 264687 66774 264696
rect 66732 263634 66760 264687
rect 66812 264240 66864 264246
rect 66812 264182 66864 264188
rect 66824 263673 66852 264182
rect 66810 263664 66866 263673
rect 66720 263628 66772 263634
rect 66810 263599 66866 263608
rect 66720 263570 66772 263576
rect 66812 262880 66864 262886
rect 66812 262822 66864 262828
rect 66824 262585 66852 262822
rect 66810 262576 66866 262585
rect 66810 262511 66866 262520
rect 66810 261488 66866 261497
rect 66810 261423 66866 261432
rect 66824 260982 66852 261423
rect 66812 260976 66864 260982
rect 66812 260918 66864 260924
rect 66260 258120 66312 258126
rect 66258 258088 66260 258097
rect 66312 258088 66314 258097
rect 66258 258023 66314 258032
rect 66810 256320 66866 256329
rect 66810 256255 66866 256264
rect 66824 255338 66852 256255
rect 66812 255332 66864 255338
rect 66812 255274 66864 255280
rect 66810 254144 66866 254153
rect 66810 254079 66866 254088
rect 66824 253978 66852 254079
rect 66812 253972 66864 253978
rect 66812 253914 66864 253920
rect 66916 253230 66944 287026
rect 66994 285696 67050 285705
rect 66994 285631 67050 285640
rect 67008 268394 67036 285631
rect 67100 284617 67128 307702
rect 67192 307086 67220 307935
rect 67180 307080 67232 307086
rect 67180 307022 67232 307028
rect 67376 305833 67404 309106
rect 67362 305824 67418 305833
rect 67362 305759 67418 305768
rect 67560 298489 67588 330103
rect 67546 298480 67602 298489
rect 67546 298415 67602 298424
rect 67546 295216 67602 295225
rect 67546 295151 67602 295160
rect 67560 294030 67588 295151
rect 67548 294024 67600 294030
rect 67548 293966 67600 293972
rect 67086 284608 67142 284617
rect 67086 284543 67142 284552
rect 67546 282704 67602 282713
rect 67546 282639 67602 282648
rect 67178 279440 67234 279449
rect 67178 279375 67234 279384
rect 67192 278798 67220 279375
rect 67180 278792 67232 278798
rect 67180 278734 67232 278740
rect 67364 269068 67416 269074
rect 67364 269010 67416 269016
rect 66996 268388 67048 268394
rect 66996 268330 67048 268336
rect 66904 253224 66956 253230
rect 66904 253166 66956 253172
rect 66810 253056 66866 253065
rect 66810 252991 66866 253000
rect 66824 252618 66852 252991
rect 66812 252612 66864 252618
rect 66812 252554 66864 252560
rect 66442 250064 66498 250073
rect 66442 249999 66498 250008
rect 66456 249830 66484 249999
rect 66444 249824 66496 249830
rect 66444 249766 66496 249772
rect 66810 247888 66866 247897
rect 66810 247823 66866 247832
rect 66824 247110 66852 247823
rect 66812 247104 66864 247110
rect 66812 247046 66864 247052
rect 67270 246800 67326 246809
rect 67270 246735 67326 246744
rect 66628 244928 66680 244934
rect 66628 244870 66680 244876
rect 66640 244633 66668 244870
rect 66626 244624 66682 244633
rect 66626 244559 66682 244568
rect 66810 243536 66866 243545
rect 66810 243471 66866 243480
rect 66824 242962 66852 243471
rect 66812 242956 66864 242962
rect 66812 242898 66864 242904
rect 67086 242856 67142 242865
rect 67086 242791 67142 242800
rect 66166 235920 66222 235929
rect 66166 235855 66222 235864
rect 66074 230480 66130 230489
rect 66074 230415 66130 230424
rect 64788 229084 64840 229090
rect 64788 229026 64840 229032
rect 64694 217288 64750 217297
rect 64694 217223 64750 217232
rect 67100 200705 67128 242791
rect 67284 215937 67312 246735
rect 67376 236609 67404 269010
rect 67454 255232 67510 255241
rect 67454 255167 67510 255176
rect 67468 241777 67496 255167
rect 67454 241768 67510 241777
rect 67454 241703 67510 241712
rect 67560 240106 67588 282639
rect 67652 269074 67680 380151
rect 67744 374678 67772 442031
rect 68296 440910 68324 452678
rect 68468 447840 68520 447846
rect 68468 447782 68520 447788
rect 68480 447234 68508 447782
rect 68468 447228 68520 447234
rect 68468 447170 68520 447176
rect 68652 447228 68704 447234
rect 68652 447170 68704 447176
rect 68284 440904 68336 440910
rect 68284 440846 68336 440852
rect 68664 391241 68692 447170
rect 68756 444825 68784 453290
rect 71056 449954 71084 454650
rect 72068 452674 72096 454718
rect 72056 452668 72108 452674
rect 72056 452610 72108 452616
rect 71044 449948 71096 449954
rect 71044 449890 71096 449896
rect 70306 449168 70362 449177
rect 70306 449103 70362 449112
rect 68742 444816 68798 444825
rect 68742 444751 68798 444760
rect 68756 444666 68784 444751
rect 68756 444638 68830 444666
rect 68802 444380 68830 444638
rect 70320 444530 70348 449103
rect 70274 444502 70348 444530
rect 70274 444380 70302 444502
rect 72068 444394 72096 452610
rect 72436 451994 72464 537474
rect 73172 536110 73200 539158
rect 73160 536104 73212 536110
rect 73160 536046 73212 536052
rect 74000 535498 74028 539158
rect 73160 535492 73212 535498
rect 73160 535434 73212 535440
rect 73988 535492 74040 535498
rect 73988 535434 74040 535440
rect 73172 457570 73200 535434
rect 73160 457564 73212 457570
rect 73160 457506 73212 457512
rect 72424 451988 72476 451994
rect 72424 451930 72476 451936
rect 73252 449948 73304 449954
rect 73252 449890 73304 449896
rect 73264 444666 73292 449890
rect 74644 449274 74672 539158
rect 74724 538960 74776 538966
rect 74724 538902 74776 538908
rect 74632 449268 74684 449274
rect 74632 449210 74684 449216
rect 74736 447166 74764 538902
rect 76024 536790 76052 539158
rect 76760 538121 76788 539158
rect 76746 538112 76802 538121
rect 76746 538047 76802 538056
rect 76012 536784 76064 536790
rect 76012 536726 76064 536732
rect 76024 536178 76052 536726
rect 76012 536172 76064 536178
rect 76012 536114 76064 536120
rect 76760 535537 76788 538047
rect 75918 535528 75974 535537
rect 75918 535463 75974 535472
rect 76746 535528 76802 535537
rect 76746 535463 76802 535472
rect 75932 463010 75960 535463
rect 77312 468518 77340 539158
rect 78680 533452 78732 533458
rect 78680 533394 78732 533400
rect 77944 532024 77996 532030
rect 77944 531966 77996 531972
rect 77300 468512 77352 468518
rect 77300 468454 77352 468460
rect 76562 467800 76618 467809
rect 76562 467735 76618 467744
rect 75920 463004 75972 463010
rect 75920 462946 75972 462952
rect 74724 447160 74776 447166
rect 74724 447102 74776 447108
rect 71760 444366 72096 444394
rect 73218 444638 73292 444666
rect 73218 444380 73246 444638
rect 74736 444394 74764 447102
rect 76576 445806 76604 467735
rect 77956 458250 77984 531966
rect 78692 461650 78720 533394
rect 78680 461644 78732 461650
rect 78680 461586 78732 461592
rect 78680 460216 78732 460222
rect 78680 460158 78732 460164
rect 77300 458244 77352 458250
rect 77300 458186 77352 458192
rect 77944 458244 77996 458250
rect 77944 458186 77996 458192
rect 76564 445800 76616 445806
rect 76564 445742 76616 445748
rect 76576 444394 76604 445742
rect 74736 444366 74888 444394
rect 76360 444366 76604 444394
rect 77312 444394 77340 458186
rect 78692 446962 78720 460158
rect 78784 447817 78812 539158
rect 79520 533458 79548 539158
rect 80808 538286 80836 539158
rect 81452 539158 81696 539186
rect 82616 539158 82768 539186
rect 83536 539158 84148 539186
rect 84456 539158 84792 539186
rect 85376 539158 85528 539186
rect 86296 539158 86632 539186
rect 80336 538280 80388 538286
rect 80336 538222 80388 538228
rect 80796 538280 80848 538286
rect 80796 538222 80848 538228
rect 79508 533452 79560 533458
rect 79508 533394 79560 533400
rect 80348 528554 80376 538222
rect 80072 528526 80376 528554
rect 80072 464370 80100 528526
rect 80060 464364 80112 464370
rect 80060 464306 80112 464312
rect 81452 462913 81480 539158
rect 82740 536761 82768 539158
rect 82726 536752 82782 536761
rect 82726 536687 82782 536696
rect 81438 462904 81494 462913
rect 81438 462839 81494 462848
rect 82740 453257 82768 536687
rect 83464 457496 83516 457502
rect 83464 457438 83516 457444
rect 82726 453248 82782 453257
rect 82726 453183 82782 453192
rect 82084 452736 82136 452742
rect 82084 452678 82136 452684
rect 80060 449200 80112 449206
rect 80060 449142 80112 449148
rect 80072 448594 80100 449142
rect 80060 448588 80112 448594
rect 80060 448530 80112 448536
rect 80888 448588 80940 448594
rect 80888 448530 80940 448536
rect 78770 447808 78826 447817
rect 78770 447743 78826 447752
rect 78680 446956 78732 446962
rect 78680 446898 78732 446904
rect 79140 446956 79192 446962
rect 79140 446898 79192 446904
rect 79152 445874 79180 446898
rect 79140 445868 79192 445874
rect 79140 445810 79192 445816
rect 79152 444394 79180 445810
rect 80900 444530 80928 448530
rect 80900 444502 80974 444530
rect 77312 444366 77832 444394
rect 79152 444366 79488 444394
rect 80946 444380 80974 444502
rect 82096 444394 82124 452678
rect 83476 451353 83504 457438
rect 84120 454753 84148 539158
rect 84764 536081 84792 539158
rect 85500 536246 85528 539158
rect 86604 538214 86632 539158
rect 86972 539158 87400 539186
rect 88320 539158 88380 539186
rect 86868 538214 86920 538218
rect 86604 538212 86920 538214
rect 86604 538186 86868 538212
rect 86868 538154 86920 538160
rect 85488 536240 85540 536246
rect 85488 536182 85540 536188
rect 86224 536240 86276 536246
rect 86224 536182 86276 536188
rect 84750 536072 84806 536081
rect 84750 536007 84806 536016
rect 85580 458856 85632 458862
rect 85580 458798 85632 458804
rect 84106 454744 84162 454753
rect 84106 454679 84162 454688
rect 83462 451344 83518 451353
rect 83462 451279 83518 451288
rect 83476 444394 83504 451279
rect 85592 445913 85620 458798
rect 86236 447817 86264 536182
rect 86880 457473 86908 538154
rect 86972 461553 87000 539158
rect 86958 461544 87014 461553
rect 86958 461479 87014 461488
rect 86960 460964 87012 460970
rect 86960 460906 87012 460912
rect 86866 457464 86922 457473
rect 86866 457399 86922 457408
rect 86222 447808 86278 447817
rect 86222 447743 86278 447752
rect 85578 445904 85634 445913
rect 85578 445839 85634 445848
rect 85592 444666 85620 445839
rect 85546 444638 85620 444666
rect 86972 444666 87000 460906
rect 88352 456113 88380 539158
rect 88338 456104 88394 456113
rect 88338 456039 88394 456048
rect 88996 451274 89024 588610
rect 89088 575550 89116 700266
rect 89166 593464 89222 593473
rect 89166 593399 89222 593408
rect 89180 588470 89208 593399
rect 89720 589416 89772 589422
rect 89720 589358 89772 589364
rect 89168 588464 89220 588470
rect 89168 588406 89220 588412
rect 89180 585818 89208 588406
rect 89168 585812 89220 585818
rect 89168 585754 89220 585760
rect 89076 575544 89128 575550
rect 89076 575486 89128 575492
rect 88812 451246 89024 451274
rect 88812 445777 88840 451246
rect 88798 445768 88854 445777
rect 88798 445703 88854 445712
rect 86972 444638 87046 444666
rect 82096 444366 82432 444394
rect 83476 444366 83904 444394
rect 85546 444380 85574 444638
rect 87018 444380 87046 444638
rect 88812 444394 88840 445703
rect 88504 444366 88840 444394
rect 89732 444394 89760 589358
rect 89824 560153 89852 702578
rect 91192 594584 91244 594590
rect 91192 594526 91244 594532
rect 89902 585712 89958 585721
rect 89902 585647 89958 585656
rect 89810 560144 89866 560153
rect 89810 560079 89866 560088
rect 89916 538898 89944 585647
rect 91098 581632 91154 581641
rect 91098 581567 91154 581576
rect 91112 581058 91140 581567
rect 91100 581052 91152 581058
rect 91100 580994 91152 581000
rect 91098 578912 91154 578921
rect 91098 578847 91154 578856
rect 91112 578270 91140 578847
rect 91100 578264 91152 578270
rect 91100 578206 91152 578212
rect 91098 577552 91154 577561
rect 91098 577487 91154 577496
rect 91112 576910 91140 577487
rect 91100 576904 91152 576910
rect 91100 576846 91152 576852
rect 91204 576745 91232 594526
rect 92480 587852 92532 587858
rect 92480 587794 92532 587800
rect 91926 584624 91982 584633
rect 91926 584559 91982 584568
rect 91940 584458 91968 584559
rect 91928 584452 91980 584458
rect 91928 584394 91980 584400
rect 91928 583704 91980 583710
rect 91926 583672 91928 583681
rect 91980 583672 91982 583681
rect 91926 583607 91982 583616
rect 91190 576736 91246 576745
rect 91190 576671 91246 576680
rect 91204 576162 91232 576671
rect 91192 576156 91244 576162
rect 91192 576098 91244 576104
rect 91284 575544 91336 575550
rect 91284 575486 91336 575492
rect 91098 573472 91154 573481
rect 91098 573407 91154 573416
rect 91112 572762 91140 573407
rect 91100 572756 91152 572762
rect 91100 572698 91152 572704
rect 91190 572112 91246 572121
rect 91190 572047 91246 572056
rect 91100 571464 91152 571470
rect 91098 571432 91100 571441
rect 91152 571432 91154 571441
rect 91204 571402 91232 572047
rect 91098 571367 91154 571376
rect 91192 571396 91244 571402
rect 91192 571338 91244 571344
rect 91098 570072 91154 570081
rect 91098 570007 91154 570016
rect 91112 569974 91140 570007
rect 91100 569968 91152 569974
rect 91100 569910 91152 569916
rect 91296 567905 91324 575486
rect 91926 574832 91982 574841
rect 91926 574767 91928 574776
rect 91980 574767 91982 574776
rect 91928 574738 91980 574744
rect 91742 568712 91798 568721
rect 91742 568647 91798 568656
rect 91282 567896 91338 567905
rect 91282 567831 91284 567840
rect 91336 567831 91338 567840
rect 91284 567802 91336 567808
rect 91296 567771 91324 567802
rect 91100 565888 91152 565894
rect 91098 565856 91100 565865
rect 91152 565856 91154 565865
rect 91098 565791 91154 565800
rect 91098 564496 91154 564505
rect 91098 564431 91100 564440
rect 91152 564431 91154 564440
rect 91100 564402 91152 564408
rect 91098 563136 91154 563145
rect 91098 563071 91100 563080
rect 91152 563071 91154 563080
rect 91100 563042 91152 563048
rect 91098 560960 91154 560969
rect 91098 560895 91154 560904
rect 89904 538892 89956 538898
rect 89904 538834 89956 538840
rect 91112 530602 91140 560895
rect 91190 558240 91246 558249
rect 91190 558175 91246 558184
rect 91204 557598 91232 558175
rect 91192 557592 91244 557598
rect 91192 557534 91244 557540
rect 91190 556880 91246 556889
rect 91190 556815 91246 556824
rect 91204 556238 91232 556815
rect 91192 556232 91244 556238
rect 91192 556174 91244 556180
rect 91190 555520 91246 555529
rect 91190 555455 91246 555464
rect 91204 554810 91232 555455
rect 91192 554804 91244 554810
rect 91192 554746 91244 554752
rect 91282 552800 91338 552809
rect 91282 552735 91338 552744
rect 91192 552152 91244 552158
rect 91190 552120 91192 552129
rect 91244 552120 91246 552129
rect 91296 552090 91324 552735
rect 91190 552055 91246 552064
rect 91284 552084 91336 552090
rect 91284 552026 91336 552032
rect 91190 549400 91246 549409
rect 91190 549335 91246 549344
rect 91204 549302 91232 549335
rect 91192 549296 91244 549302
rect 91192 549238 91244 549244
rect 91190 547904 91246 547913
rect 91190 547839 91246 547848
rect 91204 533390 91232 547839
rect 91282 546544 91338 546553
rect 91282 546479 91284 546488
rect 91336 546479 91338 546488
rect 91284 546450 91336 546456
rect 91296 545850 91324 546450
rect 91296 545822 91416 545850
rect 91284 545760 91336 545766
rect 91284 545702 91336 545708
rect 91296 545465 91324 545702
rect 91282 545456 91338 545465
rect 91282 545391 91338 545400
rect 91284 544400 91336 544406
rect 91284 544342 91336 544348
rect 91296 544105 91324 544342
rect 91282 544096 91338 544105
rect 91282 544031 91338 544040
rect 91282 542464 91338 542473
rect 91282 542399 91284 542408
rect 91336 542399 91338 542408
rect 91284 542370 91336 542376
rect 91284 541680 91336 541686
rect 91284 541622 91336 541628
rect 91296 541385 91324 541622
rect 91282 541376 91338 541385
rect 91282 541311 91338 541320
rect 91282 539744 91338 539753
rect 91282 539679 91284 539688
rect 91336 539679 91338 539688
rect 91284 539650 91336 539656
rect 91388 534750 91416 545822
rect 91376 534744 91428 534750
rect 91376 534686 91428 534692
rect 91192 533384 91244 533390
rect 91192 533326 91244 533332
rect 91100 530596 91152 530602
rect 91100 530538 91152 530544
rect 91100 456068 91152 456074
rect 91100 456010 91152 456016
rect 91112 454102 91140 456010
rect 91100 454096 91152 454102
rect 91100 454038 91152 454044
rect 91112 451274 91140 454038
rect 91756 453354 91784 568647
rect 91834 560144 91890 560153
rect 91834 560079 91890 560088
rect 91848 548554 91876 560079
rect 91836 548548 91888 548554
rect 91836 548490 91888 548496
rect 91744 453348 91796 453354
rect 91744 453290 91796 453296
rect 91112 451246 91232 451274
rect 90132 444544 90188 444553
rect 90132 444479 90188 444488
rect 90146 444394 90174 444479
rect 89732 444380 90174 444394
rect 91204 444394 91232 451246
rect 92492 444514 92520 587794
rect 93780 584458 93808 703394
rect 101496 703112 101548 703118
rect 101496 703054 101548 703060
rect 97908 702772 97960 702778
rect 97908 702714 97960 702720
rect 94504 702636 94556 702642
rect 94504 702578 94556 702584
rect 93768 584452 93820 584458
rect 93768 584394 93820 584400
rect 94516 583710 94544 702578
rect 96620 592136 96672 592142
rect 96620 592078 96672 592084
rect 95882 590880 95938 590889
rect 95882 590815 95938 590824
rect 93768 583704 93820 583710
rect 93768 583646 93820 583652
rect 94504 583704 94556 583710
rect 94504 583646 94556 583652
rect 93780 581641 93808 583646
rect 93766 581632 93822 581641
rect 93766 581567 93822 581576
rect 93768 574796 93820 574802
rect 93768 574738 93820 574744
rect 93780 569226 93808 574738
rect 94504 571464 94556 571470
rect 94504 571406 94556 571412
rect 93768 569220 93820 569226
rect 93768 569162 93820 569168
rect 93124 539708 93176 539714
rect 93124 539650 93176 539656
rect 93136 512689 93164 539650
rect 93122 512680 93178 512689
rect 93122 512615 93178 512624
rect 94516 463010 94544 571406
rect 95896 543046 95924 590815
rect 96436 545760 96488 545766
rect 96436 545702 96488 545708
rect 95884 543040 95936 543046
rect 95884 542982 95936 542988
rect 96448 467129 96476 545702
rect 96528 544400 96580 544406
rect 96528 544342 96580 544348
rect 96434 467120 96490 467129
rect 96434 467055 96490 467064
rect 95884 465724 95936 465730
rect 95884 465666 95936 465672
rect 94504 463004 94556 463010
rect 94504 462946 94556 462952
rect 95896 447166 95924 465666
rect 96540 464409 96568 544342
rect 96526 464400 96582 464409
rect 96526 464335 96582 464344
rect 95884 447160 95936 447166
rect 95884 447102 95936 447108
rect 94410 445768 94466 445777
rect 94410 445703 94466 445712
rect 92480 444508 92532 444514
rect 92480 444450 92532 444456
rect 93078 444508 93130 444514
rect 93078 444450 93130 444456
rect 89732 444366 90160 444380
rect 91204 444366 91632 444394
rect 93090 444380 93118 444450
rect 94424 444394 94452 445703
rect 95896 444394 95924 447102
rect 96632 445777 96660 592078
rect 97920 580961 97948 702714
rect 101404 594856 101456 594862
rect 101404 594798 101456 594804
rect 98642 592104 98698 592113
rect 98642 592039 98698 592048
rect 97906 580952 97962 580961
rect 97906 580887 97962 580896
rect 97920 580281 97948 580887
rect 97906 580272 97962 580281
rect 97906 580207 97962 580216
rect 97264 542428 97316 542434
rect 97264 542370 97316 542376
rect 97276 458153 97304 542370
rect 97262 458144 97318 458153
rect 97262 458079 97318 458088
rect 98552 456816 98604 456822
rect 98552 456758 98604 456764
rect 96618 445768 96674 445777
rect 96618 445703 96674 445712
rect 97354 445768 97410 445777
rect 97354 445703 97410 445712
rect 97368 444394 97396 445703
rect 98564 444394 98592 456758
rect 98656 445777 98684 592039
rect 98734 588704 98790 588713
rect 98734 588639 98790 588648
rect 98748 456822 98776 588639
rect 100668 577516 100720 577522
rect 100668 577458 100720 577464
rect 100680 576910 100708 577458
rect 100668 576904 100720 576910
rect 100668 576846 100720 576852
rect 98736 456816 98788 456822
rect 98736 456758 98788 456764
rect 100680 447817 100708 576846
rect 100666 447808 100722 447817
rect 100666 447743 100722 447752
rect 98642 445768 98698 445777
rect 98642 445703 98698 445712
rect 101416 444514 101444 594798
rect 101508 574802 101536 703054
rect 104912 599622 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 122104 703656 122156 703662
rect 122104 703598 122156 703604
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 104900 599616 104952 599622
rect 104900 599558 104952 599564
rect 106924 597576 106976 597582
rect 106924 597518 106976 597524
rect 105544 592068 105596 592074
rect 105544 592010 105596 592016
rect 103520 590844 103572 590850
rect 103520 590786 103572 590792
rect 102784 581052 102836 581058
rect 102784 580994 102836 581000
rect 101496 574796 101548 574802
rect 101496 574738 101548 574744
rect 101496 565888 101548 565894
rect 101496 565830 101548 565836
rect 101508 456074 101536 565830
rect 102796 512650 102824 580994
rect 102784 512644 102836 512650
rect 102784 512586 102836 512592
rect 101496 456068 101548 456074
rect 101496 456010 101548 456016
rect 103532 447234 103560 590786
rect 104256 549296 104308 549302
rect 104256 549238 104308 549244
rect 104164 546508 104216 546514
rect 104164 546450 104216 546456
rect 104176 458289 104204 546450
rect 104268 463593 104296 549238
rect 104254 463584 104310 463593
rect 104254 463519 104310 463528
rect 104162 458280 104218 458289
rect 104162 458215 104218 458224
rect 103520 447228 103572 447234
rect 103520 447170 103572 447176
rect 102138 445768 102194 445777
rect 102138 445703 102194 445712
rect 101404 444508 101456 444514
rect 101404 444450 101456 444456
rect 101416 444394 101444 444450
rect 94424 444366 94760 444394
rect 95896 444366 96232 444394
rect 97368 444366 97704 444394
rect 98564 444366 99176 444394
rect 100832 444366 101444 444394
rect 102152 444394 102180 445703
rect 103532 444394 103560 447170
rect 105556 445913 105584 592010
rect 105636 576156 105688 576162
rect 105636 576098 105688 576104
rect 105648 457502 105676 576098
rect 105636 457496 105688 457502
rect 105636 457438 105688 457444
rect 105542 445904 105598 445913
rect 106936 445874 106964 597518
rect 108304 595468 108356 595474
rect 108304 595410 108356 595416
rect 107106 591016 107162 591025
rect 107106 590951 107162 590960
rect 107120 553110 107148 590951
rect 108316 589354 108344 595410
rect 110420 593428 110472 593434
rect 110420 593370 110472 593376
rect 108304 589348 108356 589354
rect 108304 589290 108356 589296
rect 107108 553104 107160 553110
rect 107108 553046 107160 553052
rect 107016 552152 107068 552158
rect 107016 552094 107068 552100
rect 107028 461553 107056 552094
rect 107014 461544 107070 461553
rect 107014 461479 107070 461488
rect 108316 449993 108344 589290
rect 108948 554804 109000 554810
rect 108948 554746 109000 554752
rect 108302 449984 108358 449993
rect 108302 449919 108358 449928
rect 105542 445839 105598 445848
rect 106924 445868 106976 445874
rect 105556 444394 105584 445839
rect 106924 445810 106976 445816
rect 106936 444666 106964 445810
rect 102152 444366 102304 444394
rect 103532 444366 103776 444394
rect 105432 444366 105584 444394
rect 106890 444638 106964 444666
rect 108316 444666 108344 449919
rect 108960 447953 108988 554746
rect 109040 553104 109092 553110
rect 109040 553046 109092 553052
rect 108946 447944 109002 447953
rect 108946 447879 109002 447888
rect 108316 444638 108390 444666
rect 106890 444380 106918 444638
rect 108362 444380 108390 444638
rect 109052 444394 109080 553046
rect 110432 445777 110460 593370
rect 114468 588600 114520 588606
rect 114468 588542 114520 588548
rect 114480 587858 114508 588542
rect 122116 587858 122144 703598
rect 136652 703582 137692 703610
rect 130384 703248 130436 703254
rect 130384 703190 130436 703196
rect 124864 703044 124916 703050
rect 124864 702986 124916 702992
rect 114468 587852 114520 587858
rect 114468 587794 114520 587800
rect 122104 587852 122156 587858
rect 122104 587794 122156 587800
rect 112442 585440 112498 585449
rect 112442 585375 112498 585384
rect 112456 455462 112484 585375
rect 112444 455456 112496 455462
rect 112444 455398 112496 455404
rect 112456 451246 112484 455398
rect 112444 451240 112496 451246
rect 112444 451182 112496 451188
rect 110418 445768 110474 445777
rect 110418 445703 110474 445712
rect 111430 445768 111486 445777
rect 111430 445703 111486 445712
rect 109498 444680 109554 444689
rect 109498 444615 109554 444624
rect 109512 444394 109540 444615
rect 111444 444530 111472 445703
rect 111444 444502 111518 444530
rect 109052 444366 109848 444394
rect 111490 444380 111518 444502
rect 112456 444394 112484 451182
rect 114480 444825 114508 587794
rect 116584 585812 116636 585818
rect 116584 585754 116636 585760
rect 115204 584452 115256 584458
rect 115204 584394 115256 584400
rect 115216 447846 115244 584394
rect 116596 450022 116624 585754
rect 121552 578264 121604 578270
rect 121552 578206 121604 578212
rect 120724 572756 120776 572762
rect 120724 572698 120776 572704
rect 120632 564460 120684 564466
rect 120632 564402 120684 564408
rect 117320 543040 117372 543046
rect 117320 542982 117372 542988
rect 116584 450016 116636 450022
rect 116584 449958 116636 449964
rect 115204 447840 115256 447846
rect 115204 447782 115256 447788
rect 114466 444816 114522 444825
rect 114466 444751 114522 444760
rect 114480 444666 114508 444751
rect 114434 444638 114508 444666
rect 112456 444366 112976 444394
rect 114434 444380 114462 444638
rect 116596 444394 116624 449958
rect 117332 445777 117360 542982
rect 118698 460184 118754 460193
rect 118698 460119 118754 460128
rect 117318 445768 117374 445777
rect 117318 445703 117374 445712
rect 116104 444366 116624 444394
rect 117332 444394 117360 445703
rect 118712 444446 118740 460119
rect 119020 444680 119076 444689
rect 119020 444615 119076 444624
rect 118700 444440 118752 444446
rect 117332 444366 117576 444394
rect 119034 444394 119062 444615
rect 118752 444388 119062 444394
rect 118700 444382 119062 444388
rect 118712 444380 119062 444382
rect 118712 444366 119048 444380
rect 120644 404297 120672 564402
rect 120736 418985 120764 572698
rect 121460 548548 121512 548554
rect 121460 548490 121512 548496
rect 120816 451920 120868 451926
rect 120816 451862 120868 451868
rect 120828 439929 120856 451862
rect 120814 439920 120870 439929
rect 120814 439855 120870 439864
rect 120814 435296 120870 435305
rect 120814 435231 120870 435240
rect 120722 418976 120778 418985
rect 120722 418911 120778 418920
rect 120630 404288 120686 404297
rect 120630 404223 120686 404232
rect 120644 403034 120672 404223
rect 120632 403028 120684 403034
rect 120632 402970 120684 402976
rect 68650 391232 68706 391241
rect 68650 391167 68706 391176
rect 86314 390960 86370 390969
rect 86314 390895 86370 390904
rect 92846 390960 92902 390969
rect 102138 390960 102194 390969
rect 92902 390918 93440 390946
rect 92846 390895 92902 390904
rect 69938 390416 69994 390425
rect 68480 390374 68816 390402
rect 68480 389065 68508 390374
rect 71870 390416 71926 390425
rect 69994 390388 70288 390402
rect 69994 390374 70302 390388
rect 71760 390374 71870 390402
rect 69938 390351 69994 390360
rect 70274 390130 70302 390374
rect 80058 390416 80114 390425
rect 71926 390374 72096 390402
rect 71870 390351 71926 390360
rect 71884 390291 71912 390351
rect 70274 390102 70348 390130
rect 68466 389056 68522 389065
rect 68466 388991 68522 389000
rect 67732 374672 67784 374678
rect 67732 374614 67784 374620
rect 70320 371890 70348 390102
rect 72068 389065 72096 390374
rect 73218 390130 73246 390388
rect 73172 390102 73246 390130
rect 74644 390374 74888 390402
rect 76360 390374 76604 390402
rect 72054 389056 72110 389065
rect 72054 388991 72110 389000
rect 73066 389056 73122 389065
rect 73066 388991 73122 389000
rect 71780 388476 71832 388482
rect 71780 388418 71832 388424
rect 71792 387870 71820 388418
rect 71780 387864 71832 387870
rect 71780 387806 71832 387812
rect 71792 378026 71820 387806
rect 73080 379574 73108 388991
rect 73172 387870 73200 390102
rect 73160 387864 73212 387870
rect 73160 387806 73212 387812
rect 74644 386374 74672 390374
rect 76576 387802 76604 390374
rect 77404 390374 77832 390402
rect 79336 390374 79488 390402
rect 77404 389298 77432 390374
rect 77392 389292 77444 389298
rect 77392 389234 77444 389240
rect 76564 387796 76616 387802
rect 76564 387738 76616 387744
rect 74632 386368 74684 386374
rect 74632 386310 74684 386316
rect 72424 379568 72476 379574
rect 72424 379510 72476 379516
rect 73068 379568 73120 379574
rect 73068 379510 73120 379516
rect 71700 377998 71820 378026
rect 70308 371884 70360 371890
rect 70308 371826 70360 371832
rect 71700 356658 71728 377998
rect 70400 356652 70452 356658
rect 70400 356594 70452 356600
rect 71688 356652 71740 356658
rect 71688 356594 71740 356600
rect 70412 345014 70440 356594
rect 71700 356114 71728 356594
rect 71688 356108 71740 356114
rect 71688 356050 71740 356056
rect 71042 355328 71098 355337
rect 71042 355263 71098 355272
rect 70412 344986 70808 345014
rect 67732 338564 67784 338570
rect 67732 338506 67784 338512
rect 67744 306921 67772 338506
rect 67824 334620 67876 334626
rect 67824 334562 67876 334568
rect 67836 321609 67864 334562
rect 70030 334248 70086 334257
rect 70030 334183 70086 334192
rect 69294 331256 69350 331265
rect 69294 331191 69350 331200
rect 69112 329860 69164 329866
rect 69112 329802 69164 329808
rect 69124 327434 69152 329802
rect 69000 327406 69152 327434
rect 69308 327049 69336 331191
rect 70044 327570 70072 334183
rect 70676 330812 70728 330818
rect 70676 330754 70728 330760
rect 70688 327570 70716 330754
rect 69736 327542 70072 327570
rect 70472 327542 70716 327570
rect 70780 327162 70808 344986
rect 70780 327134 70992 327162
rect 69294 327040 69350 327049
rect 69294 326975 69350 326984
rect 69938 327040 69994 327049
rect 69938 326975 69940 326984
rect 69992 326975 69994 326984
rect 69940 326946 69992 326952
rect 70964 326890 70992 327134
rect 71056 327010 71084 355263
rect 72436 338570 72464 379510
rect 74644 373994 74672 386310
rect 74552 373966 74672 373994
rect 73804 343664 73856 343670
rect 73804 343606 73856 343612
rect 73066 339688 73122 339697
rect 73066 339623 73122 339632
rect 72424 338564 72476 338570
rect 72424 338506 72476 338512
rect 72240 331288 72292 331294
rect 72240 331230 72292 331236
rect 72252 327570 72280 331230
rect 73080 327570 73108 339623
rect 73160 335368 73212 335374
rect 73160 335310 73212 335316
rect 71944 327542 72280 327570
rect 72680 327542 73108 327570
rect 73172 327570 73200 335310
rect 73816 330818 73844 343606
rect 74552 333402 74580 373966
rect 76576 362273 76604 387738
rect 77208 385688 77260 385694
rect 77208 385630 77260 385636
rect 76562 362264 76618 362273
rect 76562 362199 76618 362208
rect 77220 359281 77248 385630
rect 77404 373994 77432 389234
rect 79336 387705 79364 390374
rect 80058 390351 80114 390360
rect 80610 390416 80666 390425
rect 80666 390374 80960 390402
rect 81452 390374 82432 390402
rect 82832 390374 83904 390402
rect 80610 390351 80666 390360
rect 80072 389201 80100 390351
rect 80058 389192 80114 389201
rect 80058 389127 80114 389136
rect 79322 387696 79378 387705
rect 79322 387631 79378 387640
rect 77312 373966 77432 373994
rect 76562 359272 76618 359281
rect 76562 359207 76618 359216
rect 77206 359272 77262 359281
rect 77206 359207 77262 359216
rect 74630 335608 74686 335617
rect 74630 335543 74686 335552
rect 74540 333396 74592 333402
rect 74540 333338 74592 333344
rect 73804 330812 73856 330818
rect 73804 330754 73856 330760
rect 74172 329996 74224 330002
rect 74172 329938 74224 329944
rect 74184 327570 74212 329938
rect 74644 327842 74672 335543
rect 76472 334688 76524 334694
rect 76472 334630 76524 334636
rect 75736 333260 75788 333266
rect 75736 333202 75788 333208
rect 74644 327814 74718 327842
rect 73172 327542 73416 327570
rect 73968 327542 74212 327570
rect 74690 327556 74718 327814
rect 75748 327570 75776 333202
rect 76484 327570 76512 334630
rect 76576 330002 76604 359207
rect 77220 358873 77248 359207
rect 77206 358864 77262 358873
rect 77206 358799 77262 358808
rect 77312 349761 77340 373966
rect 77298 349752 77354 349761
rect 77298 349687 77354 349696
rect 77208 347812 77260 347818
rect 77208 347754 77260 347760
rect 76564 329996 76616 330002
rect 76564 329938 76616 329944
rect 77220 327570 77248 347754
rect 79336 347750 79364 387631
rect 80072 364993 80100 389127
rect 81452 380866 81480 390374
rect 81440 380860 81492 380866
rect 81440 380802 81492 380808
rect 81452 379642 81480 380802
rect 81440 379636 81492 379642
rect 81440 379578 81492 379584
rect 82084 379636 82136 379642
rect 82084 379578 82136 379584
rect 81348 366376 81400 366382
rect 81348 366318 81400 366324
rect 80058 364984 80114 364993
rect 80058 364919 80114 364928
rect 79968 349852 80020 349858
rect 79968 349794 80020 349800
rect 79324 347744 79376 347750
rect 79324 347686 79376 347692
rect 78586 342272 78642 342281
rect 78586 342207 78642 342216
rect 78496 340196 78548 340202
rect 78496 340138 78548 340144
rect 77944 330268 77996 330274
rect 77944 330210 77996 330216
rect 77956 327570 77984 330210
rect 78508 327570 78536 340138
rect 78600 330274 78628 342207
rect 79876 338768 79928 338774
rect 79876 338710 79928 338716
rect 78588 330268 78640 330274
rect 78588 330210 78640 330216
rect 79416 330268 79468 330274
rect 79416 330210 79468 330216
rect 79428 327570 79456 330210
rect 79888 327570 79916 338710
rect 79980 330274 80008 349794
rect 80794 341048 80850 341057
rect 80794 340983 80850 340992
rect 80704 331152 80756 331158
rect 80704 331094 80756 331100
rect 79968 330268 80020 330274
rect 79968 330210 80020 330216
rect 80716 327570 80744 331094
rect 75440 327542 75776 327570
rect 76176 327542 76512 327570
rect 76912 327542 77248 327570
rect 77648 327542 77984 327570
rect 78384 327542 78536 327570
rect 79120 327542 79456 327570
rect 79672 327542 79916 327570
rect 80408 327542 80744 327570
rect 80808 327570 80836 340983
rect 81360 331158 81388 366318
rect 82096 365702 82124 379578
rect 81440 365696 81492 365702
rect 81440 365638 81492 365644
rect 82084 365696 82136 365702
rect 82084 365638 82136 365644
rect 81452 364410 81480 365638
rect 81440 364404 81492 364410
rect 81440 364346 81492 364352
rect 81348 331152 81400 331158
rect 81348 331094 81400 331100
rect 81452 327570 81480 364346
rect 82832 361554 82860 390374
rect 85546 390130 85574 390388
rect 85546 390102 85620 390130
rect 85592 385014 85620 390102
rect 85580 385008 85632 385014
rect 85580 384950 85632 384956
rect 86224 385008 86276 385014
rect 86224 384950 86276 384956
rect 86236 374066 86264 384950
rect 86224 374060 86276 374066
rect 86224 374002 86276 374008
rect 82820 361548 82872 361554
rect 82820 361490 82872 361496
rect 84106 360904 84162 360913
rect 84106 360839 84162 360848
rect 83464 348424 83516 348430
rect 83464 348366 83516 348372
rect 83476 331158 83504 348366
rect 82728 331152 82780 331158
rect 82728 331094 82780 331100
rect 83464 331152 83516 331158
rect 83464 331094 83516 331100
rect 82740 327570 82768 331094
rect 84120 330313 84148 360839
rect 85488 351960 85540 351966
rect 85488 351902 85540 351908
rect 85500 335354 85528 351902
rect 86236 351121 86264 374002
rect 86222 351112 86278 351121
rect 86222 351047 86278 351056
rect 86328 347002 86356 390895
rect 89810 390416 89866 390425
rect 87018 390130 87046 390388
rect 88504 390374 88932 390402
rect 86972 390102 87046 390130
rect 86972 378146 87000 390102
rect 88904 388929 88932 390374
rect 91282 390416 91338 390425
rect 89866 390374 90404 390402
rect 89810 390351 89866 390360
rect 89718 389056 89774 389065
rect 89718 388991 89774 389000
rect 88890 388920 88946 388929
rect 88890 388855 88946 388864
rect 88904 383654 88932 388855
rect 89732 387122 89760 388991
rect 90376 388793 90404 390374
rect 91338 390374 92060 390402
rect 91282 390351 91338 390360
rect 90362 388784 90418 388793
rect 90362 388719 90418 388728
rect 89720 387116 89772 387122
rect 89720 387058 89772 387064
rect 88904 383626 89024 383654
rect 86960 378140 87012 378146
rect 86960 378082 87012 378088
rect 86972 352578 87000 378082
rect 87052 362228 87104 362234
rect 87052 362170 87104 362176
rect 87972 362228 88024 362234
rect 87972 362170 88024 362176
rect 86960 352572 87012 352578
rect 86960 352514 87012 352520
rect 86866 351112 86922 351121
rect 86866 351047 86922 351056
rect 85580 346996 85632 347002
rect 85580 346938 85632 346944
rect 86316 346996 86368 347002
rect 86316 346938 86368 346944
rect 85224 335326 85528 335354
rect 84106 330304 84162 330313
rect 84106 330239 84162 330248
rect 83646 327584 83702 327593
rect 80808 327542 81144 327570
rect 81452 327542 81880 327570
rect 82616 327542 82768 327570
rect 83352 327542 83646 327570
rect 85224 327570 85252 335326
rect 85592 331158 85620 346938
rect 85670 338328 85726 338337
rect 85670 338263 85726 338272
rect 85580 331152 85632 331158
rect 85580 331094 85632 331100
rect 85684 327570 85712 338263
rect 86880 335354 86908 351047
rect 86512 335326 86908 335354
rect 86512 327593 86540 335326
rect 87064 334694 87092 362170
rect 87984 361622 88012 362170
rect 87972 361616 88024 361622
rect 87972 361558 88024 361564
rect 88996 351898 89024 383626
rect 90376 362982 90404 388719
rect 92032 383654 92060 390374
rect 93412 388482 93440 390918
rect 118698 390960 118754 390969
rect 102194 390918 102640 390946
rect 102138 390895 102194 390904
rect 97354 390416 97410 390425
rect 94240 390374 94576 390402
rect 95896 390374 96232 390402
rect 93400 388476 93452 388482
rect 93400 388418 93452 388424
rect 94240 388414 94268 390374
rect 95896 389065 95924 390374
rect 98826 390416 98882 390425
rect 97410 390374 97856 390402
rect 97354 390351 97410 390360
rect 95882 389056 95938 389065
rect 95882 388991 95938 389000
rect 93768 388408 93820 388414
rect 93768 388350 93820 388356
rect 94228 388408 94280 388414
rect 94228 388350 94280 388356
rect 92032 383626 92336 383654
rect 90364 362976 90416 362982
rect 90364 362918 90416 362924
rect 89076 352028 89128 352034
rect 89076 351970 89128 351976
rect 88984 351892 89036 351898
rect 88984 351834 89036 351840
rect 87972 343732 88024 343738
rect 87972 343674 88024 343680
rect 87052 334688 87104 334694
rect 87052 334630 87104 334636
rect 86592 331152 86644 331158
rect 86592 331094 86644 331100
rect 86498 327584 86554 327593
rect 84824 327542 85252 327570
rect 85560 327542 85712 327570
rect 86112 327542 86498 327570
rect 83646 327519 83702 327528
rect 86604 327570 86632 331094
rect 87984 327570 88012 343674
rect 89088 338774 89116 351970
rect 90376 351966 90404 362918
rect 92308 360874 92336 383626
rect 93780 364313 93808 388350
rect 96434 369608 96490 369617
rect 96434 369543 96490 369552
rect 96448 368529 96476 369543
rect 96434 368520 96490 368529
rect 96434 368455 96490 368464
rect 96448 366382 96476 368455
rect 96436 366376 96488 366382
rect 96436 366318 96488 366324
rect 93766 364304 93822 364313
rect 93766 364239 93822 364248
rect 93780 363089 93808 364239
rect 93122 363080 93178 363089
rect 93122 363015 93178 363024
rect 93766 363080 93822 363089
rect 93766 363015 93822 363024
rect 92296 360868 92348 360874
rect 92296 360810 92348 360816
rect 92386 356688 92442 356697
rect 92386 356623 92442 356632
rect 90364 351960 90416 351966
rect 90364 351902 90416 351908
rect 91008 345092 91060 345098
rect 91008 345034 91060 345040
rect 89076 338768 89128 338774
rect 89076 338710 89128 338716
rect 89442 338464 89498 338473
rect 89442 338399 89498 338408
rect 88614 334112 88670 334121
rect 88614 334047 88670 334056
rect 88628 327570 88656 334047
rect 89456 327570 89484 338399
rect 89810 335472 89866 335481
rect 89810 335407 89866 335416
rect 89824 327842 89852 335407
rect 91020 335354 91048 345034
rect 91742 336832 91798 336841
rect 91742 336767 91798 336776
rect 86604 327542 86848 327570
rect 87584 327542 88012 327570
rect 88320 327542 88656 327570
rect 89056 327542 89484 327570
rect 89778 327814 89852 327842
rect 90928 335326 91048 335354
rect 89778 327556 89806 327814
rect 90928 327570 90956 335326
rect 91756 327826 91784 336767
rect 92400 335354 92428 356623
rect 92662 353288 92718 353297
rect 92662 353223 92718 353232
rect 92676 352034 92704 353223
rect 92664 352028 92716 352034
rect 92664 351970 92716 351976
rect 93136 340202 93164 363015
rect 93768 358080 93820 358086
rect 93768 358022 93820 358028
rect 96526 358048 96582 358057
rect 93676 342304 93728 342310
rect 93676 342246 93728 342252
rect 93124 340196 93176 340202
rect 93124 340138 93176 340144
rect 92216 335326 92428 335354
rect 91744 327820 91796 327826
rect 91744 327762 91796 327768
rect 91236 327720 91292 327729
rect 91236 327655 91292 327664
rect 90528 327542 90956 327570
rect 91250 327556 91278 327655
rect 92216 327570 92244 335326
rect 92386 332480 92442 332489
rect 92386 332415 92442 332424
rect 92400 327729 92428 332415
rect 92848 330064 92900 330070
rect 92848 330006 92900 330012
rect 92386 327720 92442 327729
rect 92386 327655 92442 327664
rect 92860 327570 92888 330006
rect 93688 327570 93716 342246
rect 93780 330070 93808 358022
rect 96526 357983 96582 357992
rect 93858 353560 93914 353569
rect 93858 353495 93914 353504
rect 93768 330064 93820 330070
rect 93768 330006 93820 330012
rect 91816 327542 92244 327570
rect 92552 327542 92888 327570
rect 93288 327542 93716 327570
rect 93872 327570 93900 353495
rect 95054 333296 95110 333305
rect 95054 333231 95110 333240
rect 95068 327570 95096 333231
rect 96436 330540 96488 330546
rect 96436 330482 96488 330488
rect 95792 329996 95844 330002
rect 95792 329938 95844 329944
rect 95804 327570 95832 329938
rect 96448 327570 96476 330482
rect 96540 330002 96568 357983
rect 97828 355366 97856 390374
rect 100666 390416 100722 390425
rect 98882 390374 99328 390402
rect 98826 390351 98882 390360
rect 99300 378826 99328 390374
rect 100722 390374 101168 390402
rect 100666 390351 100722 390360
rect 101140 389065 101168 390374
rect 102612 389162 102640 390918
rect 118754 390918 119048 390946
rect 118698 390895 118754 390904
rect 115754 390688 115810 390697
rect 115810 390646 115888 390674
rect 115754 390623 115810 390632
rect 111504 390510 111656 390538
rect 105082 390416 105138 390425
rect 103776 390374 104112 390402
rect 102600 389156 102652 389162
rect 102600 389098 102652 389104
rect 101126 389056 101182 389065
rect 101126 388991 101182 389000
rect 101954 389056 102010 389065
rect 101954 388991 102010 389000
rect 100024 388476 100076 388482
rect 100024 388418 100076 388424
rect 101404 388476 101456 388482
rect 101404 388418 101456 388424
rect 99288 378820 99340 378826
rect 99288 378762 99340 378768
rect 99286 364440 99342 364449
rect 99286 364375 99342 364384
rect 99300 364334 99328 364375
rect 99300 364306 99420 364334
rect 99288 360256 99340 360262
rect 99288 360198 99340 360204
rect 97816 355360 97868 355366
rect 97816 355302 97868 355308
rect 99194 350704 99250 350713
rect 99194 350639 99250 350648
rect 97906 339552 97962 339561
rect 97906 339487 97962 339496
rect 97264 332716 97316 332722
rect 97264 332658 97316 332664
rect 96528 329996 96580 330002
rect 96528 329938 96580 329944
rect 97276 327570 97304 332658
rect 97920 327570 97948 339487
rect 98552 330404 98604 330410
rect 98552 330346 98604 330352
rect 98564 327570 98592 330346
rect 99208 327570 99236 350639
rect 99300 330410 99328 360198
rect 99392 331226 99420 364306
rect 100036 363769 100064 388418
rect 100022 363760 100078 363769
rect 100022 363695 100078 363704
rect 101416 360913 101444 388418
rect 101402 360904 101458 360913
rect 101402 360839 101458 360848
rect 101968 359009 101996 388991
rect 104084 387122 104112 390374
rect 106554 390416 106610 390425
rect 105138 390374 105676 390402
rect 105082 390351 105138 390360
rect 105544 389156 105596 389162
rect 105544 389098 105596 389104
rect 104072 387116 104124 387122
rect 104072 387058 104124 387064
rect 102046 371376 102102 371385
rect 102046 371311 102102 371320
rect 101402 359000 101458 359009
rect 101402 358935 101458 358944
rect 101954 359000 102010 359009
rect 101954 358935 102010 358944
rect 101416 333266 101444 358935
rect 101496 334008 101548 334014
rect 101496 333950 101548 333956
rect 101404 333260 101456 333266
rect 101404 333202 101456 333208
rect 99380 331220 99432 331226
rect 99380 331162 99432 331168
rect 99288 330404 99340 330410
rect 99288 330346 99340 330352
rect 99392 329866 99420 331162
rect 100022 330440 100078 330449
rect 100022 330375 100078 330384
rect 99380 329860 99432 329866
rect 99380 329802 99432 329808
rect 100036 327570 100064 330375
rect 100116 329860 100168 329866
rect 100116 329802 100168 329808
rect 93872 327542 94024 327570
rect 94760 327542 95096 327570
rect 95496 327542 95832 327570
rect 96232 327542 96476 327570
rect 96968 327542 97304 327570
rect 97520 327542 97948 327570
rect 98256 327542 98592 327570
rect 98992 327542 99236 327570
rect 99728 327542 100064 327570
rect 100128 327570 100156 329802
rect 101508 327570 101536 333950
rect 102060 327570 102088 371311
rect 104900 365764 104952 365770
rect 104900 365706 104952 365712
rect 104808 352572 104860 352578
rect 104808 352514 104860 352520
rect 102784 340944 102836 340950
rect 102784 340886 102836 340892
rect 102690 331392 102746 331401
rect 102690 331327 102746 331336
rect 102704 327842 102732 331327
rect 100128 327542 100464 327570
rect 101200 327542 101536 327570
rect 101936 327542 102088 327570
rect 102658 327814 102732 327842
rect 102658 327556 102686 327814
rect 102796 327570 102824 340886
rect 104164 329860 104216 329866
rect 104164 329802 104216 329808
rect 104176 327570 104204 329802
rect 104820 327570 104848 352514
rect 104912 345014 104940 365706
rect 105556 345681 105584 389098
rect 105648 381546 105676 390374
rect 108026 390416 108082 390425
rect 106610 390374 107332 390402
rect 106554 390351 106610 390360
rect 107304 383654 107332 390374
rect 109498 390416 109554 390425
rect 108082 390374 108804 390402
rect 108026 390351 108082 390360
rect 108776 383654 108804 390374
rect 109554 390374 110276 390402
rect 109498 390351 109554 390360
rect 107304 383626 107516 383654
rect 108776 383626 108896 383654
rect 105636 381540 105688 381546
rect 105636 381482 105688 381488
rect 107488 351121 107516 383626
rect 108304 378888 108356 378894
rect 108304 378830 108356 378836
rect 107474 351112 107530 351121
rect 107474 351047 107530 351056
rect 105542 345672 105598 345681
rect 105542 345607 105598 345616
rect 108316 345014 108344 378830
rect 108868 370705 108896 383626
rect 110248 382974 110276 390374
rect 111628 389230 111656 390510
rect 112640 390374 112976 390402
rect 114112 390374 114448 390402
rect 111708 389836 111760 389842
rect 111708 389778 111760 389784
rect 111616 389224 111668 389230
rect 111616 389166 111668 389172
rect 111628 387870 111656 389166
rect 111616 387864 111668 387870
rect 111616 387806 111668 387812
rect 110236 382968 110288 382974
rect 110236 382910 110288 382916
rect 108854 370696 108910 370705
rect 108854 370631 108910 370640
rect 109682 358728 109738 358737
rect 109682 358663 109738 358672
rect 109696 357513 109724 358663
rect 109682 357504 109738 357513
rect 109682 357439 109738 357448
rect 108946 349344 109002 349353
rect 108946 349279 109002 349288
rect 104912 344986 105032 345014
rect 102796 327542 103224 327570
rect 103960 327542 104204 327570
rect 104696 327542 104848 327570
rect 105004 327570 105032 344986
rect 107856 344986 108344 345014
rect 105542 342408 105598 342417
rect 105542 342343 105598 342352
rect 105556 329866 105584 342343
rect 107856 339833 107884 344986
rect 108854 343768 108910 343777
rect 108854 343703 108910 343712
rect 107842 339824 107898 339833
rect 107842 339759 107898 339768
rect 106464 338156 106516 338162
rect 106464 338098 106516 338104
rect 106002 332616 106058 332625
rect 106002 332551 106058 332560
rect 105544 329860 105596 329866
rect 105544 329802 105596 329808
rect 106016 327570 106044 332551
rect 106476 327570 106504 338098
rect 107856 327570 107884 339759
rect 108580 329860 108632 329866
rect 108580 329802 108632 329808
rect 108592 327570 108620 329802
rect 108868 327842 108896 343703
rect 108960 329866 108988 349279
rect 109696 348430 109724 357439
rect 111338 356144 111394 356153
rect 111338 356079 111394 356088
rect 110418 355872 110474 355881
rect 110418 355807 110474 355816
rect 109684 348424 109736 348430
rect 109684 348366 109736 348372
rect 110432 345014 110460 355807
rect 111352 349858 111380 356079
rect 111720 355881 111748 389778
rect 112640 389065 112668 390374
rect 111798 389056 111854 389065
rect 111798 388991 111854 389000
rect 112626 389056 112682 389065
rect 112626 388991 112682 389000
rect 111812 356726 111840 388991
rect 114112 388657 114140 390374
rect 113178 388648 113234 388657
rect 113178 388583 113234 388592
rect 114098 388648 114154 388657
rect 114098 388583 114154 388592
rect 112444 387864 112496 387870
rect 112444 387806 112496 387812
rect 111800 356720 111852 356726
rect 111800 356662 111852 356668
rect 111706 355872 111762 355881
rect 111706 355807 111762 355816
rect 111720 354793 111748 355807
rect 111706 354784 111762 354793
rect 111706 354719 111762 354728
rect 112456 349858 112484 387806
rect 113192 385694 113220 388583
rect 113180 385688 113232 385694
rect 113180 385630 113232 385636
rect 115860 352073 115888 390646
rect 115938 390416 115994 390425
rect 115994 390374 116104 390402
rect 117576 390374 117912 390402
rect 115938 390351 115994 390360
rect 114558 352064 114614 352073
rect 114558 351999 114614 352008
rect 115846 352064 115902 352073
rect 115846 351999 115902 352008
rect 111340 349852 111392 349858
rect 111340 349794 111392 349800
rect 112444 349852 112496 349858
rect 112444 349794 112496 349800
rect 113086 347984 113142 347993
rect 113086 347919 113142 347928
rect 110432 344986 110736 345014
rect 109958 330304 110014 330313
rect 109958 330239 110014 330248
rect 108948 329860 109000 329866
rect 108948 329802 109000 329808
rect 108868 327814 108942 327842
rect 105004 327542 105432 327570
rect 106016 327542 106168 327570
rect 106476 327542 106904 327570
rect 107640 327542 107884 327570
rect 108376 327542 108620 327570
rect 108914 327556 108942 327814
rect 109972 327570 110000 330239
rect 110604 330132 110656 330138
rect 110604 330074 110656 330080
rect 110616 327570 110644 330074
rect 109664 327542 110000 327570
rect 110400 327542 110644 327570
rect 110708 327570 110736 344986
rect 111706 340912 111762 340921
rect 111706 340847 111762 340856
rect 111720 330138 111748 340847
rect 113100 335354 113128 347919
rect 114572 345014 114600 351999
rect 115952 345817 115980 390351
rect 117884 389162 117912 390374
rect 117872 389156 117924 389162
rect 117872 389098 117924 389104
rect 118712 382294 118740 390895
rect 120736 390697 120764 418911
rect 120722 390688 120778 390697
rect 120722 390623 120778 390632
rect 120170 390416 120226 390425
rect 120226 390374 120520 390402
rect 120170 390351 120226 390360
rect 120184 388482 120212 390351
rect 120172 388476 120224 388482
rect 120172 388418 120224 388424
rect 118700 382288 118752 382294
rect 118700 382230 118752 382236
rect 119436 382288 119488 382294
rect 119436 382230 119488 382236
rect 119342 368384 119398 368393
rect 119342 368319 119398 368328
rect 118700 360868 118752 360874
rect 118700 360810 118752 360816
rect 118712 357474 118740 360810
rect 118700 357468 118752 357474
rect 118700 357410 118752 357416
rect 117318 349208 117374 349217
rect 117318 349143 117374 349152
rect 115938 345808 115994 345817
rect 115938 345743 115994 345752
rect 115204 345160 115256 345166
rect 115204 345102 115256 345108
rect 114572 344986 114692 345014
rect 114468 339584 114520 339590
rect 114468 339526 114520 339532
rect 113008 335326 113128 335354
rect 112166 334384 112222 334393
rect 112166 334319 112222 334328
rect 111708 330132 111760 330138
rect 111708 330074 111760 330080
rect 112180 327570 112208 334319
rect 113008 327570 113036 335326
rect 114376 331152 114428 331158
rect 114376 331094 114428 331100
rect 113640 329996 113692 330002
rect 113640 329938 113692 329944
rect 113652 327570 113680 329938
rect 114388 327570 114416 331094
rect 114480 330002 114508 339526
rect 114468 329996 114520 330002
rect 114468 329938 114520 329944
rect 114664 327842 114692 344986
rect 114742 335744 114798 335753
rect 114742 335679 114798 335688
rect 114756 331158 114784 335679
rect 115216 334626 115244 345102
rect 117332 345014 117360 349143
rect 118606 345128 118662 345137
rect 118606 345063 118662 345072
rect 117332 344986 117912 345014
rect 115940 336864 115992 336870
rect 115940 336806 115992 336812
rect 115296 335436 115348 335442
rect 115296 335378 115348 335384
rect 115204 334620 115256 334626
rect 115204 334562 115256 334568
rect 114744 331152 114796 331158
rect 114744 331094 114796 331100
rect 115308 328438 115336 335378
rect 115664 332648 115716 332654
rect 115664 332590 115716 332596
rect 115296 328432 115348 328438
rect 115296 328374 115348 328380
rect 114618 327814 114692 327842
rect 114618 327570 114646 327814
rect 115676 327570 115704 332590
rect 110708 327542 111136 327570
rect 111872 327542 112208 327570
rect 112608 327542 113036 327570
rect 113344 327542 113680 327570
rect 114080 327542 114416 327570
rect 114480 327556 114646 327570
rect 114480 327542 114632 327556
rect 115368 327542 115704 327570
rect 115952 327570 115980 336806
rect 117134 332752 117190 332761
rect 117134 332687 117190 332696
rect 117148 327570 117176 332687
rect 117780 330268 117832 330274
rect 117780 330210 117832 330216
rect 117792 327570 117820 330210
rect 115952 327542 116104 327570
rect 116840 327542 117176 327570
rect 117576 327542 117820 327570
rect 117884 327570 117912 344986
rect 118620 330274 118648 345063
rect 118608 330268 118660 330274
rect 118608 330210 118660 330216
rect 118712 327570 118740 357410
rect 119356 350606 119384 368319
rect 119448 367810 119476 382230
rect 120828 375465 120856 435231
rect 121472 396953 121500 548490
rect 121564 428505 121592 578206
rect 123484 569220 123536 569226
rect 123484 569162 123536 569168
rect 122104 556232 122156 556238
rect 122104 556174 122156 556180
rect 121644 453348 121696 453354
rect 121644 453290 121696 453296
rect 121550 428496 121606 428505
rect 121550 428431 121606 428440
rect 121552 418124 121604 418130
rect 121552 418066 121604 418072
rect 121564 417353 121592 418066
rect 121550 417344 121606 417353
rect 121550 417279 121606 417288
rect 121458 396944 121514 396953
rect 121458 396879 121514 396888
rect 121472 396098 121500 396879
rect 121460 396092 121512 396098
rect 121460 396034 121512 396040
rect 121564 389842 121592 417279
rect 121656 410553 121684 453290
rect 121642 410544 121698 410553
rect 121642 410479 121698 410488
rect 121656 409902 121684 410479
rect 121644 409896 121696 409902
rect 121644 409838 121696 409844
rect 122116 407114 122144 556174
rect 122932 512644 122984 512650
rect 122932 512586 122984 512592
rect 122944 433129 122972 512586
rect 123024 457496 123076 457502
rect 123024 457438 123076 457444
rect 122930 433120 122986 433129
rect 122930 433055 122986 433064
rect 122838 428496 122894 428505
rect 122838 428431 122894 428440
rect 122104 407108 122156 407114
rect 122104 407050 122156 407056
rect 122654 393272 122710 393281
rect 122654 393207 122710 393216
rect 121552 389836 121604 389842
rect 121552 389778 121604 389784
rect 122668 385665 122696 393207
rect 122746 392592 122802 392601
rect 122746 392527 122802 392536
rect 122654 385656 122710 385665
rect 122654 385591 122710 385600
rect 120814 375456 120870 375465
rect 120814 375391 120870 375400
rect 120828 373994 120856 375391
rect 120736 373966 120856 373994
rect 119436 367804 119488 367810
rect 119436 367746 119488 367752
rect 120080 354748 120132 354754
rect 120080 354690 120132 354696
rect 118792 350600 118844 350606
rect 118792 350542 118844 350548
rect 119344 350600 119396 350606
rect 119344 350542 119396 350548
rect 118804 345014 118832 350542
rect 118804 344986 119292 345014
rect 119264 327570 119292 344986
rect 119342 343904 119398 343913
rect 119342 343839 119398 343848
rect 119356 330449 119384 343839
rect 119342 330440 119398 330449
rect 119342 330375 119398 330384
rect 120092 327570 120120 354690
rect 120736 352578 120764 373966
rect 122760 372638 122788 392527
rect 122104 372632 122156 372638
rect 122104 372574 122156 372580
rect 122748 372632 122800 372638
rect 122748 372574 122800 372580
rect 121368 368552 121420 368558
rect 121368 368494 121420 368500
rect 120724 352572 120776 352578
rect 120724 352514 120776 352520
rect 121380 327570 121408 368494
rect 121458 361720 121514 361729
rect 121458 361655 121514 361664
rect 121472 356697 121500 361655
rect 121458 356688 121514 356697
rect 121458 356623 121514 356632
rect 121644 347880 121696 347886
rect 121644 347822 121696 347828
rect 121656 347750 121684 347822
rect 121644 347744 121696 347750
rect 121644 347686 121696 347692
rect 122116 331906 122144 372574
rect 122852 370569 122880 428431
rect 123036 424153 123064 457438
rect 123208 456068 123260 456074
rect 123208 456010 123260 456016
rect 123022 424144 123078 424153
rect 122944 424102 123022 424130
rect 122944 412634 122972 424102
rect 123022 424079 123078 424088
rect 123024 422340 123076 422346
rect 123024 422282 123076 422288
rect 123036 421977 123064 422282
rect 123022 421968 123078 421977
rect 123022 421903 123078 421912
rect 123116 413976 123168 413982
rect 123116 413918 123168 413924
rect 123128 412729 123156 413918
rect 123114 412720 123170 412729
rect 123114 412655 123170 412664
rect 122944 412606 123064 412634
rect 122932 407108 122984 407114
rect 122932 407050 122984 407056
rect 122944 392601 122972 407050
rect 122930 392592 122986 392601
rect 122930 392527 122986 392536
rect 123036 380225 123064 412606
rect 123128 384334 123156 412655
rect 123220 406201 123248 456010
rect 123496 422346 123524 569162
rect 124220 567860 124272 567866
rect 124220 567802 124272 567808
rect 124128 444372 124180 444378
rect 124128 444314 124180 444320
rect 124140 444281 124168 444314
rect 124126 444272 124182 444281
rect 124126 444207 124182 444216
rect 124126 442096 124182 442105
rect 124126 442031 124182 442040
rect 124140 441658 124168 442031
rect 124128 441652 124180 441658
rect 124128 441594 124180 441600
rect 124126 439920 124182 439929
rect 124126 439855 124182 439864
rect 124140 438938 124168 439855
rect 124128 438932 124180 438938
rect 124128 438874 124180 438880
rect 124128 438184 124180 438190
rect 124128 438126 124180 438132
rect 124140 437753 124168 438126
rect 124126 437744 124182 437753
rect 124126 437679 124182 437688
rect 124126 433120 124182 433129
rect 124126 433055 124182 433064
rect 124140 432614 124168 433055
rect 124128 432608 124180 432614
rect 124128 432550 124180 432556
rect 123484 422340 123536 422346
rect 123484 422282 123536 422288
rect 124128 415200 124180 415206
rect 124126 415168 124128 415177
rect 124180 415168 124182 415177
rect 124126 415103 124182 415112
rect 124126 408368 124182 408377
rect 124232 408354 124260 567802
rect 124876 536790 124904 702986
rect 126244 702908 126296 702914
rect 126244 702850 126296 702856
rect 125600 557592 125652 557598
rect 125600 557534 125652 557540
rect 124864 536784 124916 536790
rect 124864 536726 124916 536732
rect 124864 458244 124916 458250
rect 124864 458186 124916 458192
rect 124312 447840 124364 447846
rect 124312 447782 124364 447788
rect 124324 438190 124352 447782
rect 124312 438184 124364 438190
rect 124312 438126 124364 438132
rect 124182 408326 124260 408354
rect 124126 408303 124182 408312
rect 124140 407794 124168 408303
rect 124128 407788 124180 407794
rect 124128 407730 124180 407736
rect 123206 406192 123262 406201
rect 123206 406127 123208 406136
rect 123260 406127 123262 406136
rect 123208 406098 123260 406104
rect 123220 406067 123248 406098
rect 124126 401568 124182 401577
rect 124126 401503 124128 401512
rect 124180 401503 124182 401512
rect 124128 401474 124180 401480
rect 123482 399392 123538 399401
rect 123482 399327 123538 399336
rect 123496 398886 123524 399327
rect 123484 398880 123536 398886
rect 123484 398822 123536 398828
rect 123668 395548 123720 395554
rect 123668 395490 123720 395496
rect 123680 394777 123708 395490
rect 123666 394768 123722 394777
rect 123666 394703 123722 394712
rect 123116 384328 123168 384334
rect 123116 384270 123168 384276
rect 123022 380216 123078 380225
rect 123022 380151 123078 380160
rect 122838 370560 122894 370569
rect 122838 370495 122894 370504
rect 122930 367704 122986 367713
rect 122930 367639 122986 367648
rect 122656 354000 122708 354006
rect 122656 353942 122708 353948
rect 122196 339516 122248 339522
rect 122196 339458 122248 339464
rect 122104 331900 122156 331906
rect 122104 331842 122156 331848
rect 122104 330608 122156 330614
rect 122104 330550 122156 330556
rect 122116 327570 122144 330550
rect 122208 329798 122236 339458
rect 122196 329792 122248 329798
rect 122196 329734 122248 329740
rect 122668 327570 122696 353942
rect 122748 347880 122800 347886
rect 122748 347822 122800 347828
rect 122760 347774 122788 347822
rect 122760 347746 122880 347774
rect 117884 327542 118312 327570
rect 118712 327542 119048 327570
rect 119264 327542 119784 327570
rect 120092 327542 120336 327570
rect 121072 327542 121408 327570
rect 121808 327542 122144 327570
rect 122544 327542 122696 327570
rect 86498 327519 86554 327528
rect 86512 327459 86540 327519
rect 83922 327176 83978 327185
rect 83978 327134 84088 327162
rect 83922 327111 83978 327120
rect 93872 327078 93900 327542
rect 114480 327457 114508 327542
rect 114466 327448 114522 327457
rect 114466 327383 114522 327392
rect 122852 327321 122880 347746
rect 122944 328681 122972 367639
rect 124876 365838 124904 458186
rect 124956 445868 125008 445874
rect 124956 445810 125008 445816
rect 124968 406337 124996 445810
rect 124954 406328 125010 406337
rect 124954 406263 125010 406272
rect 125048 406156 125100 406162
rect 125048 406098 125100 406104
rect 124956 398880 125008 398886
rect 124956 398822 125008 398828
rect 124968 392018 124996 398822
rect 124956 392012 125008 392018
rect 124956 391954 125008 391960
rect 124968 391406 124996 391954
rect 124956 391400 125008 391406
rect 124956 391342 125008 391348
rect 124956 374672 125008 374678
rect 124956 374614 125008 374620
rect 124864 365832 124916 365838
rect 124864 365774 124916 365780
rect 123298 360224 123354 360233
rect 123298 360159 123354 360168
rect 123312 355337 123340 360159
rect 123298 355328 123354 355337
rect 123298 355263 123354 355272
rect 124876 330546 124904 365774
rect 124968 360330 124996 374614
rect 125060 371278 125088 406098
rect 125612 395554 125640 557534
rect 126256 545766 126284 702850
rect 129004 702704 129056 702710
rect 129004 702646 129056 702652
rect 126980 571396 127032 571402
rect 126980 571338 127032 571344
rect 126244 545760 126296 545766
rect 126244 545702 126296 545708
rect 125692 463004 125744 463010
rect 125692 462946 125744 462952
rect 125704 415206 125732 462946
rect 126244 444508 126296 444514
rect 126244 444450 126296 444456
rect 125692 415200 125744 415206
rect 125692 415142 125744 415148
rect 125600 395548 125652 395554
rect 125600 395490 125652 395496
rect 125048 371272 125100 371278
rect 125048 371214 125100 371220
rect 125508 371272 125560 371278
rect 125508 371214 125560 371220
rect 124956 360324 125008 360330
rect 124956 360266 125008 360272
rect 124864 330540 124916 330546
rect 124864 330482 124916 330488
rect 122930 328672 122986 328681
rect 122930 328607 122986 328616
rect 122944 327434 122972 328607
rect 124968 328545 124996 360266
rect 125520 352034 125548 371214
rect 125600 369912 125652 369918
rect 125600 369854 125652 369860
rect 125508 352028 125560 352034
rect 125508 351970 125560 351976
rect 125506 338192 125562 338201
rect 125506 338127 125562 338136
rect 124954 328536 125010 328545
rect 124954 328471 125010 328480
rect 124968 327570 124996 328471
rect 125520 327842 125548 338127
rect 124752 327542 124996 327570
rect 125474 327814 125548 327842
rect 125474 327556 125502 327814
rect 125612 327570 125640 369854
rect 125704 358057 125732 415142
rect 126256 369918 126284 444450
rect 126992 418130 127020 571338
rect 128360 569968 128412 569974
rect 128360 569910 128412 569916
rect 127624 452668 127676 452674
rect 127624 452610 127676 452616
rect 126980 418124 127032 418130
rect 126980 418066 127032 418072
rect 126244 369912 126296 369918
rect 126244 369854 126296 369860
rect 127636 367169 127664 452610
rect 128372 413982 128400 569910
rect 129016 544406 129044 702646
rect 129740 563100 129792 563106
rect 129740 563042 129792 563048
rect 129004 544400 129056 544406
rect 129004 544342 129056 544348
rect 129002 536072 129058 536081
rect 129002 536007 129058 536016
rect 128360 413976 128412 413982
rect 128360 413918 128412 413924
rect 127622 367160 127678 367169
rect 127622 367095 127678 367104
rect 125690 358048 125746 358057
rect 125690 357983 125746 357992
rect 127636 354006 127664 367095
rect 129016 364313 129044 536007
rect 129096 409896 129148 409902
rect 129096 409838 129148 409844
rect 129002 364304 129058 364313
rect 129002 364239 129058 364248
rect 129016 363633 129044 364239
rect 129002 363624 129058 363633
rect 129002 363559 129058 363568
rect 127716 359508 127768 359514
rect 127716 359450 127768 359456
rect 127624 354000 127676 354006
rect 127624 353942 127676 353948
rect 125692 352028 125744 352034
rect 125692 351970 125744 351976
rect 125704 345014 125732 351970
rect 127728 350577 127756 359450
rect 128360 358896 128412 358902
rect 128360 358838 128412 358844
rect 126978 350568 127034 350577
rect 126978 350503 127034 350512
rect 127714 350568 127770 350577
rect 127714 350503 127770 350512
rect 125704 344986 126376 345014
rect 126348 327570 126376 344986
rect 126992 331158 127020 350503
rect 128372 345014 128400 358838
rect 129108 356697 129136 409838
rect 129752 401538 129780 563042
rect 130396 536761 130424 703190
rect 133144 700324 133196 700330
rect 133144 700266 133196 700272
rect 132498 582992 132554 583001
rect 132498 582927 132554 582936
rect 130382 536752 130438 536761
rect 130382 536687 130438 536696
rect 132512 444378 132540 582927
rect 133156 538218 133184 700266
rect 134524 552084 134576 552090
rect 134524 552026 134576 552032
rect 133144 538212 133196 538218
rect 133144 538154 133196 538160
rect 132500 444372 132552 444378
rect 132500 444314 132552 444320
rect 133788 444372 133840 444378
rect 133788 444314 133840 444320
rect 133800 443698 133828 444314
rect 133788 443692 133840 443698
rect 133788 443634 133840 443640
rect 133144 441652 133196 441658
rect 133144 441594 133196 441600
rect 129740 401532 129792 401538
rect 129740 401474 129792 401480
rect 129752 400246 129780 401474
rect 129740 400240 129792 400246
rect 129740 400182 129792 400188
rect 130384 400240 130436 400246
rect 130384 400182 130436 400188
rect 130396 358193 130424 400182
rect 133156 377369 133184 441594
rect 134536 389162 134564 552026
rect 136652 541686 136680 703582
rect 137664 703474 137692 703582
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202604 703588 202656 703594
rect 202604 703530 202656 703536
rect 137848 703474 137876 703520
rect 137664 703446 137876 703474
rect 154132 702545 154160 703520
rect 154118 702536 154174 702545
rect 154118 702471 154174 702480
rect 170324 702434 170352 703520
rect 202616 703474 202644 703530
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234988 703656 235040 703662
rect 234988 703598 235040 703604
rect 202800 703474 202828 703520
rect 202616 703446 202828 703474
rect 169772 702406 170352 702434
rect 169772 596834 169800 702406
rect 218992 700330 219020 703520
rect 235000 703474 235028 703598
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267464 703520 267516 703526
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 703474 267688 703520
rect 267516 703468 267688 703474
rect 267464 703462 267688 703468
rect 267476 703446 267688 703462
rect 283852 703390 283880 703520
rect 300136 703458 300164 703520
rect 300124 703452 300176 703458
rect 300124 703394 300176 703400
rect 283840 703384 283892 703390
rect 283840 703326 283892 703332
rect 332520 703322 332548 703520
rect 332508 703316 332560 703322
rect 332508 703258 332560 703264
rect 348804 703186 348832 703520
rect 348792 703180 348844 703186
rect 348792 703122 348844 703128
rect 364996 702982 365024 703520
rect 397472 703118 397500 703520
rect 413664 703254 413692 703520
rect 413652 703248 413704 703254
rect 413652 703190 413704 703196
rect 397460 703112 397512 703118
rect 397460 703054 397512 703060
rect 429856 703050 429884 703520
rect 429844 703044 429896 703050
rect 429844 702986 429896 702992
rect 364984 702976 365036 702982
rect 364984 702918 365036 702924
rect 462332 702914 462360 703520
rect 462320 702908 462372 702914
rect 462320 702850 462372 702856
rect 478524 702778 478552 703520
rect 494808 702846 494836 703520
rect 494796 702840 494848 702846
rect 494796 702782 494848 702788
rect 478512 702772 478564 702778
rect 478512 702714 478564 702720
rect 527192 702642 527220 703520
rect 543476 702710 543504 703520
rect 543464 702704 543516 702710
rect 543464 702646 543516 702652
rect 527180 702636 527232 702642
rect 527180 702578 527232 702584
rect 559668 702506 559696 703520
rect 580264 702568 580316 702574
rect 580264 702510 580316 702516
rect 559656 702500 559708 702506
rect 559656 702442 559708 702448
rect 218980 700324 219032 700330
rect 218980 700266 219032 700272
rect 580276 670721 580304 702510
rect 582378 697232 582434 697241
rect 582378 697167 582434 697176
rect 580262 670712 580318 670721
rect 580262 670647 580318 670656
rect 169760 596828 169812 596834
rect 169760 596770 169812 596776
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580184 589937 580212 590951
rect 580170 589928 580226 589937
rect 580170 589863 580226 589872
rect 580262 577688 580318 577697
rect 580262 577623 580318 577632
rect 136640 541680 136692 541686
rect 136640 541622 136692 541628
rect 135168 432608 135220 432614
rect 135168 432550 135220 432556
rect 134524 389156 134576 389162
rect 134524 389098 134576 389104
rect 135076 387116 135128 387122
rect 135076 387058 135128 387064
rect 133142 377360 133198 377369
rect 133142 377295 133198 377304
rect 131120 363044 131172 363050
rect 131120 362986 131172 362992
rect 130382 358184 130438 358193
rect 130382 358119 130438 358128
rect 131132 358086 131160 362986
rect 131120 358080 131172 358086
rect 131120 358022 131172 358028
rect 129094 356688 129150 356697
rect 129094 356623 129150 356632
rect 129646 354920 129702 354929
rect 129646 354855 129702 354864
rect 129660 351898 129688 354855
rect 132408 353320 132460 353326
rect 132408 353262 132460 353268
rect 129648 351892 129700 351898
rect 129648 351834 129700 351840
rect 129660 350554 129688 351834
rect 129660 350526 129780 350554
rect 128372 344986 128584 345014
rect 127072 335436 127124 335442
rect 127072 335378 127124 335384
rect 126980 331152 127032 331158
rect 126980 331094 127032 331100
rect 127084 327570 127112 335378
rect 127900 331152 127952 331158
rect 127900 331094 127952 331100
rect 127912 327570 127940 331094
rect 128556 327570 128584 344986
rect 129752 327842 129780 350526
rect 130016 341012 130068 341018
rect 130016 340954 130068 340960
rect 129706 327814 129780 327842
rect 125612 327542 126040 327570
rect 126348 327542 126776 327570
rect 127084 327542 127512 327570
rect 127912 327542 128248 327570
rect 128556 327542 128984 327570
rect 129706 327556 129734 327814
rect 130028 327570 130056 340954
rect 132038 330440 132094 330449
rect 132038 330375 132094 330384
rect 131488 329860 131540 329866
rect 131488 329802 131540 329808
rect 131500 327570 131528 329802
rect 132052 327570 132080 330375
rect 132420 329866 132448 353262
rect 133880 349172 133932 349178
rect 133880 349114 133932 349120
rect 133892 345014 133920 349114
rect 133892 344986 134288 345014
rect 132776 339516 132828 339522
rect 132776 339458 132828 339464
rect 132684 329928 132736 329934
rect 132684 329870 132736 329876
rect 132408 329860 132460 329866
rect 132408 329802 132460 329808
rect 132696 327570 132724 329870
rect 130028 327542 130456 327570
rect 131192 327542 131528 327570
rect 131744 327542 132080 327570
rect 132480 327542 132724 327570
rect 132788 327570 132816 339458
rect 133788 331356 133840 331362
rect 133788 331298 133840 331304
rect 133800 329798 133828 331298
rect 134156 329860 134208 329866
rect 134156 329802 134208 329808
rect 133788 329792 133840 329798
rect 133788 329734 133840 329740
rect 133878 328536 133934 328545
rect 133878 328471 133934 328480
rect 133892 327758 133920 328471
rect 133880 327752 133932 327758
rect 133880 327694 133932 327700
rect 134168 327570 134196 329802
rect 132788 327542 133216 327570
rect 133952 327542 134196 327570
rect 134260 327570 134288 344986
rect 135088 328681 135116 387058
rect 135180 347041 135208 432550
rect 135904 407788 135956 407794
rect 135904 407730 135956 407736
rect 135916 367033 135944 407730
rect 136652 387122 136680 541622
rect 579802 537840 579858 537849
rect 579802 537775 579858 537784
rect 579816 537538 579844 537775
rect 579804 537532 579856 537538
rect 579804 537474 579856 537480
rect 580276 534070 580304 577623
rect 582392 536081 582420 697167
rect 582470 683904 582526 683913
rect 582470 683839 582526 683848
rect 582484 577522 582512 683839
rect 582562 644056 582618 644065
rect 582562 643991 582618 644000
rect 582472 577516 582524 577522
rect 582472 577458 582524 577464
rect 582472 554804 582524 554810
rect 582472 554746 582524 554752
rect 582378 536072 582434 536081
rect 582378 536007 582434 536016
rect 580264 534064 580316 534070
rect 580264 534006 580316 534012
rect 582484 524521 582512 554746
rect 582576 538286 582604 643991
rect 582654 630864 582710 630873
rect 582654 630799 582710 630808
rect 582668 540938 582696 630799
rect 582746 617536 582802 617545
rect 582746 617471 582802 617480
rect 582760 595474 582788 617471
rect 582748 595468 582800 595474
rect 582748 595410 582800 595416
rect 582746 593464 582802 593473
rect 582746 593399 582802 593408
rect 582760 564369 582788 593399
rect 582746 564360 582802 564369
rect 582746 564295 582802 564304
rect 582656 540932 582708 540938
rect 582656 540874 582708 540880
rect 582564 538280 582616 538286
rect 582564 538222 582616 538228
rect 582470 524512 582526 524521
rect 582470 524447 582526 524456
rect 580170 511320 580226 511329
rect 580170 511255 580172 511264
rect 580224 511255 580226 511264
rect 580172 511226 580224 511232
rect 582378 484664 582434 484673
rect 582378 484599 582434 484608
rect 151084 456816 151136 456822
rect 151084 456758 151136 456764
rect 144184 449948 144236 449954
rect 144184 449890 144236 449896
rect 142802 448624 142858 448633
rect 142802 448559 142858 448568
rect 137282 444544 137338 444553
rect 137282 444479 137338 444488
rect 136640 387116 136692 387122
rect 136640 387058 136692 387064
rect 135902 367024 135958 367033
rect 135902 366959 135958 366968
rect 136546 367024 136602 367033
rect 136546 366959 136602 366968
rect 136560 365809 136588 366959
rect 136546 365800 136602 365809
rect 136546 365735 136602 365744
rect 136560 349897 136588 365735
rect 137296 362710 137324 444479
rect 139308 369980 139360 369986
rect 139308 369922 139360 369928
rect 137928 367124 137980 367130
rect 137928 367066 137980 367072
rect 137284 362704 137336 362710
rect 137284 362646 137336 362652
rect 137836 362704 137888 362710
rect 137836 362646 137888 362652
rect 137848 361690 137876 362646
rect 137836 361684 137888 361690
rect 137836 361626 137888 361632
rect 136640 358828 136692 358834
rect 136640 358770 136692 358776
rect 136546 349888 136602 349897
rect 136546 349823 136602 349832
rect 135166 347032 135222 347041
rect 135166 346967 135222 346976
rect 136652 345014 136680 358770
rect 137282 345264 137338 345273
rect 137282 345199 137338 345208
rect 136652 344986 137048 345014
rect 135166 342544 135222 342553
rect 135166 342479 135222 342488
rect 135180 329866 135208 342479
rect 135258 337104 135314 337113
rect 135258 337039 135314 337048
rect 135272 329866 135300 337039
rect 136916 329928 136968 329934
rect 136916 329870 136968 329876
rect 135168 329860 135220 329866
rect 135168 329802 135220 329808
rect 135260 329860 135312 329866
rect 135260 329802 135312 329808
rect 135812 329860 135864 329866
rect 135812 329802 135864 329808
rect 135260 329112 135312 329118
rect 135260 329054 135312 329060
rect 135074 328672 135130 328681
rect 135074 328607 135130 328616
rect 135272 327570 135300 329054
rect 135824 327570 135852 329802
rect 136928 327706 136956 329870
rect 136882 327678 136956 327706
rect 134260 327542 134688 327570
rect 135272 327542 135576 327570
rect 135824 327542 136160 327570
rect 136882 327556 136910 327678
rect 137020 327570 137048 344986
rect 137296 330614 137324 345199
rect 137848 331158 137876 361626
rect 137836 331152 137888 331158
rect 137836 331094 137888 331100
rect 137284 330608 137336 330614
rect 137284 330550 137336 330556
rect 137940 329934 137968 367066
rect 138018 349888 138074 349897
rect 138018 349823 138074 349832
rect 137928 329928 137980 329934
rect 137928 329870 137980 329876
rect 138032 327570 138060 349823
rect 139320 327570 139348 369922
rect 142816 369170 142844 448559
rect 142804 369164 142856 369170
rect 142804 369106 142856 369112
rect 143448 364472 143500 364478
rect 143448 364414 143500 364420
rect 141424 356176 141476 356182
rect 141424 356118 141476 356124
rect 141332 334076 141384 334082
rect 141332 334018 141384 334024
rect 139400 331152 139452 331158
rect 139400 331094 139452 331100
rect 137020 327542 137448 327570
rect 138032 327542 138184 327570
rect 138920 327542 139348 327570
rect 139412 327570 139440 331094
rect 140688 329860 140740 329866
rect 140688 329802 140740 329808
rect 140700 327570 140728 329802
rect 141344 327570 141372 334018
rect 141436 329866 141464 356118
rect 142066 353424 142122 353433
rect 142066 353359 142122 353368
rect 141424 329860 141476 329866
rect 141424 329802 141476 329808
rect 141974 328808 142030 328817
rect 141974 328743 142030 328752
rect 141988 328438 142016 328743
rect 141976 328432 142028 328438
rect 141976 328374 142028 328380
rect 142080 327570 142108 353359
rect 143354 331528 143410 331537
rect 143354 331463 143410 331472
rect 143368 330449 143396 331463
rect 143354 330440 143410 330449
rect 143354 330375 143410 330384
rect 142802 330168 142858 330177
rect 142802 330103 142858 330112
rect 142816 329089 142844 330103
rect 142894 330032 142950 330041
rect 142894 329967 142950 329976
rect 142802 329080 142858 329089
rect 142802 329015 142858 329024
rect 142908 327570 142936 329967
rect 143460 327570 143488 364414
rect 144196 352034 144224 449890
rect 145562 376000 145618 376009
rect 145562 375935 145618 375944
rect 144184 352028 144236 352034
rect 144184 351970 144236 351976
rect 145576 349761 145604 375935
rect 151096 360913 151124 456758
rect 152464 455456 152516 455462
rect 152464 455398 152516 455404
rect 151726 363760 151782 363769
rect 151726 363695 151782 363704
rect 151082 360904 151138 360913
rect 151082 360839 151138 360848
rect 151740 357377 151768 363695
rect 151174 357368 151230 357377
rect 151174 357303 151230 357312
rect 151726 357368 151782 357377
rect 151726 357303 151782 357312
rect 146300 352028 146352 352034
rect 146300 351970 146352 351976
rect 144918 349752 144974 349761
rect 144918 349687 144974 349696
rect 145562 349752 145618 349761
rect 145562 349687 145618 349696
rect 144182 330168 144238 330177
rect 144182 330103 144238 330112
rect 143540 329928 143592 329934
rect 143540 329870 143592 329876
rect 139412 327542 139656 327570
rect 140392 327542 140728 327570
rect 141128 327542 141372 327570
rect 141864 327542 142108 327570
rect 142600 327542 142936 327570
rect 143152 327542 143488 327570
rect 123574 327448 123630 327457
rect 122944 327406 123574 327434
rect 123574 327383 123630 327392
rect 122838 327312 122894 327321
rect 122838 327247 122894 327256
rect 123666 327312 123722 327321
rect 123722 327270 124016 327298
rect 123666 327247 123722 327256
rect 135548 327146 135576 327542
rect 135536 327140 135588 327146
rect 135536 327082 135588 327088
rect 143552 327078 143580 329870
rect 144196 327570 144224 330103
rect 144828 328500 144880 328506
rect 144828 328442 144880 328448
rect 144840 327570 144868 328442
rect 143888 327542 144224 327570
rect 144624 327542 144868 327570
rect 144932 327570 144960 349687
rect 146312 345014 146340 351970
rect 146312 344986 146432 345014
rect 146206 327720 146262 327729
rect 146206 327655 146262 327664
rect 146220 327570 146248 327655
rect 144932 327542 145360 327570
rect 146096 327542 146248 327570
rect 146404 327570 146432 344986
rect 148416 338224 148468 338230
rect 148416 338166 148468 338172
rect 147588 329996 147640 330002
rect 147588 329938 147640 329944
rect 147600 327706 147628 329938
rect 147554 327678 147628 327706
rect 146404 327542 146832 327570
rect 147554 327556 147582 327678
rect 148428 327570 148456 338166
rect 150348 329112 150400 329118
rect 150348 329054 150400 329060
rect 150360 327706 150388 329054
rect 150314 327678 150388 327706
rect 148428 327542 148856 327570
rect 150314 327556 150342 327678
rect 149886 327448 149942 327457
rect 149592 327406 149886 327434
rect 149886 327383 149942 327392
rect 148304 327282 148640 327298
rect 148304 327276 148652 327282
rect 148304 327270 148600 327276
rect 148600 327218 148652 327224
rect 150714 327176 150770 327185
rect 151188 327162 151216 357303
rect 152476 347138 152504 455398
rect 158720 454096 158772 454102
rect 158720 454038 158772 454044
rect 155224 445800 155276 445806
rect 155224 445742 155276 445748
rect 155236 356046 155264 445742
rect 157984 438184 158036 438190
rect 157984 438126 158036 438132
rect 157338 364984 157394 364993
rect 157338 364919 157394 364928
rect 155224 356040 155276 356046
rect 155224 355982 155276 355988
rect 155960 356040 156012 356046
rect 155960 355982 156012 355988
rect 155316 355360 155368 355366
rect 155316 355302 155368 355308
rect 152464 347132 152516 347138
rect 152464 347074 152516 347080
rect 153842 345672 153898 345681
rect 153842 345607 153898 345616
rect 153856 335354 153884 345607
rect 155224 338224 155276 338230
rect 155224 338166 155276 338172
rect 153580 335326 153884 335354
rect 153580 331214 153608 335326
rect 153304 331186 153608 331214
rect 153304 329866 153332 331186
rect 153292 329860 153344 329866
rect 153292 329802 153344 329808
rect 153304 327842 153332 329802
rect 153382 328808 153438 328817
rect 153382 328743 153438 328752
rect 153258 327814 153332 327842
rect 153258 327556 153286 327814
rect 152924 327276 152976 327282
rect 152924 327218 152976 327224
rect 152096 327208 152148 327214
rect 150770 327134 151216 327162
rect 151800 327156 152096 327162
rect 152830 327176 152886 327185
rect 151800 327150 152148 327156
rect 151800 327134 152136 327150
rect 152536 327134 152830 327162
rect 150714 327111 150770 327120
rect 152830 327111 152886 327120
rect 93860 327072 93912 327078
rect 93860 327014 93912 327020
rect 143540 327072 143592 327078
rect 143540 327014 143592 327020
rect 71044 327004 71096 327010
rect 71044 326946 71096 326952
rect 152936 326942 152964 327218
rect 153396 327049 153424 328743
rect 155236 327729 155264 338166
rect 155222 327720 155278 327729
rect 155222 327655 155278 327664
rect 154856 327072 154908 327078
rect 153382 327040 153438 327049
rect 154856 327014 154908 327020
rect 153382 326975 153438 326984
rect 152924 326936 152976 326942
rect 70964 326862 71208 326890
rect 154304 326936 154356 326942
rect 152924 326878 152976 326884
rect 154008 326884 154304 326890
rect 154868 326913 154896 327014
rect 155224 326936 155276 326942
rect 154854 326904 154910 326913
rect 154008 326878 154356 326884
rect 154008 326862 154344 326878
rect 154560 326862 154712 326890
rect 67822 321600 67878 321609
rect 67822 321535 67878 321544
rect 154684 318345 154712 326862
rect 155224 326878 155276 326884
rect 154854 326839 154910 326848
rect 154670 318336 154726 318345
rect 154670 318271 154726 318280
rect 67730 306912 67786 306921
rect 67730 306847 67786 306856
rect 155236 298858 155264 326878
rect 155224 298852 155276 298858
rect 155224 298794 155276 298800
rect 155224 296064 155276 296070
rect 155224 296006 155276 296012
rect 67640 269068 67692 269074
rect 67640 269010 67692 269016
rect 67652 268841 67680 269010
rect 67638 268832 67694 268841
rect 67638 268767 67694 268776
rect 155236 264217 155264 296006
rect 155328 279313 155356 355302
rect 155406 332888 155462 332897
rect 155406 332823 155462 332832
rect 155420 305697 155448 332823
rect 155972 318073 156000 355982
rect 156694 353968 156750 353977
rect 156694 353903 156750 353912
rect 156052 349852 156104 349858
rect 156052 349794 156104 349800
rect 156064 331214 156092 349794
rect 156064 331186 156184 331214
rect 156050 326496 156106 326505
rect 156050 326431 156106 326440
rect 156064 326058 156092 326431
rect 156052 326052 156104 326058
rect 156052 325994 156104 326000
rect 156156 325417 156184 331186
rect 156142 325408 156198 325417
rect 156142 325343 156198 325352
rect 156156 325038 156184 325343
rect 156144 325032 156196 325038
rect 156144 324974 156196 324980
rect 156050 324320 156106 324329
rect 156050 324255 156106 324264
rect 156064 322998 156092 324255
rect 156052 322992 156104 322998
rect 156052 322934 156104 322940
rect 156050 322144 156106 322153
rect 156050 322079 156106 322088
rect 156064 321638 156092 322079
rect 156052 321632 156104 321638
rect 156052 321574 156104 321580
rect 155958 318064 156014 318073
rect 155958 317999 156014 318008
rect 156602 318064 156658 318073
rect 156602 317999 156658 318008
rect 155406 305688 155462 305697
rect 155406 305623 155462 305632
rect 156050 304192 156106 304201
rect 156050 304127 156106 304136
rect 156064 303686 156092 304127
rect 156052 303680 156104 303686
rect 156052 303622 156104 303628
rect 156418 297936 156474 297945
rect 156418 297871 156474 297880
rect 156432 296002 156460 297871
rect 156420 295996 156472 296002
rect 156420 295938 156472 295944
rect 156328 295316 156380 295322
rect 156328 295258 156380 295264
rect 156340 294681 156368 295258
rect 156326 294672 156382 294681
rect 156326 294607 156382 294616
rect 156510 293584 156566 293593
rect 156510 293519 156566 293528
rect 156524 292670 156552 293519
rect 156512 292664 156564 292670
rect 156512 292606 156564 292612
rect 156050 291680 156106 291689
rect 156050 291615 156106 291624
rect 156064 291242 156092 291615
rect 156052 291236 156104 291242
rect 156052 291178 156104 291184
rect 156418 285152 156474 285161
rect 156418 285087 156474 285096
rect 156432 284374 156460 285087
rect 156420 284368 156472 284374
rect 156420 284310 156472 284316
rect 155314 279304 155370 279313
rect 155314 279239 155370 279248
rect 155328 276729 155356 279239
rect 155314 276720 155370 276729
rect 155314 276655 155370 276664
rect 155316 276616 155368 276622
rect 155316 276558 155368 276564
rect 155222 264208 155278 264217
rect 155222 264143 155278 264152
rect 67822 260400 67878 260409
rect 67822 260335 67878 260344
rect 67730 250880 67786 250889
rect 67730 250815 67786 250824
rect 67638 245712 67694 245721
rect 67638 245647 67694 245656
rect 67548 240100 67600 240106
rect 67548 240042 67600 240048
rect 67362 236600 67418 236609
rect 67362 236535 67418 236544
rect 67270 215928 67326 215937
rect 67270 215863 67326 215872
rect 67652 209098 67680 245647
rect 67744 218006 67772 250815
rect 67836 240174 67864 260335
rect 155224 256012 155276 256018
rect 155224 255954 155276 255960
rect 154948 243568 155000 243574
rect 154948 243510 155000 243516
rect 154960 243273 154988 243510
rect 154946 243264 155002 243273
rect 154946 243199 155002 243208
rect 82820 242072 82872 242078
rect 152464 242072 152516 242078
rect 135994 242040 136050 242049
rect 82820 242014 82872 242020
rect 70306 241904 70362 241913
rect 70362 241874 70440 241890
rect 70362 241868 70452 241874
rect 70362 241862 70400 241868
rect 70306 241839 70362 241848
rect 70400 241810 70452 241816
rect 71044 241868 71096 241874
rect 71044 241810 71096 241816
rect 69662 241768 69718 241777
rect 69662 241703 69718 241712
rect 67928 241590 68816 241618
rect 69032 241590 69368 241618
rect 67824 240168 67876 240174
rect 67824 240110 67876 240116
rect 67928 238066 67956 241590
rect 67916 238060 67968 238066
rect 67916 238002 67968 238008
rect 67732 218000 67784 218006
rect 67732 217942 67784 217948
rect 69032 211138 69060 241590
rect 69020 211132 69072 211138
rect 69020 211074 69072 211080
rect 67640 209092 67692 209098
rect 67640 209034 67692 209040
rect 67086 200696 67142 200705
rect 67086 200631 67142 200640
rect 69676 190466 69704 241703
rect 70104 241590 70348 241618
rect 70320 240106 70348 241590
rect 70412 241590 70840 241618
rect 69756 240100 69808 240106
rect 69756 240042 69808 240048
rect 70308 240100 70360 240106
rect 70308 240042 70360 240048
rect 69768 215257 69796 240042
rect 69754 215248 69810 215257
rect 69754 215183 69810 215192
rect 70412 204270 70440 241590
rect 71056 212498 71084 241810
rect 71576 241590 71728 241618
rect 72312 241590 72924 241618
rect 73048 241590 73108 241618
rect 71700 239426 71728 241590
rect 71688 239420 71740 239426
rect 71688 239362 71740 239368
rect 72896 238754 72924 241590
rect 72896 238726 73016 238754
rect 72988 230353 73016 238726
rect 72974 230344 73030 230353
rect 72974 230279 73030 230288
rect 71044 212492 71096 212498
rect 71044 212434 71096 212440
rect 70400 204264 70452 204270
rect 70400 204206 70452 204212
rect 73080 197985 73108 241590
rect 73172 241590 73784 241618
rect 74520 241590 74580 241618
rect 75072 241590 75408 241618
rect 73172 238241 73200 241590
rect 73158 238232 73214 238241
rect 73158 238167 73214 238176
rect 73804 238128 73856 238134
rect 73804 238070 73856 238076
rect 73816 220697 73844 238070
rect 73802 220688 73858 220697
rect 73802 220623 73858 220632
rect 74552 204202 74580 241590
rect 75380 240961 75408 241590
rect 75472 241590 75808 241618
rect 76544 241590 76880 241618
rect 77280 241590 77340 241618
rect 75366 240952 75422 240961
rect 75366 240887 75422 240896
rect 75472 240009 75500 241590
rect 76656 240780 76708 240786
rect 76656 240722 76708 240728
rect 76564 240168 76616 240174
rect 76564 240110 76616 240116
rect 74722 240000 74778 240009
rect 74722 239935 74778 239944
rect 75458 240000 75514 240009
rect 75458 239935 75514 239944
rect 74736 232937 74764 239935
rect 75090 237960 75146 237969
rect 75090 237895 75146 237904
rect 75104 234569 75132 237895
rect 75090 234560 75146 234569
rect 75090 234495 75146 234504
rect 75184 233912 75236 233918
rect 75184 233854 75236 233860
rect 74722 232928 74778 232937
rect 74722 232863 74778 232872
rect 75196 213926 75224 233854
rect 75184 213920 75236 213926
rect 75184 213862 75236 213868
rect 76576 209681 76604 240110
rect 76668 224942 76696 240722
rect 76852 238754 76880 241590
rect 77312 240145 77340 241590
rect 77404 241590 78016 241618
rect 78752 241590 79088 241618
rect 79488 241590 80008 241618
rect 80224 241590 80560 241618
rect 80776 241590 81296 241618
rect 81512 241590 81572 241618
rect 77298 240136 77354 240145
rect 77298 240071 77354 240080
rect 76852 238726 77248 238754
rect 76656 224936 76708 224942
rect 76656 224878 76708 224884
rect 77220 222873 77248 238726
rect 77404 231130 77432 241590
rect 77942 240136 77998 240145
rect 77942 240071 77998 240080
rect 77392 231124 77444 231130
rect 77392 231066 77444 231072
rect 77206 222864 77262 222873
rect 77206 222799 77262 222808
rect 76562 209672 76618 209681
rect 76562 209607 76618 209616
rect 74540 204196 74592 204202
rect 74540 204138 74592 204144
rect 73066 197976 73122 197985
rect 73066 197911 73122 197920
rect 77956 197305 77984 240071
rect 79060 240038 79088 241590
rect 79048 240032 79100 240038
rect 79048 239974 79100 239980
rect 79876 240032 79928 240038
rect 79876 239974 79928 239980
rect 79324 239420 79376 239426
rect 79324 239362 79376 239368
rect 79336 228721 79364 239362
rect 79322 228712 79378 228721
rect 79322 228647 79378 228656
rect 79888 206281 79916 239974
rect 79874 206272 79930 206281
rect 79874 206207 79930 206216
rect 77942 197296 77998 197305
rect 77942 197231 77998 197240
rect 79980 195906 80008 241590
rect 80532 240038 80560 241590
rect 80520 240032 80572 240038
rect 80520 239974 80572 239980
rect 81268 211993 81296 241590
rect 81544 240038 81572 241590
rect 81636 241590 82248 241618
rect 81348 240032 81400 240038
rect 81348 239974 81400 239980
rect 81532 240032 81584 240038
rect 81532 239974 81584 239980
rect 81254 211984 81310 211993
rect 81254 211919 81310 211928
rect 81360 205630 81388 239974
rect 81636 216646 81664 241590
rect 82832 240786 82860 242014
rect 135272 241998 135994 242026
rect 82970 241505 82998 241604
rect 83720 241590 84056 241618
rect 82956 241496 83012 241505
rect 82956 241431 83012 241440
rect 82820 240780 82872 240786
rect 82820 240722 82872 240728
rect 82728 240032 82780 240038
rect 82728 239974 82780 239980
rect 82740 218793 82768 239974
rect 84028 239873 84056 241590
rect 84212 241590 84456 241618
rect 85192 241590 85528 241618
rect 85928 241590 86080 241618
rect 84106 241496 84162 241505
rect 84106 241431 84162 241440
rect 84014 239864 84070 239873
rect 84014 239799 84070 239808
rect 84120 224777 84148 241431
rect 84212 237726 84240 241590
rect 84200 237720 84252 237726
rect 84200 237662 84252 237668
rect 84106 224768 84162 224777
rect 84106 224703 84162 224712
rect 82726 218784 82782 218793
rect 82726 218719 82782 218728
rect 81624 216640 81676 216646
rect 81624 216582 81676 216588
rect 81348 205624 81400 205630
rect 81348 205566 81400 205572
rect 79968 195900 80020 195906
rect 79968 195842 80020 195848
rect 85500 192545 85528 241590
rect 86052 240038 86080 241590
rect 86144 241590 86480 241618
rect 86972 241590 87216 241618
rect 87952 241590 88288 241618
rect 88688 241590 89024 241618
rect 89424 241590 89668 241618
rect 90160 241590 90496 241618
rect 90896 241590 91048 241618
rect 86040 240032 86092 240038
rect 86040 239974 86092 239980
rect 86144 238754 86172 241590
rect 86868 240032 86920 240038
rect 86868 239974 86920 239980
rect 85592 238726 86172 238754
rect 85592 208350 85620 238726
rect 86224 236700 86276 236706
rect 86224 236642 86276 236648
rect 86236 226302 86264 236642
rect 86224 226296 86276 226302
rect 86224 226238 86276 226244
rect 85580 208344 85632 208350
rect 85580 208286 85632 208292
rect 86880 194546 86908 239974
rect 86972 222902 87000 241590
rect 86960 222896 87012 222902
rect 86960 222838 87012 222844
rect 88260 210361 88288 241590
rect 88996 239562 89024 241590
rect 88984 239556 89036 239562
rect 88984 239498 89036 239504
rect 89536 239556 89588 239562
rect 89536 239498 89588 239504
rect 88246 210352 88302 210361
rect 88246 210287 88302 210296
rect 89548 196654 89576 239498
rect 89536 196648 89588 196654
rect 89536 196590 89588 196596
rect 86868 194540 86920 194546
rect 86868 194482 86920 194488
rect 85486 192536 85542 192545
rect 85486 192471 85542 192480
rect 69664 190460 69716 190466
rect 69664 190402 69716 190408
rect 89640 189825 89668 241590
rect 90468 240038 90496 241590
rect 90456 240032 90508 240038
rect 90456 239974 90508 239980
rect 90916 240032 90968 240038
rect 90916 239974 90968 239980
rect 90928 220153 90956 239974
rect 90914 220144 90970 220153
rect 90914 220079 90970 220088
rect 89626 189816 89682 189825
rect 89626 189751 89682 189760
rect 91020 185745 91048 241590
rect 91112 241590 91632 241618
rect 92184 241590 92428 241618
rect 91112 236706 91140 241590
rect 91100 236700 91152 236706
rect 91100 236642 91152 236648
rect 92400 213217 92428 241590
rect 92492 241590 92920 241618
rect 93656 241590 93808 241618
rect 92492 234598 92520 241590
rect 93124 237720 93176 237726
rect 93124 237662 93176 237668
rect 92480 234592 92532 234598
rect 92480 234534 92532 234540
rect 92492 233918 92520 234534
rect 92480 233912 92532 233918
rect 92480 233854 92532 233860
rect 92386 213208 92442 213217
rect 92386 213143 92442 213152
rect 93136 206990 93164 237662
rect 93780 214577 93808 241590
rect 93872 241590 94392 241618
rect 95128 241590 95188 241618
rect 93872 222086 93900 241590
rect 93860 222080 93912 222086
rect 93860 222022 93912 222028
rect 93872 217841 93900 222022
rect 93858 217832 93914 217841
rect 93858 217767 93914 217776
rect 93766 214568 93822 214577
rect 93766 214503 93822 214512
rect 95160 211857 95188 241590
rect 95252 241590 95864 241618
rect 96600 241590 96660 241618
rect 97336 241590 97672 241618
rect 97888 241590 97948 241618
rect 98624 241590 99052 241618
rect 99360 241590 99420 241618
rect 95146 211848 95202 211857
rect 95146 211783 95202 211792
rect 93124 206984 93176 206990
rect 93124 206926 93176 206932
rect 95252 204950 95280 241590
rect 96632 238513 96660 241590
rect 97644 239358 97672 241590
rect 97632 239352 97684 239358
rect 97632 239294 97684 239300
rect 96618 238504 96674 238513
rect 96618 238439 96674 238448
rect 95240 204944 95292 204950
rect 95240 204886 95292 204892
rect 97920 191185 97948 241590
rect 99024 238754 99052 241590
rect 99392 239562 99420 241590
rect 99484 241590 100096 241618
rect 100832 241590 101168 241618
rect 101568 241590 101996 241618
rect 99380 239556 99432 239562
rect 99380 239498 99432 239504
rect 99024 238726 99328 238754
rect 97906 191176 97962 191185
rect 97906 191111 97962 191120
rect 99300 188329 99328 238726
rect 99484 222086 99512 241590
rect 101140 239698 101168 241590
rect 101128 239692 101180 239698
rect 101128 239634 101180 239640
rect 100668 239556 100720 239562
rect 100668 239498 100720 239504
rect 99472 222080 99524 222086
rect 99472 222022 99524 222028
rect 100680 215966 100708 239498
rect 101968 221513 101996 241590
rect 102152 241590 102304 241618
rect 103040 241590 103468 241618
rect 102048 239692 102100 239698
rect 102048 239634 102100 239640
rect 101954 221504 102010 221513
rect 101954 221439 102010 221448
rect 100668 215960 100720 215966
rect 100668 215902 100720 215908
rect 102060 210497 102088 239634
rect 102152 235657 102180 241590
rect 102138 235648 102194 235657
rect 102138 235583 102194 235592
rect 102152 234705 102180 235583
rect 102138 234696 102194 234705
rect 102138 234631 102194 234640
rect 102782 234696 102838 234705
rect 102782 234631 102838 234640
rect 102796 228857 102824 234631
rect 102782 228848 102838 228857
rect 102782 228783 102838 228792
rect 102046 210488 102102 210497
rect 102046 210423 102102 210432
rect 103440 209166 103468 241590
rect 103532 241590 103592 241618
rect 103716 241590 104328 241618
rect 105004 241590 105064 241618
rect 105464 241590 105800 241618
rect 106536 241590 106872 241618
rect 107272 241590 107516 241618
rect 103532 237386 103560 241590
rect 103520 237380 103572 237386
rect 103520 237322 103572 237328
rect 103716 235346 103744 241590
rect 104900 240168 104952 240174
rect 104900 240110 104952 240116
rect 104164 239352 104216 239358
rect 104164 239294 104216 239300
rect 103704 235340 103756 235346
rect 103704 235282 103756 235288
rect 103428 209160 103480 209166
rect 103428 209102 103480 209108
rect 104176 198529 104204 239294
rect 104256 236700 104308 236706
rect 104256 236642 104308 236648
rect 104268 212537 104296 236642
rect 104254 212528 104310 212537
rect 104254 212463 104310 212472
rect 104162 198520 104218 198529
rect 104162 198455 104218 198464
rect 104912 191146 104940 240110
rect 105004 220114 105032 241590
rect 105464 240174 105492 241590
rect 105452 240168 105504 240174
rect 105452 240110 105504 240116
rect 106844 239834 106872 241590
rect 106832 239828 106884 239834
rect 106832 239770 106884 239776
rect 104992 220108 105044 220114
rect 104992 220050 105044 220056
rect 107488 195809 107516 241590
rect 107672 241590 108008 241618
rect 108408 241590 108744 241618
rect 109296 241590 109632 241618
rect 110032 241590 110368 241618
rect 110768 241590 111104 241618
rect 111504 241590 111748 241618
rect 112240 241590 112576 241618
rect 112976 241590 113128 241618
rect 113712 241590 114140 241618
rect 114448 241590 114508 241618
rect 115000 241590 115336 241618
rect 115736 241590 115796 241618
rect 107568 239828 107620 239834
rect 107568 239770 107620 239776
rect 107474 195800 107530 195809
rect 107474 195735 107530 195744
rect 107580 193905 107608 239770
rect 107672 238678 107700 241590
rect 108408 239562 108436 241590
rect 109604 239562 109632 241590
rect 107752 239556 107804 239562
rect 107752 239498 107804 239504
rect 108396 239556 108448 239562
rect 108396 239498 108448 239504
rect 109592 239556 109644 239562
rect 109592 239498 109644 239504
rect 110236 239556 110288 239562
rect 110236 239498 110288 239504
rect 107660 238672 107712 238678
rect 107660 238614 107712 238620
rect 107764 232558 107792 239498
rect 108304 238060 108356 238066
rect 108304 238002 108356 238008
rect 107752 232552 107804 232558
rect 107752 232494 107804 232500
rect 108316 216617 108344 238002
rect 108302 216608 108358 216617
rect 108302 216543 108358 216552
rect 110248 206922 110276 239498
rect 110236 206916 110288 206922
rect 110236 206858 110288 206864
rect 110340 198694 110368 241590
rect 111076 239562 111104 241590
rect 111064 239556 111116 239562
rect 111064 239498 111116 239504
rect 111616 239556 111668 239562
rect 111616 239498 111668 239504
rect 111064 233912 111116 233918
rect 111064 233854 111116 233860
rect 110328 198688 110380 198694
rect 110328 198630 110380 198636
rect 107566 193896 107622 193905
rect 107566 193831 107622 193840
rect 111076 193225 111104 233854
rect 111628 218657 111656 239498
rect 111614 218648 111670 218657
rect 111614 218583 111670 218592
rect 111720 214713 111748 241590
rect 112548 240009 112576 241590
rect 112534 240000 112590 240009
rect 112534 239935 112590 239944
rect 111706 214704 111762 214713
rect 111706 214639 111762 214648
rect 113100 207670 113128 241590
rect 114112 238754 114140 241590
rect 114112 238726 114416 238754
rect 114388 231169 114416 238726
rect 114374 231160 114430 231169
rect 114374 231095 114430 231104
rect 113088 207664 113140 207670
rect 113088 207606 113140 207612
rect 114480 204241 114508 241590
rect 115308 239290 115336 241590
rect 115296 239284 115348 239290
rect 115296 239226 115348 239232
rect 115768 227730 115796 241590
rect 115952 241590 116472 241618
rect 117208 241590 117268 241618
rect 117944 241590 118372 241618
rect 118680 241590 118740 241618
rect 115848 240848 115900 240854
rect 115848 240790 115900 240796
rect 115860 240106 115888 240790
rect 115848 240100 115900 240106
rect 115848 240042 115900 240048
rect 115848 239284 115900 239290
rect 115848 239226 115900 239232
rect 115756 227724 115808 227730
rect 115756 227666 115808 227672
rect 115204 227044 115256 227050
rect 115204 226986 115256 226992
rect 114466 204232 114522 204241
rect 114466 204167 114522 204176
rect 111062 193216 111118 193225
rect 115216 193186 115244 226986
rect 115296 214600 115348 214606
rect 115296 214542 115348 214548
rect 115308 205601 115336 214542
rect 115860 209001 115888 239226
rect 115952 235278 115980 241590
rect 117240 240106 117268 241590
rect 117228 240100 117280 240106
rect 117228 240042 117280 240048
rect 118344 238754 118372 241590
rect 118344 238726 118648 238754
rect 115940 235272 115992 235278
rect 115940 235214 115992 235220
rect 115846 208992 115902 209001
rect 115846 208927 115902 208936
rect 115294 205592 115350 205601
rect 115294 205527 115350 205536
rect 118620 199481 118648 238726
rect 118712 237318 118740 241590
rect 119356 241590 119416 241618
rect 120152 241590 120212 241618
rect 118700 237312 118752 237318
rect 118700 237254 118752 237260
rect 119356 235793 119384 241590
rect 120184 239698 120212 241590
rect 120276 241590 120704 241618
rect 121440 241590 121776 241618
rect 122176 241590 122696 241618
rect 120172 239692 120224 239698
rect 120172 239634 120224 239640
rect 120276 238377 120304 241590
rect 121748 240038 121776 241590
rect 121736 240032 121788 240038
rect 121736 239974 121788 239980
rect 121368 239692 121420 239698
rect 121368 239634 121420 239640
rect 120262 238368 120318 238377
rect 120262 238303 120318 238312
rect 119342 235784 119398 235793
rect 119342 235719 119398 235728
rect 119356 201385 119384 235719
rect 119436 235340 119488 235346
rect 119436 235282 119488 235288
rect 119448 227050 119476 235282
rect 119436 227044 119488 227050
rect 119436 226986 119488 226992
rect 119434 225040 119490 225049
rect 119434 224975 119490 224984
rect 119448 202842 119476 224975
rect 121380 202842 121408 239634
rect 122668 217977 122696 241590
rect 122852 241590 122912 241618
rect 123036 241590 123648 241618
rect 124384 241590 124720 241618
rect 125120 241590 125548 241618
rect 125856 241590 126192 241618
rect 126408 241590 126928 241618
rect 127144 241590 127480 241618
rect 127880 241590 128216 241618
rect 128616 241590 128952 241618
rect 129352 241590 129596 241618
rect 130088 241590 130424 241618
rect 130824 241590 131068 241618
rect 131560 241590 131896 241618
rect 132112 241590 132448 241618
rect 132848 241590 133184 241618
rect 133584 241590 133828 241618
rect 134320 241590 134656 241618
rect 122748 240032 122800 240038
rect 122748 239974 122800 239980
rect 122654 217968 122710 217977
rect 122654 217903 122710 217912
rect 122760 213353 122788 239974
rect 122746 213344 122802 213353
rect 122746 213279 122802 213288
rect 122852 208321 122880 241590
rect 122930 240816 122986 240825
rect 122930 240751 122986 240760
rect 122944 234598 122972 240751
rect 122932 234592 122984 234598
rect 122932 234534 122984 234540
rect 123036 229022 123064 241590
rect 124310 240272 124366 240281
rect 124310 240207 124366 240216
rect 124324 233238 124352 240207
rect 124692 239426 124720 241590
rect 124680 239420 124732 239426
rect 124680 239362 124732 239368
rect 125416 239420 125468 239426
rect 125416 239362 125468 239368
rect 124312 233232 124364 233238
rect 124312 233174 124364 233180
rect 123024 229016 123076 229022
rect 123024 228958 123076 228964
rect 125428 222193 125456 239362
rect 125414 222184 125470 222193
rect 125414 222119 125470 222128
rect 122838 208312 122894 208321
rect 122838 208247 122894 208256
rect 119436 202836 119488 202842
rect 119436 202778 119488 202784
rect 121368 202836 121420 202842
rect 121368 202778 121420 202784
rect 125520 202162 125548 241590
rect 126164 239902 126192 241590
rect 126702 240952 126758 240961
rect 126702 240887 126758 240896
rect 126242 240816 126298 240825
rect 126242 240751 126298 240760
rect 126152 239896 126204 239902
rect 126152 239838 126204 239844
rect 126256 231810 126284 240751
rect 126716 233238 126744 240887
rect 126704 233232 126756 233238
rect 126704 233174 126756 233180
rect 126244 231804 126296 231810
rect 126244 231746 126296 231752
rect 126900 214606 126928 241590
rect 127452 240038 127480 241590
rect 127440 240032 127492 240038
rect 127440 239974 127492 239980
rect 128188 231713 128216 241590
rect 128820 240780 128872 240786
rect 128820 240722 128872 240728
rect 128268 240032 128320 240038
rect 128268 239974 128320 239980
rect 128174 231704 128230 231713
rect 128174 231639 128230 231648
rect 128280 219337 128308 239974
rect 128832 235958 128860 240722
rect 128924 239970 128952 241590
rect 128912 239964 128964 239970
rect 128912 239906 128964 239912
rect 128820 235952 128872 235958
rect 128820 235894 128872 235900
rect 129004 232552 129056 232558
rect 129004 232494 129056 232500
rect 129016 227361 129044 232494
rect 129568 230217 129596 241590
rect 129648 239964 129700 239970
rect 129648 239906 129700 239912
rect 129554 230208 129610 230217
rect 129554 230143 129610 230152
rect 129002 227352 129058 227361
rect 129002 227287 129058 227296
rect 128266 219328 128322 219337
rect 128266 219263 128322 219272
rect 126888 214600 126940 214606
rect 126888 214542 126940 214548
rect 125508 202156 125560 202162
rect 125508 202098 125560 202104
rect 119342 201376 119398 201385
rect 119342 201311 119398 201320
rect 129660 200841 129688 239906
rect 130396 239290 130424 241590
rect 130384 239284 130436 239290
rect 130384 239226 130436 239232
rect 130936 239284 130988 239290
rect 130936 239226 130988 239232
rect 130382 233064 130438 233073
rect 130382 232999 130438 233008
rect 130396 227730 130424 232999
rect 130384 227724 130436 227730
rect 130384 227666 130436 227672
rect 129646 200832 129702 200841
rect 129646 200767 129702 200776
rect 118606 199472 118662 199481
rect 118606 199407 118662 199416
rect 130396 195945 130424 227666
rect 130948 217938 130976 239226
rect 130936 217932 130988 217938
rect 130936 217874 130988 217880
rect 131040 200054 131068 241590
rect 131868 240038 131896 241590
rect 131856 240032 131908 240038
rect 131856 239974 131908 239980
rect 132316 240032 132368 240038
rect 132316 239974 132368 239980
rect 132328 224262 132356 239974
rect 132316 224256 132368 224262
rect 132316 224198 132368 224204
rect 132420 205057 132448 241590
rect 133156 239222 133184 241590
rect 133144 239216 133196 239222
rect 133144 239158 133196 239164
rect 133696 239216 133748 239222
rect 133696 239158 133748 239164
rect 133602 236600 133658 236609
rect 133602 236535 133658 236544
rect 133616 234530 133644 236535
rect 133604 234524 133656 234530
rect 133604 234466 133656 234472
rect 133708 209166 133736 239158
rect 133144 209160 133196 209166
rect 133144 209102 133196 209108
rect 133696 209160 133748 209166
rect 133696 209102 133748 209108
rect 132406 205048 132462 205057
rect 132406 204983 132462 204992
rect 131028 200048 131080 200054
rect 131028 199990 131080 199996
rect 130382 195936 130438 195945
rect 130382 195871 130438 195880
rect 111062 193151 111118 193160
rect 115204 193180 115256 193186
rect 115204 193122 115256 193128
rect 104900 191140 104952 191146
rect 104900 191082 104952 191088
rect 133156 191049 133184 209102
rect 133800 206417 133828 241590
rect 134628 239222 134656 241590
rect 134720 241590 135056 241618
rect 134616 239216 134668 239222
rect 134616 239158 134668 239164
rect 134720 238754 134748 241590
rect 135168 239216 135220 239222
rect 135168 239158 135220 239164
rect 133892 238726 134748 238754
rect 133892 213858 133920 238726
rect 135180 227118 135208 239158
rect 135168 227112 135220 227118
rect 135168 227054 135220 227060
rect 135166 225040 135222 225049
rect 135272 225026 135300 241998
rect 138202 242040 138258 242049
rect 135994 241975 136050 241984
rect 138032 241998 138202 242026
rect 136528 241590 136588 241618
rect 135222 224998 135300 225026
rect 135166 224975 135222 224984
rect 133880 213852 133932 213858
rect 133880 213794 133932 213800
rect 133786 206408 133842 206417
rect 133786 206343 133842 206352
rect 135180 198665 135208 224975
rect 136560 222970 136588 241590
rect 136652 241590 137264 241618
rect 137816 241590 137968 241618
rect 136652 235657 136680 241590
rect 137100 237380 137152 237386
rect 137100 237322 137152 237328
rect 137112 237289 137140 237322
rect 137098 237280 137154 237289
rect 137098 237215 137154 237224
rect 137112 236881 137140 237215
rect 137098 236872 137154 236881
rect 137098 236807 137154 236816
rect 136638 235648 136694 235657
rect 136638 235583 136694 235592
rect 136652 234705 136680 235583
rect 137284 235272 137336 235278
rect 137284 235214 137336 235220
rect 136638 234696 136694 234705
rect 136638 234631 136694 234640
rect 136548 222964 136600 222970
rect 136548 222906 136600 222912
rect 137296 222057 137324 235214
rect 137374 234696 137430 234705
rect 137374 234631 137430 234640
rect 137388 226302 137416 234631
rect 137376 226296 137428 226302
rect 137376 226238 137428 226244
rect 137466 225584 137522 225593
rect 137466 225519 137522 225528
rect 137282 222048 137338 222057
rect 137282 221983 137338 221992
rect 137480 218006 137508 225519
rect 137940 219366 137968 241590
rect 138032 237386 138060 241998
rect 146758 242040 146814 242049
rect 138258 241998 138552 242026
rect 146464 241998 146758 242026
rect 138202 241975 138258 241984
rect 154120 242072 154172 242078
rect 152464 242014 152516 242020
rect 152554 242040 152610 242049
rect 146758 241975 146814 241984
rect 138952 241590 139288 241618
rect 140024 241590 140544 241618
rect 140760 241590 141096 241618
rect 138952 239970 138980 241590
rect 138112 239964 138164 239970
rect 138112 239906 138164 239912
rect 138940 239964 138992 239970
rect 138940 239906 138992 239912
rect 138020 237380 138072 237386
rect 138020 237322 138072 237328
rect 138124 232558 138152 239906
rect 140516 238754 140544 241590
rect 141068 239154 141096 241590
rect 141482 241466 141510 241604
rect 142232 241590 142292 241618
rect 141470 241460 141522 241466
rect 141470 241402 141522 241408
rect 142264 239970 142292 241590
rect 142356 241590 142968 241618
rect 143704 241590 144040 241618
rect 144256 241590 144868 241618
rect 144992 241590 145328 241618
rect 145728 241590 146248 241618
rect 147200 241590 147628 241618
rect 147936 241590 148272 241618
rect 148672 241590 148916 241618
rect 142252 239964 142304 239970
rect 142252 239906 142304 239912
rect 141056 239148 141108 239154
rect 141056 239090 141108 239096
rect 142068 239148 142120 239154
rect 142068 239090 142120 239096
rect 140516 238726 140728 238754
rect 138112 232552 138164 232558
rect 138112 232494 138164 232500
rect 137928 219360 137980 219366
rect 137928 219302 137980 219308
rect 137468 218000 137520 218006
rect 137468 217942 137520 217948
rect 135166 198656 135222 198665
rect 135166 198591 135222 198600
rect 133788 198008 133840 198014
rect 133788 197950 133840 197956
rect 133800 197334 133828 197950
rect 133788 197328 133840 197334
rect 133788 197270 133840 197276
rect 140700 196625 140728 238726
rect 142080 230382 142108 239090
rect 142356 235793 142384 241590
rect 143356 239964 143408 239970
rect 143356 239906 143408 239912
rect 142342 235784 142398 235793
rect 142342 235719 142398 235728
rect 142068 230376 142120 230382
rect 142068 230318 142120 230324
rect 143368 225622 143396 239906
rect 144012 239154 144040 241590
rect 144000 239148 144052 239154
rect 144000 239090 144052 239096
rect 144736 239148 144788 239154
rect 144736 239090 144788 239096
rect 143446 231160 143502 231169
rect 143446 231095 143502 231104
rect 142896 225616 142948 225622
rect 142896 225558 142948 225564
rect 143356 225616 143408 225622
rect 143356 225558 143408 225564
rect 142908 217326 142936 225558
rect 143356 218748 143408 218754
rect 143356 218690 143408 218696
rect 142896 217320 142948 217326
rect 142896 217262 142948 217268
rect 143368 211041 143396 218690
rect 143354 211032 143410 211041
rect 143354 210967 143410 210976
rect 140686 196616 140742 196625
rect 140686 196551 140742 196560
rect 143460 191826 143488 231095
rect 144748 226302 144776 239090
rect 144736 226296 144788 226302
rect 144736 226238 144788 226244
rect 144840 220794 144868 241590
rect 145300 239970 145328 241590
rect 145930 240408 145986 240417
rect 145930 240343 145986 240352
rect 145288 239964 145340 239970
rect 145288 239906 145340 239912
rect 145944 234598 145972 240343
rect 146024 239964 146076 239970
rect 146024 239906 146076 239912
rect 146036 234598 146064 239906
rect 145932 234592 145984 234598
rect 145932 234534 145984 234540
rect 146024 234592 146076 234598
rect 146024 234534 146076 234540
rect 144828 220788 144880 220794
rect 144828 220730 144880 220736
rect 146220 212430 146248 241590
rect 147600 231742 147628 241590
rect 148244 239834 148272 241590
rect 148232 239828 148284 239834
rect 148232 239770 148284 239776
rect 148888 231810 148916 241590
rect 149152 241596 149204 241602
rect 149408 241590 149560 241618
rect 149152 241538 149204 241544
rect 149058 241496 149114 241505
rect 149058 241431 149060 241440
rect 149112 241431 149114 241440
rect 149060 241402 149112 241408
rect 149164 240825 149192 241538
rect 149150 240816 149206 240825
rect 149532 240786 149560 241590
rect 149624 241590 149960 241618
rect 150452 241590 150696 241618
rect 151432 241590 151768 241618
rect 149150 240751 149206 240760
rect 149520 240780 149572 240786
rect 149520 240722 149572 240728
rect 148968 239828 149020 239834
rect 148968 239770 149020 239776
rect 148876 231804 148928 231810
rect 148876 231746 148928 231752
rect 147588 231736 147640 231742
rect 147588 231678 147640 231684
rect 148508 231124 148560 231130
rect 148508 231066 148560 231072
rect 148520 227118 148548 231066
rect 146760 227112 146812 227118
rect 146760 227054 146812 227060
rect 148508 227112 148560 227118
rect 148508 227054 148560 227060
rect 146772 226137 146800 227054
rect 146758 226128 146814 226137
rect 146758 226063 146814 226072
rect 146208 212424 146260 212430
rect 146208 212366 146260 212372
rect 143448 191820 143500 191826
rect 143448 191762 143500 191768
rect 133142 191040 133198 191049
rect 133142 190975 133198 190984
rect 148980 189961 149008 239770
rect 149624 239154 149652 241590
rect 149060 239148 149112 239154
rect 149060 239090 149112 239096
rect 149612 239148 149664 239154
rect 149612 239090 149664 239096
rect 149072 237289 149100 239090
rect 149058 237280 149114 237289
rect 149058 237215 149114 237224
rect 150452 234433 150480 241590
rect 150438 234424 150494 234433
rect 150438 234359 150494 234368
rect 151082 208992 151138 209001
rect 151082 208927 151138 208936
rect 148966 189952 149022 189961
rect 148966 189887 149022 189896
rect 129648 189100 129700 189106
rect 129648 189042 129700 189048
rect 99286 188320 99342 188329
rect 99286 188255 99342 188264
rect 122748 186448 122800 186454
rect 122748 186390 122800 186396
rect 108948 186380 109000 186386
rect 108948 186322 109000 186328
rect 91006 185736 91062 185745
rect 91006 185671 91062 185680
rect 106188 184952 106240 184958
rect 106188 184894 106240 184900
rect 100666 183696 100722 183705
rect 100666 183631 100722 183640
rect 103428 183660 103480 183666
rect 98918 182200 98974 182209
rect 98918 182135 98974 182144
rect 98932 177585 98960 182135
rect 98918 177576 98974 177585
rect 98918 177511 98974 177520
rect 100680 176769 100708 183631
rect 103428 183602 103480 183608
rect 100758 180976 100814 180985
rect 100758 180911 100814 180920
rect 100772 177585 100800 180911
rect 100758 177576 100814 177585
rect 100758 177511 100814 177520
rect 103440 176769 103468 183602
rect 106200 177585 106228 184894
rect 108960 177585 108988 186322
rect 119526 182336 119582 182345
rect 119526 182271 119582 182280
rect 115846 180840 115902 180849
rect 115846 180775 115902 180784
rect 110234 179480 110290 179489
rect 110234 179415 110290 179424
rect 112260 179444 112312 179450
rect 106186 177576 106242 177585
rect 106186 177511 106242 177520
rect 108946 177576 109002 177585
rect 108946 177511 109002 177520
rect 110248 177041 110276 179415
rect 112260 179386 112312 179392
rect 112272 177041 112300 179386
rect 115860 177585 115888 180775
rect 116952 178084 117004 178090
rect 116952 178026 117004 178032
rect 115846 177576 115902 177585
rect 115846 177511 115902 177520
rect 110234 177032 110290 177041
rect 110234 176967 110290 176976
rect 112258 177032 112314 177041
rect 112258 176967 112314 176976
rect 116964 176769 116992 178026
rect 119540 177585 119568 182271
rect 121000 179512 121052 179518
rect 121000 179454 121052 179460
rect 119526 177576 119582 177585
rect 119526 177511 119582 177520
rect 121012 176769 121040 179454
rect 122760 177585 122788 186390
rect 124128 185020 124180 185026
rect 124128 184962 124180 184968
rect 124140 177585 124168 184962
rect 128268 183592 128320 183598
rect 128268 183534 128320 183540
rect 125968 180940 126020 180946
rect 125968 180882 126020 180888
rect 124496 178152 124548 178158
rect 124496 178094 124548 178100
rect 122746 177576 122802 177585
rect 122746 177511 122802 177520
rect 124126 177576 124182 177585
rect 124126 177511 124182 177520
rect 124508 176769 124536 178094
rect 125980 177585 126008 180882
rect 128280 177585 128308 183534
rect 129660 177585 129688 189042
rect 135168 187740 135220 187746
rect 135168 187682 135220 187688
rect 133144 182300 133196 182306
rect 133144 182242 133196 182248
rect 132408 180872 132460 180878
rect 132408 180814 132460 180820
rect 132420 177585 132448 180814
rect 133156 177585 133184 182242
rect 135180 177585 135208 187682
rect 151096 187105 151124 208927
rect 151740 195265 151768 241590
rect 151832 241590 152168 241618
rect 151832 233073 151860 241590
rect 152476 237318 152504 242014
rect 152610 241998 153056 242026
rect 154120 242014 154172 242020
rect 152554 241975 152610 241984
rect 152464 237312 152516 237318
rect 152464 237254 152516 237260
rect 152464 236700 152516 236706
rect 152464 236642 152516 236648
rect 151818 233064 151874 233073
rect 151818 232999 151874 233008
rect 152476 219337 152504 236642
rect 152462 219328 152518 219337
rect 152462 219263 152518 219272
rect 153028 204105 153056 241998
rect 154026 241632 154082 241641
rect 153640 241590 153976 241618
rect 153948 239154 153976 241590
rect 154026 241567 154028 241576
rect 154080 241567 154082 241576
rect 154028 241538 154080 241544
rect 153936 239148 153988 239154
rect 153936 239090 153988 239096
rect 154132 238754 154160 242014
rect 154376 241590 154436 241618
rect 153856 238726 154160 238754
rect 153856 234297 153884 238726
rect 153842 234288 153898 234297
rect 153842 234223 153898 234232
rect 153108 232552 153160 232558
rect 153108 232494 153160 232500
rect 153014 204096 153070 204105
rect 153014 204031 153070 204040
rect 151726 195256 151782 195265
rect 151726 195191 151782 195200
rect 151082 187096 151138 187105
rect 151082 187031 151138 187040
rect 153120 186969 153148 232494
rect 154408 209137 154436 241590
rect 154488 239148 154540 239154
rect 154488 239090 154540 239096
rect 154394 209128 154450 209137
rect 154394 209063 154450 209072
rect 154500 202201 154528 239090
rect 155236 202842 155264 255954
rect 155328 232558 155356 276558
rect 156512 274644 156564 274650
rect 156512 274586 156564 274592
rect 156524 273737 156552 274586
rect 156510 273728 156566 273737
rect 156510 273663 156566 273672
rect 156420 269068 156472 269074
rect 156420 269010 156472 269016
rect 156432 268297 156460 269010
rect 156418 268288 156474 268297
rect 156418 268223 156474 268232
rect 156326 267472 156382 267481
rect 156326 267407 156382 267416
rect 156340 260166 156368 267407
rect 156418 263120 156474 263129
rect 156418 263055 156474 263064
rect 156432 262342 156460 263055
rect 156420 262336 156472 262342
rect 156420 262278 156472 262284
rect 156328 260160 156380 260166
rect 156328 260102 156380 260108
rect 156510 255776 156566 255785
rect 156510 255711 156566 255720
rect 156524 254590 156552 255711
rect 156512 254584 156564 254590
rect 156512 254526 156564 254532
rect 156510 249520 156566 249529
rect 156510 249455 156566 249464
rect 156524 248470 156552 249455
rect 156512 248464 156564 248470
rect 156512 248406 156564 248412
rect 156236 247716 156288 247722
rect 156236 247658 156288 247664
rect 155684 244316 155736 244322
rect 155684 244258 155736 244264
rect 155406 242992 155462 243001
rect 155406 242927 155462 242936
rect 155316 232552 155368 232558
rect 155316 232494 155368 232500
rect 155420 219434 155448 242927
rect 155696 240854 155724 244258
rect 156050 244080 156106 244089
rect 156050 244015 156106 244024
rect 156064 242962 156092 244015
rect 156052 242956 156104 242962
rect 156052 242898 156104 242904
rect 156248 242185 156276 247658
rect 156234 242176 156290 242185
rect 156234 242111 156290 242120
rect 155684 240848 155736 240854
rect 155684 240790 155736 240796
rect 155500 233164 155552 233170
rect 155500 233106 155552 233112
rect 155512 225593 155540 233106
rect 155498 225584 155554 225593
rect 155498 225519 155554 225528
rect 156616 224641 156644 317999
rect 156708 316062 156736 353903
rect 156970 326904 157026 326913
rect 156970 326839 157026 326848
rect 156984 320890 157012 326839
rect 156972 320884 157024 320890
rect 156972 320826 157024 320832
rect 157248 320000 157300 320006
rect 157246 319968 157248 319977
rect 157300 319968 157302 319977
rect 157246 319903 157302 319912
rect 157246 318880 157302 318889
rect 157246 318815 157248 318824
rect 157300 318815 157302 318824
rect 157248 318786 157300 318792
rect 157246 316976 157302 316985
rect 157352 316962 157380 364919
rect 157302 316934 157380 316962
rect 157246 316911 157302 316920
rect 157260 316742 157288 316911
rect 157248 316736 157300 316742
rect 157248 316678 157300 316684
rect 156696 316056 156748 316062
rect 156696 315998 156748 316004
rect 156708 296857 156736 315998
rect 157248 315988 157300 315994
rect 157248 315930 157300 315936
rect 157154 315888 157210 315897
rect 157154 315823 157210 315832
rect 157168 312594 157196 315823
rect 157260 314809 157288 315930
rect 157246 314800 157302 314809
rect 157246 314735 157302 314744
rect 157246 312624 157302 312633
rect 157156 312588 157208 312594
rect 157246 312559 157302 312568
rect 157156 312530 157208 312536
rect 157260 311914 157288 312559
rect 157248 311908 157300 311914
rect 157248 311850 157300 311856
rect 157246 311536 157302 311545
rect 157246 311471 157302 311480
rect 157260 310554 157288 311471
rect 157248 310548 157300 310554
rect 157248 310490 157300 310496
rect 157246 310448 157302 310457
rect 157246 310383 157302 310392
rect 157154 309632 157210 309641
rect 157154 309567 157210 309576
rect 157168 309194 157196 309567
rect 157260 309233 157288 310383
rect 157246 309224 157302 309233
rect 157156 309188 157208 309194
rect 157246 309159 157302 309168
rect 157156 309130 157208 309136
rect 157248 309120 157300 309126
rect 157248 309062 157300 309068
rect 157260 308553 157288 309062
rect 157246 308544 157302 308553
rect 157246 308479 157302 308488
rect 157246 306368 157302 306377
rect 157246 306303 157248 306312
rect 157300 306303 157302 306312
rect 157248 306274 157300 306280
rect 157246 305280 157302 305289
rect 157246 305215 157248 305224
rect 157300 305215 157302 305224
rect 157248 305186 157300 305192
rect 157246 303104 157302 303113
rect 157246 303039 157302 303048
rect 157260 302258 157288 303039
rect 157248 302252 157300 302258
rect 157248 302194 157300 302200
rect 157248 299192 157300 299198
rect 157248 299134 157300 299140
rect 157260 299033 157288 299134
rect 157246 299024 157302 299033
rect 157246 298959 157302 298968
rect 156694 296848 156750 296857
rect 156694 296783 156750 296792
rect 157246 292768 157302 292777
rect 157246 292703 157302 292712
rect 157260 292602 157288 292703
rect 157248 292596 157300 292602
rect 157248 292538 157300 292544
rect 156786 291136 156842 291145
rect 156786 291071 156842 291080
rect 156800 290193 156828 291071
rect 157246 290592 157302 290601
rect 157246 290527 157302 290536
rect 156786 290184 156842 290193
rect 156786 290119 156842 290128
rect 156694 259856 156750 259865
rect 156694 259791 156750 259800
rect 156602 224632 156658 224641
rect 156602 224567 156658 224576
rect 156616 223009 156644 224567
rect 156602 223000 156658 223009
rect 156602 222935 156658 222944
rect 155408 219428 155460 219434
rect 155408 219370 155460 219376
rect 156602 213888 156658 213897
rect 156602 213823 156658 213832
rect 155224 202836 155276 202842
rect 155224 202778 155276 202784
rect 154486 202192 154542 202201
rect 154486 202127 154542 202136
rect 156616 194177 156644 213823
rect 156708 209001 156736 259791
rect 156800 247353 156828 290119
rect 157260 289882 157288 290527
rect 157248 289876 157300 289882
rect 157248 289818 157300 289824
rect 157246 289504 157302 289513
rect 157246 289439 157302 289448
rect 157260 288522 157288 289439
rect 157248 288516 157300 288522
rect 157248 288458 157300 288464
rect 157246 288416 157302 288425
rect 157246 288351 157302 288360
rect 157260 287094 157288 288351
rect 157248 287088 157300 287094
rect 157248 287030 157300 287036
rect 157062 286240 157118 286249
rect 157062 286175 157118 286184
rect 156880 280832 156932 280838
rect 156880 280774 156932 280780
rect 156892 275913 156920 280774
rect 157076 278118 157104 286175
rect 157154 285560 157210 285569
rect 157154 285495 157210 285504
rect 157168 284345 157196 285495
rect 157154 284336 157210 284345
rect 157154 284271 157210 284280
rect 157246 283248 157302 283257
rect 157246 283183 157248 283192
rect 157300 283183 157302 283192
rect 157248 283154 157300 283160
rect 157248 281512 157300 281518
rect 157248 281454 157300 281460
rect 157260 281081 157288 281454
rect 157246 281072 157302 281081
rect 157246 281007 157302 281016
rect 157246 279984 157302 279993
rect 157302 279942 157380 279970
rect 157246 279919 157302 279928
rect 157248 279540 157300 279546
rect 157248 279482 157300 279488
rect 157260 278905 157288 279482
rect 157246 278896 157302 278905
rect 157246 278831 157302 278840
rect 157064 278112 157116 278118
rect 157064 278054 157116 278060
rect 157246 277808 157302 277817
rect 157246 277743 157302 277752
rect 156878 275904 156934 275913
rect 156878 275839 156934 275848
rect 157260 275330 157288 277743
rect 157352 276758 157380 279942
rect 157340 276752 157392 276758
rect 157340 276694 157392 276700
rect 157248 275324 157300 275330
rect 157248 275266 157300 275272
rect 157246 274816 157302 274825
rect 157246 274751 157302 274760
rect 157260 274718 157288 274751
rect 157248 274712 157300 274718
rect 157248 274654 157300 274660
rect 156970 272640 157026 272649
rect 156970 272575 157026 272584
rect 156984 271182 157012 272575
rect 156972 271176 157024 271182
rect 156972 271118 157024 271124
rect 157246 270464 157302 270473
rect 157246 270399 157302 270408
rect 157260 269142 157288 270399
rect 157248 269136 157300 269142
rect 157248 269078 157300 269084
rect 157248 266416 157300 266422
rect 157246 266384 157248 266393
rect 157300 266384 157302 266393
rect 157246 266319 157302 266328
rect 157246 265296 157302 265305
rect 157246 265231 157302 265240
rect 157260 264994 157288 265231
rect 157248 264988 157300 264994
rect 157248 264930 157300 264936
rect 156970 262032 157026 262041
rect 156970 261967 157026 261976
rect 156984 260846 157012 261967
rect 157246 260944 157302 260953
rect 157246 260879 157248 260888
rect 157300 260879 157302 260888
rect 157248 260850 157300 260856
rect 156972 260840 157024 260846
rect 156972 260782 157024 260788
rect 156880 257984 156932 257990
rect 156878 257952 156880 257961
rect 156932 257952 156934 257961
rect 156878 257887 156934 257896
rect 157248 257372 157300 257378
rect 157248 257314 157300 257320
rect 157260 256873 157288 257314
rect 157246 256864 157302 256873
rect 157246 256799 157302 256808
rect 157246 254688 157302 254697
rect 157246 254623 157248 254632
rect 157300 254623 157302 254632
rect 157248 254594 157300 254600
rect 157248 253632 157300 253638
rect 157246 253600 157248 253609
rect 157300 253600 157302 253609
rect 157246 253535 157302 253544
rect 157154 252512 157210 252521
rect 157154 252447 157210 252456
rect 157168 251258 157196 252447
rect 157246 251424 157302 251433
rect 157246 251359 157302 251368
rect 157260 251326 157288 251359
rect 157248 251320 157300 251326
rect 157248 251262 157300 251268
rect 157156 251252 157208 251258
rect 157156 251194 157208 251200
rect 157246 250608 157302 250617
rect 157246 250543 157302 250552
rect 157260 249830 157288 250543
rect 157248 249824 157300 249830
rect 157248 249766 157300 249772
rect 156972 249416 157024 249422
rect 156972 249358 157024 249364
rect 156984 248441 157012 249358
rect 156970 248432 157026 248441
rect 156970 248367 157026 248376
rect 156786 247344 156842 247353
rect 156786 247279 156842 247288
rect 157246 246256 157302 246265
rect 157246 246191 157302 246200
rect 156786 246120 156842 246129
rect 157260 246090 157288 246191
rect 156786 246055 156842 246064
rect 157248 246084 157300 246090
rect 156800 213897 156828 246055
rect 157248 246026 157300 246032
rect 157996 244390 158024 438126
rect 158074 358184 158130 358193
rect 158074 358119 158130 358128
rect 157984 244384 158036 244390
rect 157984 244326 158036 244332
rect 157338 232928 157394 232937
rect 157338 232863 157394 232872
rect 157352 232558 157380 232863
rect 157340 232552 157392 232558
rect 157340 232494 157392 232500
rect 156786 213888 156842 213897
rect 156786 213823 156842 213832
rect 156694 208992 156750 209001
rect 156694 208927 156750 208936
rect 157338 207088 157394 207097
rect 157338 207023 157394 207032
rect 157352 205630 157380 207023
rect 157340 205624 157392 205630
rect 157340 205566 157392 205572
rect 157996 198529 158024 244326
rect 158088 223145 158116 358119
rect 158168 328500 158220 328506
rect 158168 328442 158220 328448
rect 158180 279682 158208 328442
rect 158168 279676 158220 279682
rect 158168 279618 158220 279624
rect 158732 279546 158760 454038
rect 161572 450016 161624 450022
rect 161572 449958 161624 449964
rect 161478 370696 161534 370705
rect 161478 370631 161534 370640
rect 160098 366344 160154 366353
rect 160098 366279 160154 366288
rect 159638 336968 159694 336977
rect 159638 336903 159694 336912
rect 159548 334008 159600 334014
rect 159548 333950 159600 333956
rect 159364 329860 159416 329866
rect 159364 329802 159416 329808
rect 159376 302841 159404 329802
rect 159456 326052 159508 326058
rect 159456 325994 159508 326000
rect 159468 308417 159496 325994
rect 159560 323678 159588 333950
rect 159652 326466 159680 336903
rect 159640 326460 159692 326466
rect 159640 326402 159692 326408
rect 159548 323672 159600 323678
rect 159548 323614 159600 323620
rect 159454 308408 159510 308417
rect 159454 308343 159510 308352
rect 160112 306338 160140 366279
rect 160742 357368 160798 357377
rect 160742 357303 160798 357312
rect 160756 337385 160784 357303
rect 160742 337376 160798 337385
rect 160742 337311 160798 337320
rect 160926 337104 160982 337113
rect 160926 337039 160982 337048
rect 160742 331392 160798 331401
rect 160742 331327 160798 331336
rect 160100 306332 160152 306338
rect 160100 306274 160152 306280
rect 160112 304298 160140 306274
rect 160100 304292 160152 304298
rect 160100 304234 160152 304240
rect 159362 302832 159418 302841
rect 159362 302767 159418 302776
rect 159362 293176 159418 293185
rect 159362 293111 159418 293120
rect 158720 279540 158772 279546
rect 158720 279482 158772 279488
rect 158168 278044 158220 278050
rect 158168 277986 158220 277992
rect 158180 231742 158208 277986
rect 158718 247208 158774 247217
rect 158718 247143 158774 247152
rect 158260 245676 158312 245682
rect 158260 245618 158312 245624
rect 158272 233170 158300 245618
rect 158732 241641 158760 247143
rect 158718 241632 158774 241641
rect 158718 241567 158774 241576
rect 158260 233164 158312 233170
rect 158260 233106 158312 233112
rect 158168 231736 158220 231742
rect 158168 231678 158220 231684
rect 158260 231124 158312 231130
rect 158260 231066 158312 231072
rect 158074 223136 158130 223145
rect 158074 223071 158130 223080
rect 158272 217841 158300 231066
rect 158718 223136 158774 223145
rect 158718 223071 158774 223080
rect 158258 217832 158314 217841
rect 158258 217767 158314 217776
rect 157982 198520 158038 198529
rect 157982 198455 158038 198464
rect 158732 195809 158760 223071
rect 159376 220697 159404 293111
rect 159548 284436 159600 284442
rect 159548 284378 159600 284384
rect 159454 267064 159510 267073
rect 159454 266999 159510 267008
rect 159468 227361 159496 266999
rect 159560 257990 159588 284378
rect 159640 262268 159692 262274
rect 159640 262210 159692 262216
rect 159548 257984 159600 257990
rect 159548 257926 159600 257932
rect 159652 249422 159680 262210
rect 160756 253230 160784 331327
rect 160836 327208 160888 327214
rect 160836 327150 160888 327156
rect 160848 309806 160876 327150
rect 160940 323610 160968 337039
rect 160928 323604 160980 323610
rect 160928 323546 160980 323552
rect 161020 322992 161072 322998
rect 161020 322934 161072 322940
rect 161032 311166 161060 322934
rect 161020 311160 161072 311166
rect 161020 311102 161072 311108
rect 160836 309800 160888 309806
rect 160836 309742 160888 309748
rect 160834 295352 160890 295361
rect 160834 295287 160890 295296
rect 160848 255921 160876 295287
rect 160928 274780 160980 274786
rect 160928 274722 160980 274728
rect 160834 255912 160890 255921
rect 160834 255847 160890 255856
rect 160744 253224 160796 253230
rect 160744 253166 160796 253172
rect 159640 249416 159692 249422
rect 159640 249358 159692 249364
rect 160836 246084 160888 246090
rect 160836 246026 160888 246032
rect 160742 245168 160798 245177
rect 160742 245103 160798 245112
rect 159454 227352 159510 227361
rect 159454 227287 159510 227296
rect 160008 223576 160060 223582
rect 160008 223518 160060 223524
rect 160020 222970 160048 223518
rect 160008 222964 160060 222970
rect 160008 222906 160060 222912
rect 159362 220688 159418 220697
rect 159362 220623 159418 220632
rect 158718 195800 158774 195809
rect 158718 195735 158774 195744
rect 156602 194168 156658 194177
rect 156602 194103 156658 194112
rect 153106 186960 153162 186969
rect 153106 186895 153162 186904
rect 148232 182232 148284 182238
rect 148232 182174 148284 182180
rect 148244 177585 148272 182174
rect 160020 180033 160048 222906
rect 160756 182889 160784 245103
rect 160848 188465 160876 246026
rect 160940 223582 160968 274722
rect 161020 274712 161072 274718
rect 161020 274654 161072 274660
rect 161032 261594 161060 274654
rect 161020 261588 161072 261594
rect 161020 261530 161072 261536
rect 161018 257272 161074 257281
rect 161018 257207 161074 257216
rect 161032 234598 161060 257207
rect 161492 236706 161520 370631
rect 161584 320006 161612 449958
rect 169024 449200 169076 449206
rect 169024 449142 169076 449148
rect 169668 449200 169720 449206
rect 169668 449142 169720 449148
rect 169036 448594 169064 449142
rect 169024 448588 169076 448594
rect 169024 448530 169076 448536
rect 165620 443692 165672 443698
rect 165620 443634 165672 443640
rect 163504 403640 163556 403646
rect 163504 403582 163556 403588
rect 163516 403034 163544 403582
rect 163504 403028 163556 403034
rect 163504 402970 163556 402976
rect 162124 353388 162176 353394
rect 162124 353330 162176 353336
rect 161664 347132 161716 347138
rect 161664 347074 161716 347080
rect 161572 320000 161624 320006
rect 161572 319942 161624 319948
rect 161676 254658 161704 347074
rect 162136 311137 162164 353330
rect 162216 320000 162268 320006
rect 162216 319942 162268 319948
rect 162122 311128 162178 311137
rect 162122 311063 162178 311072
rect 162124 305244 162176 305250
rect 162124 305186 162176 305192
rect 162136 283626 162164 305186
rect 162228 300150 162256 319942
rect 162216 300144 162268 300150
rect 162216 300086 162268 300092
rect 162124 283620 162176 283626
rect 162124 283562 162176 283568
rect 162768 283212 162820 283218
rect 162768 283154 162820 283160
rect 162780 282198 162808 283154
rect 162768 282192 162820 282198
rect 162768 282134 162820 282140
rect 162216 279676 162268 279682
rect 162216 279618 162268 279624
rect 161664 254652 161716 254658
rect 161664 254594 161716 254600
rect 162124 253972 162176 253978
rect 162124 253914 162176 253920
rect 161480 236700 161532 236706
rect 161480 236642 161532 236648
rect 161020 234592 161072 234598
rect 161020 234534 161072 234540
rect 160928 223576 160980 223582
rect 160928 223518 160980 223524
rect 160834 188456 160890 188465
rect 160834 188391 160890 188400
rect 162136 188358 162164 253914
rect 162228 222970 162256 279618
rect 162768 256760 162820 256766
rect 162768 256702 162820 256708
rect 162676 254652 162728 254658
rect 162676 254594 162728 254600
rect 162688 254561 162716 254594
rect 162674 254552 162730 254561
rect 162674 254487 162730 254496
rect 162780 253638 162808 256702
rect 162768 253632 162820 253638
rect 162768 253574 162820 253580
rect 162766 237008 162822 237017
rect 162766 236943 162822 236952
rect 162780 236706 162808 236943
rect 162768 236700 162820 236706
rect 162768 236642 162820 236648
rect 163516 230353 163544 402970
rect 164884 373312 164936 373318
rect 164884 373254 164936 373260
rect 164240 361684 164292 361690
rect 164240 361626 164292 361632
rect 163688 342372 163740 342378
rect 163688 342314 163740 342320
rect 163594 331528 163650 331537
rect 163594 331463 163650 331472
rect 163608 302938 163636 331463
rect 163700 319433 163728 342314
rect 163686 319424 163742 319433
rect 163686 319359 163742 319368
rect 163596 302932 163648 302938
rect 163596 302874 163648 302880
rect 164146 299432 164202 299441
rect 164146 299367 164202 299376
rect 164160 299198 164188 299367
rect 164148 299192 164200 299198
rect 164148 299134 164200 299140
rect 163596 286340 163648 286346
rect 163596 286282 163648 286288
rect 163608 234433 163636 286282
rect 164252 270502 164280 361626
rect 164896 291281 164924 373254
rect 164974 343904 165030 343913
rect 164974 343839 165030 343848
rect 164988 306950 165016 343839
rect 164976 306944 165028 306950
rect 164976 306886 165028 306892
rect 165528 302252 165580 302258
rect 165528 302194 165580 302200
rect 165540 298790 165568 302194
rect 165528 298784 165580 298790
rect 165528 298726 165580 298732
rect 164976 297356 165028 297362
rect 164976 297298 165028 297304
rect 164882 291272 164938 291281
rect 164882 291207 164938 291216
rect 164896 286385 164924 291207
rect 164882 286376 164938 286385
rect 164882 286311 164938 286320
rect 164882 275360 164938 275369
rect 164882 275295 164938 275304
rect 164240 270496 164292 270502
rect 164240 270438 164292 270444
rect 164252 270298 164280 270438
rect 163688 270292 163740 270298
rect 163688 270234 163740 270240
rect 164240 270292 164292 270298
rect 164240 270234 164292 270240
rect 163700 253978 163728 270234
rect 164240 262200 164292 262206
rect 164240 262142 164292 262148
rect 164252 260914 164280 262142
rect 164240 260908 164292 260914
rect 164240 260850 164292 260856
rect 163688 253972 163740 253978
rect 163688 253914 163740 253920
rect 164148 247104 164200 247110
rect 164148 247046 164200 247052
rect 164160 242282 164188 247046
rect 164252 243574 164280 260850
rect 164240 243568 164292 243574
rect 164240 243510 164292 243516
rect 164148 242276 164200 242282
rect 164148 242218 164200 242224
rect 163688 241528 163740 241534
rect 163688 241470 163740 241476
rect 163594 234424 163650 234433
rect 163594 234359 163650 234368
rect 163502 230344 163558 230353
rect 163502 230279 163558 230288
rect 163700 223553 163728 241470
rect 164896 237386 164924 275295
rect 164988 247722 165016 297298
rect 165068 253972 165120 253978
rect 165068 253914 165120 253920
rect 164976 247716 165028 247722
rect 164976 247658 165028 247664
rect 164976 243568 165028 243574
rect 164976 243510 165028 243516
rect 164884 237380 164936 237386
rect 164884 237322 164936 237328
rect 164988 233889 165016 243510
rect 165080 242078 165108 253914
rect 165068 242072 165120 242078
rect 165068 242014 165120 242020
rect 165632 238754 165660 443634
rect 165712 378820 165764 378826
rect 165712 378762 165764 378768
rect 165724 297401 165752 378762
rect 167000 371884 167052 371890
rect 167000 371826 167052 371832
rect 166264 341012 166316 341018
rect 166264 340954 166316 340960
rect 166276 322250 166304 340954
rect 166906 337376 166962 337385
rect 166906 337311 166962 337320
rect 166920 329186 166948 337311
rect 166908 329180 166960 329186
rect 166908 329122 166960 329128
rect 166354 329080 166410 329089
rect 166354 329015 166410 329024
rect 166264 322244 166316 322250
rect 166264 322186 166316 322192
rect 166368 318170 166396 329015
rect 166448 321632 166500 321638
rect 166448 321574 166500 321580
rect 166356 318164 166408 318170
rect 166356 318106 166408 318112
rect 166356 310548 166408 310554
rect 166356 310490 166408 310496
rect 165710 297392 165766 297401
rect 165710 297327 165712 297336
rect 165764 297327 165766 297336
rect 165712 297298 165764 297304
rect 165724 297267 165752 297298
rect 166264 292664 166316 292670
rect 166264 292606 166316 292612
rect 165540 238726 165660 238754
rect 164974 233880 165030 233889
rect 164974 233815 165030 233824
rect 165540 226137 165568 238726
rect 165526 226128 165582 226137
rect 165526 226063 165582 226072
rect 164884 224256 164936 224262
rect 164884 224198 164936 224204
rect 163686 223544 163742 223553
rect 163686 223479 163742 223488
rect 162216 222964 162268 222970
rect 162216 222906 162268 222912
rect 162306 218784 162362 218793
rect 162306 218719 162362 218728
rect 163042 218784 163098 218793
rect 163042 218719 163098 218728
rect 162320 211070 162348 218719
rect 162308 211064 162360 211070
rect 163056 211041 163084 218719
rect 162308 211006 162360 211012
rect 163042 211032 163098 211041
rect 163042 210967 163098 210976
rect 164896 205630 164924 224198
rect 166276 207641 166304 292606
rect 166368 264246 166396 310490
rect 166460 304201 166488 321574
rect 167012 315994 167040 371826
rect 169206 339824 169262 339833
rect 169206 339759 169262 339768
rect 169024 339584 169076 339590
rect 169024 339526 169076 339532
rect 167000 315988 167052 315994
rect 167000 315930 167052 315936
rect 167012 315314 167040 315930
rect 167000 315308 167052 315314
rect 167000 315250 167052 315256
rect 166446 304192 166502 304201
rect 166446 304127 166502 304136
rect 167644 302252 167696 302258
rect 167644 302194 167696 302200
rect 167656 285569 167684 302194
rect 167642 285560 167698 285569
rect 167642 285495 167698 285504
rect 166448 270564 166500 270570
rect 166448 270506 166500 270512
rect 166356 264240 166408 264246
rect 166356 264182 166408 264188
rect 166460 231810 166488 270506
rect 168380 253224 168432 253230
rect 167642 253192 167698 253201
rect 168380 253166 168432 253172
rect 167642 253127 167698 253136
rect 166448 231804 166500 231810
rect 166448 231746 166500 231752
rect 166460 219434 166488 231746
rect 167656 231130 167684 253127
rect 168392 252618 168420 253166
rect 168380 252612 168432 252618
rect 168380 252554 168432 252560
rect 169036 249082 169064 339526
rect 169114 327312 169170 327321
rect 169114 327247 169170 327256
rect 169128 259418 169156 327247
rect 169220 315353 169248 339759
rect 169206 315344 169262 315353
rect 169206 315279 169262 315288
rect 169206 284472 169262 284481
rect 169206 284407 169262 284416
rect 169116 259412 169168 259418
rect 169116 259354 169168 259360
rect 169024 249076 169076 249082
rect 169024 249018 169076 249024
rect 168380 242208 168432 242214
rect 168380 242150 168432 242156
rect 168392 241505 168420 242150
rect 168378 241496 168434 241505
rect 168378 241431 168434 241440
rect 169220 234569 169248 284407
rect 169576 252612 169628 252618
rect 169576 252554 169628 252560
rect 169206 234560 169262 234569
rect 169206 234495 169262 234504
rect 167644 231124 167696 231130
rect 167644 231066 167696 231072
rect 166368 219406 166488 219434
rect 166262 207632 166318 207641
rect 166262 207567 166318 207576
rect 164884 205624 164936 205630
rect 164884 205566 164936 205572
rect 166264 189100 166316 189106
rect 166264 189042 166316 189048
rect 162124 188352 162176 188358
rect 162124 188294 162176 188300
rect 163504 187740 163556 187746
rect 163504 187682 163556 187688
rect 160742 182880 160798 182889
rect 160742 182815 160798 182824
rect 160006 180024 160062 180033
rect 160006 179959 160062 179968
rect 125966 177576 126022 177585
rect 125966 177511 126022 177520
rect 128266 177576 128322 177585
rect 128266 177511 128322 177520
rect 129646 177576 129702 177585
rect 129646 177511 129702 177520
rect 132406 177576 132462 177585
rect 132406 177511 132462 177520
rect 133142 177576 133198 177585
rect 133142 177511 133198 177520
rect 135166 177576 135222 177585
rect 135166 177511 135222 177520
rect 148230 177576 148286 177585
rect 148230 177511 148286 177520
rect 128176 176792 128228 176798
rect 100666 176760 100722 176769
rect 100666 176695 100722 176704
rect 103426 176760 103482 176769
rect 103426 176695 103482 176704
rect 116950 176760 117006 176769
rect 116950 176695 117006 176704
rect 120998 176760 121054 176769
rect 120998 176695 121054 176704
rect 124494 176760 124550 176769
rect 124494 176695 124550 176704
rect 128174 176760 128176 176769
rect 128228 176760 128230 176769
rect 128174 176695 128230 176704
rect 136086 176760 136142 176769
rect 136086 176695 136088 176704
rect 136140 176695 136142 176704
rect 158994 176760 159050 176769
rect 158994 176695 158996 176704
rect 136088 176666 136140 176672
rect 159048 176695 159050 176704
rect 158996 176666 159048 176672
rect 130752 175976 130804 175982
rect 130752 175918 130804 175924
rect 130764 175681 130792 175918
rect 130750 175672 130806 175681
rect 130750 175607 130806 175616
rect 163516 175234 163544 187682
rect 164884 185020 164936 185026
rect 164884 184962 164936 184968
rect 164516 182300 164568 182306
rect 164516 182242 164568 182248
rect 163504 175228 163556 175234
rect 163504 175170 163556 175176
rect 164528 175166 164556 182242
rect 164896 175273 164924 184962
rect 165528 175976 165580 175982
rect 165528 175918 165580 175924
rect 164882 175264 164938 175273
rect 164882 175199 164938 175208
rect 164516 175160 164568 175166
rect 164516 175102 164568 175108
rect 165540 173874 165568 175918
rect 165528 173868 165580 173874
rect 165528 173810 165580 173816
rect 166276 172514 166304 189042
rect 166368 181393 166396 219406
rect 167644 213988 167696 213994
rect 167644 213930 167696 213936
rect 167656 204202 167684 213930
rect 167644 204196 167696 204202
rect 167644 204138 167696 204144
rect 168380 194540 168432 194546
rect 168380 194482 168432 194488
rect 168392 194449 168420 194482
rect 168378 194440 168434 194449
rect 168378 194375 168434 194384
rect 167642 186960 167698 186969
rect 167642 186895 167698 186904
rect 166354 181384 166410 181393
rect 166354 181319 166410 181328
rect 166538 180976 166594 180985
rect 166538 180911 166594 180920
rect 166448 176792 166500 176798
rect 166448 176734 166500 176740
rect 166354 175536 166410 175545
rect 166354 175471 166410 175480
rect 166264 172508 166316 172514
rect 166264 172450 166316 172456
rect 166368 165578 166396 175471
rect 166460 171086 166488 176734
rect 166448 171080 166500 171086
rect 166448 171022 166500 171028
rect 166356 165572 166408 165578
rect 166356 165514 166408 165520
rect 166552 157350 166580 180911
rect 167656 172446 167684 186895
rect 169024 183660 169076 183666
rect 169024 183602 169076 183608
rect 167828 179512 167880 179518
rect 167828 179454 167880 179460
rect 167644 172440 167696 172446
rect 167644 172382 167696 172388
rect 167734 171592 167790 171601
rect 167734 171527 167790 171536
rect 167748 159050 167776 171527
rect 167840 168366 167868 179454
rect 167828 168360 167880 168366
rect 167828 168302 167880 168308
rect 167736 159044 167788 159050
rect 167736 158986 167788 158992
rect 169036 158710 169064 183602
rect 169114 182336 169170 182345
rect 169114 182271 169170 182280
rect 169128 167006 169156 182271
rect 169588 180130 169616 252554
rect 169680 242214 169708 449142
rect 171140 447160 171192 447166
rect 171140 447102 171192 447108
rect 169760 389224 169812 389230
rect 169760 389166 169812 389172
rect 169772 262206 169800 389166
rect 170404 332716 170456 332722
rect 170404 332658 170456 332664
rect 170416 305658 170444 332658
rect 170404 305652 170456 305658
rect 170404 305594 170456 305600
rect 170496 300960 170548 300966
rect 170496 300902 170548 300908
rect 170404 262336 170456 262342
rect 170404 262278 170456 262284
rect 169760 262200 169812 262206
rect 169760 262142 169812 262148
rect 169760 251320 169812 251326
rect 169760 251262 169812 251268
rect 169668 242208 169720 242214
rect 169668 242150 169720 242156
rect 169576 180124 169628 180130
rect 169576 180066 169628 180072
rect 169206 177032 169262 177041
rect 169206 176967 169262 176976
rect 169116 167000 169168 167006
rect 169116 166942 169168 166948
rect 169220 161430 169248 176967
rect 169298 175264 169354 175273
rect 169298 175199 169354 175208
rect 169312 169726 169340 175199
rect 169300 169720 169352 169726
rect 169300 169662 169352 169668
rect 169208 161424 169260 161430
rect 169208 161366 169260 161372
rect 169208 159044 169260 159050
rect 169208 158986 169260 158992
rect 169024 158704 169076 158710
rect 169024 158646 169076 158652
rect 166540 157344 166592 157350
rect 166540 157286 166592 157292
rect 166264 151836 166316 151842
rect 166264 151778 166316 151784
rect 67454 129296 67510 129305
rect 67454 129231 67510 129240
rect 65338 128072 65394 128081
rect 65338 128007 65394 128016
rect 65352 127129 65380 128007
rect 64786 127120 64842 127129
rect 64786 127055 64842 127064
rect 65338 127120 65394 127129
rect 65338 127055 65394 127064
rect 64694 120184 64750 120193
rect 64694 120119 64750 120128
rect 64708 94518 64736 120119
rect 64696 94512 64748 94518
rect 64696 94454 64748 94460
rect 64800 71738 64828 127055
rect 66166 125216 66222 125225
rect 66166 125151 66222 125160
rect 66074 122632 66130 122641
rect 66074 122567 66130 122576
rect 65890 120864 65946 120873
rect 65890 120799 65946 120808
rect 65904 120193 65932 120799
rect 65890 120184 65946 120193
rect 65890 120119 65946 120128
rect 65982 102368 66038 102377
rect 65982 102303 66038 102312
rect 65996 85513 66024 102303
rect 66088 93129 66116 122567
rect 66074 93120 66130 93129
rect 66074 93055 66130 93064
rect 66180 90370 66208 125151
rect 67362 123584 67418 123593
rect 67362 123519 67418 123528
rect 67270 100736 67326 100745
rect 67270 100671 67326 100680
rect 66168 90364 66220 90370
rect 66168 90306 66220 90312
rect 67284 86873 67312 100671
rect 67376 91798 67404 123519
rect 67468 94586 67496 129231
rect 67546 126304 67602 126313
rect 67546 126239 67602 126248
rect 67456 94580 67508 94586
rect 67456 94522 67508 94528
rect 67364 91792 67416 91798
rect 67364 91734 67416 91740
rect 67560 89010 67588 126239
rect 164976 96008 165028 96014
rect 164976 95950 165028 95956
rect 162122 94888 162178 94897
rect 162122 94823 162178 94832
rect 110142 94752 110198 94761
rect 110142 94687 110198 94696
rect 125414 94752 125470 94761
rect 125414 94687 125470 94696
rect 108304 94580 108356 94586
rect 108304 94522 108356 94528
rect 108118 93528 108174 93537
rect 108118 93463 108174 93472
rect 108132 93158 108160 93463
rect 108120 93152 108172 93158
rect 108120 93094 108172 93100
rect 105728 92540 105780 92546
rect 105728 92482 105780 92488
rect 105740 92449 105768 92482
rect 100022 92440 100078 92449
rect 100022 92375 100078 92384
rect 105726 92440 105782 92449
rect 105726 92375 105782 92384
rect 86498 91760 86554 91769
rect 86498 91695 86554 91704
rect 75274 91216 75330 91225
rect 75274 91151 75330 91160
rect 85486 91216 85542 91225
rect 85486 91151 85542 91160
rect 67548 89004 67600 89010
rect 67548 88946 67600 88952
rect 75288 88233 75316 91151
rect 75274 88224 75330 88233
rect 75274 88159 75330 88168
rect 67270 86864 67326 86873
rect 67270 86799 67326 86808
rect 65982 85504 66038 85513
rect 65982 85439 66038 85448
rect 73066 75304 73122 75313
rect 73066 75239 73122 75248
rect 71042 73944 71098 73953
rect 71042 73879 71098 73888
rect 64788 71732 64840 71738
rect 64788 71674 64840 71680
rect 64786 68368 64842 68377
rect 64786 68303 64842 68312
rect 63406 65512 63462 65521
rect 63406 65447 63462 65456
rect 62028 29640 62080 29646
rect 62028 29582 62080 29588
rect 61948 16546 62068 16574
rect 60648 13116 60700 13122
rect 60648 13058 60700 13064
rect 60660 3534 60688 13058
rect 60830 8936 60886 8945
rect 60830 8871 60886 8880
rect 56048 3528 56100 3534
rect 56048 3470 56100 3476
rect 56508 3528 56560 3534
rect 56508 3470 56560 3476
rect 57244 3528 57296 3534
rect 57244 3470 57296 3476
rect 57888 3528 57940 3534
rect 57888 3470 57940 3476
rect 58440 3528 58492 3534
rect 58440 3470 58492 3476
rect 59176 3528 59228 3534
rect 59176 3470 59228 3476
rect 59636 3528 59688 3534
rect 59636 3470 59688 3476
rect 60648 3528 60700 3534
rect 60648 3470 60700 3476
rect 56060 480 56088 3470
rect 57256 480 57284 3470
rect 58452 480 58480 3470
rect 59648 480 59676 3470
rect 60844 480 60872 8871
rect 62040 480 62068 16546
rect 64800 3602 64828 68303
rect 68926 65648 68982 65657
rect 68926 65583 68982 65592
rect 66168 44940 66220 44946
rect 66168 44882 66220 44888
rect 64328 3596 64380 3602
rect 64328 3538 64380 3544
rect 64788 3596 64840 3602
rect 64788 3538 64840 3544
rect 63224 3528 63276 3534
rect 63224 3470 63276 3476
rect 63236 480 63264 3470
rect 64340 480 64368 3538
rect 66180 3466 66208 44882
rect 66718 7576 66774 7585
rect 66718 7511 66774 7520
rect 65524 3460 65576 3466
rect 65524 3402 65576 3408
rect 66168 3460 66220 3466
rect 66168 3402 66220 3408
rect 65536 480 65564 3402
rect 66732 480 66760 7511
rect 68940 3466 68968 65583
rect 70308 49020 70360 49026
rect 70308 48962 70360 48968
rect 70214 39400 70270 39409
rect 70214 39335 70270 39344
rect 70228 16574 70256 39335
rect 70136 16546 70256 16574
rect 69112 3596 69164 3602
rect 69112 3538 69164 3544
rect 67916 3460 67968 3466
rect 67916 3402 67968 3408
rect 68928 3460 68980 3466
rect 68928 3402 68980 3408
rect 67928 480 67956 3402
rect 69124 480 69152 3538
rect 70136 3482 70164 16546
rect 70320 6914 70348 48962
rect 70228 6886 70348 6914
rect 70228 3602 70256 6886
rect 70216 3596 70268 3602
rect 70216 3538 70268 3544
rect 70136 3454 70348 3482
rect 70320 480 70348 3454
rect 71056 3398 71084 73879
rect 71504 6248 71556 6254
rect 71504 6190 71556 6196
rect 71044 3392 71096 3398
rect 71044 3334 71096 3340
rect 71516 480 71544 6190
rect 73080 3466 73108 75239
rect 75826 64152 75882 64161
rect 75826 64087 75882 64096
rect 73802 4856 73858 4865
rect 73802 4791 73858 4800
rect 72608 3460 72660 3466
rect 72608 3402 72660 3408
rect 73068 3460 73120 3466
rect 73068 3402 73120 3408
rect 72620 480 72648 3402
rect 73816 480 73844 4791
rect 75840 3466 75868 64087
rect 77208 61396 77260 61402
rect 77208 61338 77260 61344
rect 77220 3466 77248 61338
rect 79968 60036 80020 60042
rect 79968 59978 80020 59984
rect 77392 9036 77444 9042
rect 77392 8978 77444 8984
rect 75000 3460 75052 3466
rect 75000 3402 75052 3408
rect 75828 3460 75880 3466
rect 75828 3402 75880 3408
rect 76196 3460 76248 3466
rect 76196 3402 76248 3408
rect 77208 3460 77260 3466
rect 77208 3402 77260 3408
rect 75012 480 75040 3402
rect 76208 480 76236 3402
rect 77404 480 77432 8978
rect 79980 6914 80008 59978
rect 85500 53786 85528 91151
rect 86512 89593 86540 91695
rect 95146 91352 95202 91361
rect 95146 91287 95202 91296
rect 97906 91352 97962 91361
rect 97906 91287 97962 91296
rect 86774 91216 86830 91225
rect 86774 91151 86830 91160
rect 88246 91216 88302 91225
rect 88246 91151 88302 91160
rect 89626 91216 89682 91225
rect 89626 91151 89682 91160
rect 91006 91216 91062 91225
rect 91006 91151 91062 91160
rect 91926 91216 91982 91225
rect 91926 91151 91982 91160
rect 93214 91216 93270 91225
rect 93214 91151 93270 91160
rect 95054 91216 95110 91225
rect 95054 91151 95110 91160
rect 86498 89584 86554 89593
rect 86498 89519 86554 89528
rect 85488 53780 85540 53786
rect 85488 53722 85540 53728
rect 86788 52426 86816 91151
rect 88260 82793 88288 91151
rect 88246 82784 88302 82793
rect 88246 82719 88302 82728
rect 89640 78577 89668 91151
rect 89626 78568 89682 78577
rect 89626 78503 89682 78512
rect 91020 77246 91048 91151
rect 91940 86737 91968 91151
rect 93228 86970 93256 91151
rect 93216 86964 93268 86970
rect 93216 86906 93268 86912
rect 91926 86728 91982 86737
rect 91926 86663 91982 86672
rect 91008 77240 91060 77246
rect 91008 77182 91060 77188
rect 94962 67008 95018 67017
rect 94962 66943 95018 66952
rect 93768 62824 93820 62830
rect 93768 62766 93820 62772
rect 87602 61432 87658 61441
rect 87602 61367 87658 61376
rect 86868 58676 86920 58682
rect 86868 58618 86920 58624
rect 86776 52420 86828 52426
rect 86776 52362 86828 52368
rect 85488 40792 85540 40798
rect 85488 40734 85540 40740
rect 84108 28348 84160 28354
rect 84108 28290 84160 28296
rect 81348 17264 81400 17270
rect 81348 17206 81400 17212
rect 79704 6886 80008 6914
rect 78588 3392 78640 3398
rect 78588 3334 78640 3340
rect 78600 480 78628 3334
rect 79704 480 79732 6886
rect 81360 3466 81388 17206
rect 84120 3466 84148 28290
rect 85500 3466 85528 40734
rect 85670 3496 85726 3505
rect 80888 3460 80940 3466
rect 80888 3402 80940 3408
rect 81348 3460 81400 3466
rect 81348 3402 81400 3408
rect 83280 3460 83332 3466
rect 83280 3402 83332 3408
rect 84108 3460 84160 3466
rect 84108 3402 84160 3408
rect 84476 3460 84528 3466
rect 84476 3402 84528 3408
rect 85488 3460 85540 3466
rect 85670 3431 85726 3440
rect 85488 3402 85540 3408
rect 80900 480 80928 3402
rect 82082 2000 82138 2009
rect 82082 1935 82138 1944
rect 82096 480 82124 1935
rect 83292 480 83320 3402
rect 84488 480 84516 3402
rect 85684 480 85712 3431
rect 86880 480 86908 58618
rect 87616 3398 87644 61367
rect 89626 58576 89682 58585
rect 89626 58511 89682 58520
rect 89640 3466 89668 58511
rect 91008 55888 91060 55894
rect 91008 55830 91060 55836
rect 90364 26920 90416 26926
rect 90364 26862 90416 26868
rect 90376 6914 90404 26862
rect 90284 6886 90404 6914
rect 89168 3460 89220 3466
rect 89168 3402 89220 3408
rect 89628 3460 89680 3466
rect 89628 3402 89680 3408
rect 87604 3392 87656 3398
rect 87604 3334 87656 3340
rect 87972 2100 88024 2106
rect 87972 2042 88024 2048
rect 87984 480 88012 2042
rect 89180 480 89208 3402
rect 90284 2174 90312 6886
rect 91020 3058 91048 55830
rect 92388 21412 92440 21418
rect 92388 21354 92440 21360
rect 92400 3466 92428 21354
rect 93780 3466 93808 62766
rect 91560 3460 91612 3466
rect 91560 3402 91612 3408
rect 92388 3460 92440 3466
rect 92388 3402 92440 3408
rect 92756 3460 92808 3466
rect 92756 3402 92808 3408
rect 93768 3460 93820 3466
rect 93768 3402 93820 3408
rect 90364 3052 90416 3058
rect 90364 2994 90416 3000
rect 91008 3052 91060 3058
rect 91008 2994 91060 3000
rect 90272 2168 90324 2174
rect 90272 2110 90324 2116
rect 90376 480 90404 2994
rect 91572 480 91600 3402
rect 92768 480 92796 3402
rect 94976 2990 95004 66943
rect 95068 51066 95096 91151
rect 95160 81394 95188 91287
rect 96526 91216 96582 91225
rect 96526 91151 96582 91160
rect 97814 91216 97870 91225
rect 97814 91151 97870 91160
rect 96540 84182 96568 91151
rect 96528 84176 96580 84182
rect 96528 84118 96580 84124
rect 97828 84114 97856 91151
rect 97816 84108 97868 84114
rect 97816 84050 97868 84056
rect 95148 81388 95200 81394
rect 95148 81330 95200 81336
rect 97920 80073 97948 91287
rect 99194 91216 99250 91225
rect 99194 91151 99250 91160
rect 97906 80064 97962 80073
rect 97906 79999 97962 80008
rect 99208 57934 99236 91151
rect 100036 91118 100064 92375
rect 106924 91792 106976 91798
rect 104530 91760 104586 91769
rect 106924 91734 106976 91740
rect 104530 91695 104586 91704
rect 101954 91352 102010 91361
rect 101954 91287 102010 91296
rect 100574 91216 100630 91225
rect 100574 91151 100630 91160
rect 100024 91112 100076 91118
rect 100024 91054 100076 91060
rect 100588 82822 100616 91151
rect 101968 85377 101996 91287
rect 102046 91216 102102 91225
rect 102046 91151 102102 91160
rect 103334 91216 103390 91225
rect 103334 91151 103390 91160
rect 101954 85368 102010 85377
rect 101954 85303 102010 85312
rect 100576 82816 100628 82822
rect 100576 82758 100628 82764
rect 102060 70378 102088 91151
rect 102048 70372 102100 70378
rect 102048 70314 102100 70320
rect 103348 64870 103376 91151
rect 104256 91112 104308 91118
rect 104256 91054 104308 91060
rect 104164 90364 104216 90370
rect 104164 90306 104216 90312
rect 104176 73137 104204 90306
rect 104268 75886 104296 91054
rect 104544 89729 104572 91695
rect 104714 91216 104770 91225
rect 104714 91151 104770 91160
rect 105542 91216 105598 91225
rect 105542 91151 105598 91160
rect 104530 89720 104586 89729
rect 104530 89655 104586 89664
rect 104256 75880 104308 75886
rect 104256 75822 104308 75828
rect 104162 73128 104218 73137
rect 104162 73063 104218 73072
rect 104728 66230 104756 91151
rect 105556 85542 105584 91151
rect 105544 85536 105596 85542
rect 105544 85478 105596 85484
rect 106186 76664 106242 76673
rect 106186 76599 106242 76608
rect 104806 71224 104862 71233
rect 104806 71159 104862 71168
rect 104716 66224 104768 66230
rect 104716 66166 104768 66172
rect 103336 64864 103388 64870
rect 103336 64806 103388 64812
rect 99196 57928 99248 57934
rect 99196 57870 99248 57876
rect 100668 57248 100720 57254
rect 100668 57190 100720 57196
rect 97908 54528 97960 54534
rect 97908 54470 97960 54476
rect 95056 51060 95108 51066
rect 95056 51002 95108 51008
rect 96252 11756 96304 11762
rect 96252 11698 96304 11704
rect 95148 4888 95200 4894
rect 95148 4830 95200 4836
rect 93952 2984 94004 2990
rect 93952 2926 94004 2932
rect 94964 2984 95016 2990
rect 94964 2926 95016 2932
rect 93964 480 93992 2926
rect 95160 480 95188 4830
rect 96264 480 96292 11698
rect 97816 8968 97868 8974
rect 97816 8910 97868 8916
rect 97828 3534 97856 8910
rect 97816 3528 97868 3534
rect 97816 3470 97868 3476
rect 97920 3466 97948 54470
rect 98644 46300 98696 46306
rect 98644 46242 98696 46248
rect 98656 9042 98684 46242
rect 99288 38004 99340 38010
rect 99288 37946 99340 37952
rect 98644 9036 98696 9042
rect 98644 8978 98696 8984
rect 99300 3534 99328 37946
rect 100680 3534 100708 57190
rect 102048 53100 102100 53106
rect 102048 53042 102100 53048
rect 102060 3534 102088 53042
rect 103428 18692 103480 18698
rect 103428 18634 103480 18640
rect 103440 6914 103468 18634
rect 104820 6914 104848 71159
rect 103348 6886 103468 6914
rect 104544 6886 104848 6914
rect 98644 3528 98696 3534
rect 98644 3470 98696 3476
rect 99288 3528 99340 3534
rect 99288 3470 99340 3476
rect 99840 3528 99892 3534
rect 99840 3470 99892 3476
rect 100668 3528 100720 3534
rect 100668 3470 100720 3476
rect 101036 3528 101088 3534
rect 101036 3470 101088 3476
rect 102048 3528 102100 3534
rect 102048 3470 102100 3476
rect 97448 3460 97500 3466
rect 97448 3402 97500 3408
rect 97908 3460 97960 3466
rect 97908 3402 97960 3408
rect 97460 480 97488 3402
rect 98656 480 98684 3470
rect 99852 480 99880 3470
rect 101048 480 101076 3470
rect 102232 3460 102284 3466
rect 102232 3402 102284 3408
rect 102244 480 102272 3402
rect 103348 480 103376 6886
rect 104544 480 104572 6886
rect 106200 3534 106228 76599
rect 106936 74497 106964 91734
rect 107566 91216 107622 91225
rect 107566 91151 107622 91160
rect 108026 91216 108082 91225
rect 108026 91151 108082 91160
rect 107580 82754 107608 91151
rect 108040 88097 108068 91151
rect 108026 88088 108082 88097
rect 108026 88023 108082 88032
rect 107568 82748 107620 82754
rect 107568 82690 107620 82696
rect 108316 81433 108344 94522
rect 110156 93906 110184 94687
rect 111064 94512 111116 94518
rect 111064 94454 111116 94460
rect 121458 94480 121514 94489
rect 110144 93900 110196 93906
rect 110144 93842 110196 93848
rect 110326 91352 110382 91361
rect 110326 91287 110382 91296
rect 110234 91216 110290 91225
rect 110234 91151 110290 91160
rect 108302 81424 108358 81433
rect 108302 81359 108358 81368
rect 106922 74488 106978 74497
rect 106922 74423 106978 74432
rect 110248 67590 110276 91151
rect 110236 67584 110288 67590
rect 110236 67526 110288 67532
rect 107568 60104 107620 60110
rect 107568 60046 107620 60052
rect 107580 3534 107608 60046
rect 110340 55214 110368 91287
rect 111076 78441 111104 94454
rect 121458 94415 121514 94424
rect 121472 93158 121500 94415
rect 125428 93974 125456 94687
rect 125416 93968 125468 93974
rect 125416 93910 125468 93916
rect 121734 93528 121790 93537
rect 121734 93463 121790 93472
rect 121748 93158 121776 93463
rect 121460 93152 121512 93158
rect 121460 93094 121512 93100
rect 121736 93152 121788 93158
rect 121736 93094 121788 93100
rect 122102 93120 122158 93129
rect 122102 93055 122158 93064
rect 112444 92540 112496 92546
rect 112444 92482 112496 92488
rect 111614 92440 111670 92449
rect 111614 92375 111670 92384
rect 111628 90982 111656 92375
rect 111706 91216 111762 91225
rect 111706 91151 111762 91160
rect 111616 90976 111668 90982
rect 111616 90918 111668 90924
rect 111062 78432 111118 78441
rect 111062 78367 111118 78376
rect 111720 63510 111748 91151
rect 111708 63504 111760 63510
rect 111708 63446 111760 63452
rect 112456 59362 112484 92482
rect 113454 92440 113510 92449
rect 113454 92375 113510 92384
rect 115478 92440 115534 92449
rect 115478 92375 115534 92384
rect 118054 92440 118110 92449
rect 118054 92375 118110 92384
rect 112626 91760 112682 91769
rect 112626 91695 112682 91704
rect 112640 89457 112668 91695
rect 113362 91216 113418 91225
rect 113362 91151 113418 91160
rect 112626 89448 112682 89457
rect 112626 89383 112682 89392
rect 113376 87961 113404 91151
rect 113468 91050 113496 92375
rect 114282 91216 114338 91225
rect 115492 91186 115520 92375
rect 115570 91760 115626 91769
rect 115570 91695 115626 91704
rect 114282 91151 114338 91160
rect 115480 91180 115532 91186
rect 113456 91044 113508 91050
rect 113456 90986 113508 90992
rect 113362 87952 113418 87961
rect 113362 87887 113418 87896
rect 114296 74458 114324 91151
rect 115480 91122 115532 91128
rect 115584 89690 115612 91695
rect 117134 91352 117190 91361
rect 117134 91287 117190 91296
rect 115662 91216 115718 91225
rect 115662 91151 115718 91160
rect 115572 89684 115624 89690
rect 115572 89626 115624 89632
rect 115204 89004 115256 89010
rect 115204 88946 115256 88952
rect 115216 84017 115244 88946
rect 115202 84008 115258 84017
rect 115202 83943 115258 83952
rect 114284 74452 114336 74458
rect 114284 74394 114336 74400
rect 112444 59356 112496 59362
rect 112444 59298 112496 59304
rect 115676 56574 115704 91151
rect 117042 80880 117098 80889
rect 117042 80815 117098 80824
rect 115664 56568 115716 56574
rect 115664 56510 115716 56516
rect 110328 55208 110380 55214
rect 110328 55150 110380 55156
rect 108946 51912 109002 51921
rect 108946 51847 109002 51856
rect 108960 3534 108988 51847
rect 111708 50380 111760 50386
rect 111708 50322 111760 50328
rect 111616 24132 111668 24138
rect 111616 24074 111668 24080
rect 111628 16574 111656 24074
rect 111536 16546 111656 16574
rect 110328 15904 110380 15910
rect 110328 15846 110380 15852
rect 110340 3534 110368 15846
rect 111536 3534 111564 16546
rect 111720 6914 111748 50322
rect 115848 47660 115900 47666
rect 115848 47602 115900 47608
rect 113088 25560 113140 25566
rect 113088 25502 113140 25508
rect 113100 6914 113128 25502
rect 114468 10396 114520 10402
rect 114468 10338 114520 10344
rect 111628 6886 111748 6914
rect 112824 6886 113128 6914
rect 105728 3528 105780 3534
rect 105728 3470 105780 3476
rect 106188 3528 106240 3534
rect 106188 3470 106240 3476
rect 106924 3528 106976 3534
rect 106924 3470 106976 3476
rect 107568 3528 107620 3534
rect 107568 3470 107620 3476
rect 108120 3528 108172 3534
rect 108120 3470 108172 3476
rect 108948 3528 109000 3534
rect 108948 3470 109000 3476
rect 109316 3528 109368 3534
rect 109316 3470 109368 3476
rect 110328 3528 110380 3534
rect 110328 3470 110380 3476
rect 110512 3528 110564 3534
rect 110512 3470 110564 3476
rect 111524 3528 111576 3534
rect 111524 3470 111576 3476
rect 105740 480 105768 3470
rect 106936 480 106964 3470
rect 108132 480 108160 3470
rect 109328 480 109356 3470
rect 110524 480 110552 3470
rect 111628 480 111656 6886
rect 112824 480 112852 6886
rect 114480 3534 114508 10338
rect 115860 3534 115888 47602
rect 117056 3534 117084 80815
rect 117148 73166 117176 91287
rect 117226 91216 117282 91225
rect 117226 91151 117282 91160
rect 117240 79966 117268 91151
rect 118068 91118 118096 92375
rect 121182 91760 121238 91769
rect 121182 91695 121238 91704
rect 119710 91352 119766 91361
rect 119710 91287 119766 91296
rect 118514 91216 118570 91225
rect 118514 91151 118570 91160
rect 118056 91112 118108 91118
rect 118056 91054 118108 91060
rect 117228 79960 117280 79966
rect 117228 79902 117280 79908
rect 118528 78674 118556 91151
rect 119724 88330 119752 91287
rect 119894 91216 119950 91225
rect 119894 91151 119950 91160
rect 119712 88324 119764 88330
rect 119712 88266 119764 88272
rect 118516 78668 118568 78674
rect 118516 78610 118568 78616
rect 117136 73160 117188 73166
rect 117136 73102 117188 73108
rect 119908 71670 119936 91151
rect 121196 89622 121224 91695
rect 121366 91216 121422 91225
rect 121366 91151 121422 91160
rect 121184 89616 121236 89622
rect 121184 89558 121236 89564
rect 119988 75200 120040 75206
rect 119988 75142 120040 75148
rect 119896 71664 119948 71670
rect 119896 71606 119948 71612
rect 118608 13184 118660 13190
rect 118608 13126 118660 13132
rect 118620 3534 118648 13126
rect 119896 3596 119948 3602
rect 119896 3538 119948 3544
rect 114008 3528 114060 3534
rect 114008 3470 114060 3476
rect 114468 3528 114520 3534
rect 114468 3470 114520 3476
rect 115204 3528 115256 3534
rect 115204 3470 115256 3476
rect 115848 3528 115900 3534
rect 115848 3470 115900 3476
rect 116400 3528 116452 3534
rect 116400 3470 116452 3476
rect 117044 3528 117096 3534
rect 117044 3470 117096 3476
rect 117596 3528 117648 3534
rect 117596 3470 117648 3476
rect 118608 3528 118660 3534
rect 118608 3470 118660 3476
rect 118792 3528 118844 3534
rect 118792 3470 118844 3476
rect 114020 480 114048 3470
rect 115216 480 115244 3470
rect 116412 480 116440 3470
rect 117608 480 117636 3470
rect 118804 480 118832 3470
rect 119908 480 119936 3538
rect 120000 3534 120028 75142
rect 120078 64288 120134 64297
rect 120078 64223 120134 64232
rect 120092 58721 120120 64223
rect 121380 62082 121408 91151
rect 122116 64802 122144 93055
rect 136088 92472 136140 92478
rect 136086 92440 136088 92449
rect 136140 92440 136142 92449
rect 136086 92375 136142 92384
rect 152094 92440 152150 92449
rect 152094 92375 152096 92384
rect 152148 92375 152150 92384
rect 152096 92346 152148 92352
rect 124862 92032 124918 92041
rect 124862 91967 124918 91976
rect 124034 91488 124090 91497
rect 124034 91423 124090 91432
rect 122746 91216 122802 91225
rect 122746 91151 122802 91160
rect 122760 69018 122788 91151
rect 122748 69012 122800 69018
rect 122748 68954 122800 68960
rect 124048 66162 124076 91423
rect 124126 91216 124182 91225
rect 124126 91151 124182 91160
rect 124770 91216 124826 91225
rect 124770 91151 124826 91160
rect 124036 66156 124088 66162
rect 124036 66098 124088 66104
rect 122104 64796 122156 64802
rect 122104 64738 122156 64744
rect 121368 62076 121420 62082
rect 121368 62018 121420 62024
rect 120078 58712 120134 58721
rect 120078 58647 120134 58656
rect 124140 52358 124168 91151
rect 124784 86601 124812 91151
rect 124770 86592 124826 86601
rect 124770 86527 124826 86536
rect 124876 74526 124904 91967
rect 151542 91488 151598 91497
rect 151542 91423 151598 91432
rect 126518 91216 126574 91225
rect 126518 91151 126574 91160
rect 126886 91216 126942 91225
rect 126886 91151 126942 91160
rect 129646 91216 129702 91225
rect 129646 91151 129702 91160
rect 131026 91216 131082 91225
rect 133786 91216 133842 91225
rect 131026 91151 131082 91160
rect 133144 91180 133196 91186
rect 126532 85474 126560 91151
rect 126520 85468 126572 85474
rect 126520 85410 126572 85416
rect 126900 82657 126928 91151
rect 126886 82648 126942 82657
rect 126886 82583 126942 82592
rect 129660 81326 129688 91151
rect 129648 81320 129700 81326
rect 129648 81262 129700 81268
rect 126244 76560 126296 76566
rect 126244 76502 126296 76508
rect 124864 74520 124916 74526
rect 124864 74462 124916 74468
rect 124128 52352 124180 52358
rect 124128 52294 124180 52300
rect 124864 43512 124916 43518
rect 124864 43454 124916 43460
rect 122748 42152 122800 42158
rect 122748 42094 122800 42100
rect 121092 14544 121144 14550
rect 121092 14486 121144 14492
rect 119988 3528 120040 3534
rect 119988 3470 120040 3476
rect 121104 480 121132 14486
rect 122760 3330 122788 42094
rect 124128 32496 124180 32502
rect 124128 32438 124180 32444
rect 123484 22840 123536 22846
rect 123484 22782 123536 22788
rect 123496 6914 123524 22782
rect 123404 6886 123524 6914
rect 123404 3466 123432 6886
rect 124140 3534 124168 32438
rect 123484 3528 123536 3534
rect 123484 3470 123536 3476
rect 124128 3528 124180 3534
rect 124876 3505 124904 43454
rect 126256 3602 126284 76502
rect 131040 70310 131068 91151
rect 133786 91151 133842 91160
rect 134522 91216 134578 91225
rect 134522 91151 134578 91160
rect 133144 91122 133196 91128
rect 131028 70304 131080 70310
rect 131028 70246 131080 70252
rect 130384 68332 130436 68338
rect 130384 68274 130436 68280
rect 126244 3596 126296 3602
rect 126244 3538 126296 3544
rect 130396 3534 130424 68274
rect 133156 67522 133184 91122
rect 133800 80034 133828 91151
rect 134536 85241 134564 91151
rect 135904 91112 135956 91118
rect 135904 91054 135956 91060
rect 134522 85232 134578 85241
rect 134522 85167 134578 85176
rect 135916 84153 135944 91054
rect 151556 86902 151584 91423
rect 151726 91352 151782 91361
rect 151726 91287 151782 91296
rect 151634 91216 151690 91225
rect 151634 91151 151690 91160
rect 151544 86896 151596 86902
rect 151544 86838 151596 86844
rect 135902 84144 135958 84153
rect 135902 84079 135958 84088
rect 133788 80028 133840 80034
rect 133788 79970 133840 79976
rect 151648 78606 151676 91151
rect 151636 78600 151688 78606
rect 151636 78542 151688 78548
rect 151740 73098 151768 91287
rect 162136 73166 162164 94823
rect 162768 93220 162820 93226
rect 162768 93162 162820 93168
rect 162780 92410 162808 93162
rect 162768 92404 162820 92410
rect 162768 92346 162820 92352
rect 164884 91792 164936 91798
rect 164884 91734 164936 91740
rect 164896 74458 164924 91734
rect 164988 85241 165016 95950
rect 165896 95940 165948 95946
rect 165896 95882 165948 95888
rect 165908 89622 165936 95882
rect 165896 89616 165948 89622
rect 165896 89558 165948 89564
rect 165068 87644 165120 87650
rect 165068 87586 165120 87592
rect 164974 85232 165030 85241
rect 164974 85167 165030 85176
rect 165080 78606 165108 87586
rect 166276 86902 166304 151778
rect 169116 150476 169168 150482
rect 169116 150418 169168 150424
rect 166356 147688 166408 147694
rect 166356 147630 166408 147636
rect 166368 92478 166396 147630
rect 167736 137284 167788 137290
rect 167736 137226 167788 137232
rect 167642 135280 167698 135289
rect 167642 135215 167698 135224
rect 166540 105596 166592 105602
rect 166540 105538 166592 105544
rect 166356 92472 166408 92478
rect 166356 92414 166408 92420
rect 166552 92177 166580 105538
rect 167656 93673 167684 135215
rect 167748 108769 167776 137226
rect 169024 134632 169076 134638
rect 169024 134574 169076 134580
rect 168288 111784 168340 111790
rect 168286 111752 168288 111761
rect 168340 111752 168342 111761
rect 168286 111687 168342 111696
rect 167828 110424 167880 110430
rect 167828 110366 167880 110372
rect 167840 110129 167868 110366
rect 167826 110120 167882 110129
rect 167826 110055 167882 110064
rect 167734 108760 167790 108769
rect 167734 108695 167790 108704
rect 167828 106344 167880 106350
rect 167828 106286 167880 106292
rect 167736 100020 167788 100026
rect 167736 99962 167788 99968
rect 167642 93664 167698 93673
rect 167642 93599 167698 93608
rect 166538 92168 166594 92177
rect 166538 92103 166594 92112
rect 166448 91860 166500 91866
rect 166448 91802 166500 91808
rect 166264 86896 166316 86902
rect 166264 86838 166316 86844
rect 165068 78600 165120 78606
rect 165068 78542 165120 78548
rect 164884 74452 164936 74458
rect 164884 74394 164936 74400
rect 162124 73160 162176 73166
rect 162124 73102 162176 73108
rect 151728 73092 151780 73098
rect 151728 73034 151780 73040
rect 166460 67522 166488 91802
rect 167748 71670 167776 99962
rect 167840 86970 167868 106286
rect 167920 98048 167972 98054
rect 167920 97990 167972 97996
rect 167932 89593 167960 97990
rect 167918 89584 167974 89593
rect 167918 89519 167974 89528
rect 169036 87961 169064 134574
rect 169128 111790 169156 150418
rect 169220 150414 169248 158986
rect 169208 150408 169260 150414
rect 169208 150350 169260 150356
rect 169208 125656 169260 125662
rect 169208 125598 169260 125604
rect 169116 111784 169168 111790
rect 169116 111726 169168 111732
rect 169116 99408 169168 99414
rect 169116 99350 169168 99356
rect 169022 87952 169078 87961
rect 169022 87887 169078 87896
rect 167828 86964 167880 86970
rect 167828 86906 167880 86912
rect 169128 82793 169156 99350
rect 169220 93974 169248 125598
rect 169300 120760 169352 120766
rect 169300 120702 169352 120708
rect 169312 94897 169340 120702
rect 169576 97980 169628 97986
rect 169576 97922 169628 97928
rect 169588 96665 169616 97922
rect 169574 96656 169630 96665
rect 169574 96591 169630 96600
rect 169298 94888 169354 94897
rect 169298 94823 169354 94832
rect 169208 93968 169260 93974
rect 169208 93910 169260 93916
rect 169206 93120 169262 93129
rect 169206 93055 169262 93064
rect 169114 82784 169170 82793
rect 169114 82719 169170 82728
rect 169220 78674 169248 93055
rect 169208 78668 169260 78674
rect 169208 78610 169260 78616
rect 167736 71664 167788 71670
rect 167736 71606 167788 71612
rect 169772 68338 169800 251262
rect 170416 145586 170444 262278
rect 170508 229090 170536 300902
rect 170588 278112 170640 278118
rect 170588 278054 170640 278060
rect 170600 250510 170628 278054
rect 170588 250504 170640 250510
rect 170588 250446 170640 250452
rect 170496 229084 170548 229090
rect 170496 229026 170548 229032
rect 171152 222057 171180 447102
rect 191102 445904 191158 445913
rect 191102 445839 191158 445848
rect 186964 438932 187016 438938
rect 186964 438874 187016 438880
rect 172520 422340 172572 422346
rect 172520 422282 172572 422288
rect 171232 367804 171284 367810
rect 171232 367746 171284 367752
rect 171244 299441 171272 367746
rect 171784 334076 171836 334082
rect 171784 334018 171836 334024
rect 171796 319462 171824 334018
rect 171784 319456 171836 319462
rect 171784 319398 171836 319404
rect 172532 309126 172560 422282
rect 180064 396092 180116 396098
rect 180064 396034 180116 396040
rect 172612 392012 172664 392018
rect 172612 391954 172664 391960
rect 172520 309120 172572 309126
rect 172520 309062 172572 309068
rect 171784 306944 171836 306950
rect 171784 306886 171836 306892
rect 171230 299432 171286 299441
rect 171230 299367 171286 299376
rect 171232 288448 171284 288454
rect 171232 288390 171284 288396
rect 171244 280838 171272 288390
rect 171232 280832 171284 280838
rect 171232 280774 171284 280780
rect 171138 222048 171194 222057
rect 171138 221983 171194 221992
rect 171796 202230 171824 306886
rect 172624 306374 172652 391954
rect 177488 382968 177540 382974
rect 177488 382910 177540 382916
rect 175280 381540 175332 381546
rect 175280 381482 175332 381488
rect 174636 369164 174688 369170
rect 174636 369106 174688 369112
rect 173162 360904 173218 360913
rect 173162 360839 173218 360848
rect 173176 306406 173204 360839
rect 174542 330032 174598 330041
rect 174542 329967 174598 329976
rect 173808 309120 173860 309126
rect 173808 309062 173860 309068
rect 173820 308446 173848 309062
rect 173808 308440 173860 308446
rect 173808 308382 173860 308388
rect 173164 306400 173216 306406
rect 172624 306346 172744 306374
rect 172426 299432 172482 299441
rect 172426 299367 172482 299376
rect 172440 298761 172468 299367
rect 172426 298752 172482 298761
rect 172426 298687 172482 298696
rect 172716 295322 172744 306346
rect 173164 306342 173216 306348
rect 172704 295316 172756 295322
rect 172704 295258 172756 295264
rect 171876 279472 171928 279478
rect 171876 279414 171928 279420
rect 171888 232937 171916 279414
rect 171968 264988 172020 264994
rect 171968 264930 172020 264936
rect 171980 246362 172008 264930
rect 172520 248464 172572 248470
rect 172520 248406 172572 248412
rect 171968 246356 172020 246362
rect 171968 246298 172020 246304
rect 172532 243574 172560 248406
rect 172520 243568 172572 243574
rect 172520 243510 172572 243516
rect 171874 232928 171930 232937
rect 171874 232863 171930 232872
rect 173176 232801 173204 306342
rect 173348 298852 173400 298858
rect 173348 298794 173400 298800
rect 173256 275324 173308 275330
rect 173256 275266 173308 275272
rect 173162 232792 173218 232801
rect 173162 232727 173218 232736
rect 173268 228954 173296 275266
rect 173360 261526 173388 298794
rect 173808 295316 173860 295322
rect 173808 295258 173860 295264
rect 173820 294710 173848 295258
rect 173808 294704 173860 294710
rect 173808 294646 173860 294652
rect 173532 266484 173584 266490
rect 173532 266426 173584 266432
rect 173348 261520 173400 261526
rect 173348 261462 173400 261468
rect 173544 233238 173572 266426
rect 173808 254584 173860 254590
rect 173808 254526 173860 254532
rect 173820 251870 173848 254526
rect 173808 251864 173860 251870
rect 173808 251806 173860 251812
rect 173348 233232 173400 233238
rect 173348 233174 173400 233180
rect 173532 233232 173584 233238
rect 173532 233174 173584 233180
rect 173256 228948 173308 228954
rect 173256 228890 173308 228896
rect 173164 215960 173216 215966
rect 173164 215902 173216 215908
rect 171874 205048 171930 205057
rect 171874 204983 171930 204992
rect 171784 202224 171836 202230
rect 171784 202166 171836 202172
rect 170496 180940 170548 180946
rect 170496 180882 170548 180888
rect 170508 171018 170536 180882
rect 171784 179444 171836 179450
rect 171784 179386 171836 179392
rect 170496 171012 170548 171018
rect 170496 170954 170548 170960
rect 171796 164218 171824 179386
rect 171784 164212 171836 164218
rect 171784 164154 171836 164160
rect 171888 159390 171916 204983
rect 173176 203590 173204 215902
rect 173164 203584 173216 203590
rect 173164 203526 173216 203532
rect 173360 198121 173388 233174
rect 173806 233064 173862 233073
rect 173806 232999 173862 233008
rect 173820 232558 173848 232999
rect 173808 232552 173860 232558
rect 173808 232494 173860 232500
rect 173346 198112 173402 198121
rect 173346 198047 173402 198056
rect 171966 175400 172022 175409
rect 171966 175335 172022 175344
rect 171980 162858 172008 175335
rect 171968 162852 172020 162858
rect 171968 162794 172020 162800
rect 171876 159384 171928 159390
rect 171876 159326 171928 159332
rect 170404 145580 170456 145586
rect 170404 145522 170456 145528
rect 170402 140856 170458 140865
rect 170402 140791 170458 140800
rect 170416 93537 170444 140791
rect 173164 138712 173216 138718
rect 173164 138654 173216 138660
rect 171784 129804 171836 129810
rect 171784 129746 171836 129752
rect 170588 117360 170640 117366
rect 170588 117302 170640 117308
rect 170496 110492 170548 110498
rect 170496 110434 170548 110440
rect 170402 93528 170458 93537
rect 170402 93463 170458 93472
rect 170508 75886 170536 110434
rect 170600 90982 170628 117302
rect 170588 90976 170640 90982
rect 170588 90918 170640 90924
rect 171796 85377 171824 129746
rect 171874 116512 171930 116521
rect 171874 116447 171930 116456
rect 171782 85368 171838 85377
rect 171782 85303 171838 85312
rect 171888 82657 171916 116447
rect 171968 102196 172020 102202
rect 171968 102138 172020 102144
rect 171874 82648 171930 82657
rect 171874 82583 171930 82592
rect 170496 75880 170548 75886
rect 170496 75822 170548 75828
rect 171980 74497 172008 102138
rect 171966 74488 172022 74497
rect 171966 74423 172022 74432
rect 173176 70310 173204 138654
rect 173256 127016 173308 127022
rect 173256 126958 173308 126964
rect 173268 91089 173296 126958
rect 173348 109064 173400 109070
rect 173348 109006 173400 109012
rect 173254 91080 173310 91089
rect 173254 91015 173310 91024
rect 173360 84114 173388 109006
rect 173440 102808 173492 102814
rect 173440 102750 173492 102756
rect 173348 84108 173400 84114
rect 173348 84050 173400 84056
rect 173452 79966 173480 102750
rect 173440 79960 173492 79966
rect 173440 79902 173492 79908
rect 174556 77994 174584 329967
rect 174648 291417 174676 369106
rect 175292 296070 175320 381482
rect 177394 346624 177450 346633
rect 177394 346559 177450 346568
rect 176014 342544 176070 342553
rect 176014 342479 176070 342488
rect 175280 296064 175332 296070
rect 175280 296006 175332 296012
rect 174634 291408 174690 291417
rect 174634 291343 174690 291352
rect 174648 264217 174676 291343
rect 174726 287328 174782 287337
rect 174726 287263 174782 287272
rect 174634 264208 174690 264217
rect 174634 264143 174690 264152
rect 174634 262576 174690 262585
rect 174634 262511 174690 262520
rect 174648 195974 174676 262511
rect 174740 243953 174768 287263
rect 175922 270600 175978 270609
rect 175922 270535 175978 270544
rect 174726 243944 174782 243953
rect 174726 243879 174782 243888
rect 174636 195968 174688 195974
rect 174636 195910 174688 195916
rect 174648 188358 174676 195910
rect 174636 188352 174688 188358
rect 174636 188294 174688 188300
rect 174636 186448 174688 186454
rect 174636 186390 174688 186396
rect 174648 168298 174676 186390
rect 174636 168292 174688 168298
rect 174636 168234 174688 168240
rect 174636 122868 174688 122874
rect 174636 122810 174688 122816
rect 174648 93158 174676 122810
rect 174728 104916 174780 104922
rect 174728 104858 174780 104864
rect 174636 93152 174688 93158
rect 174636 93094 174688 93100
rect 174544 77988 174596 77994
rect 174544 77930 174596 77936
rect 174740 77246 174768 104858
rect 175936 82249 175964 270535
rect 176028 236706 176056 342479
rect 177304 329996 177356 330002
rect 177304 329938 177356 329944
rect 176108 302932 176160 302938
rect 176108 302874 176160 302880
rect 176120 302297 176148 302874
rect 176106 302288 176162 302297
rect 176106 302223 176162 302232
rect 176566 302288 176622 302297
rect 176566 302223 176622 302232
rect 176580 273222 176608 302223
rect 176568 273216 176620 273222
rect 176568 273158 176620 273164
rect 176016 236700 176068 236706
rect 176016 236642 176068 236648
rect 176016 124228 176068 124234
rect 176016 124170 176068 124176
rect 175922 82240 175978 82249
rect 175922 82175 175978 82184
rect 174728 77240 174780 77246
rect 174728 77182 174780 77188
rect 173164 70304 173216 70310
rect 173164 70246 173216 70252
rect 169760 68332 169812 68338
rect 169760 68274 169812 68280
rect 133144 67516 133196 67522
rect 133144 67458 133196 67464
rect 166448 67516 166500 67522
rect 166448 67458 166500 67464
rect 160742 67144 160798 67153
rect 160742 67079 160798 67088
rect 135258 43480 135314 43489
rect 135258 43415 135314 43424
rect 135272 14754 135300 43415
rect 160756 22846 160784 67079
rect 176028 52358 176056 124170
rect 176200 113212 176252 113218
rect 176200 113154 176252 113160
rect 176212 90953 176240 113154
rect 176198 90944 176254 90953
rect 176198 90879 176254 90888
rect 176108 90432 176160 90438
rect 176108 90374 176160 90380
rect 176120 67590 176148 90374
rect 176108 67584 176160 67590
rect 176108 67526 176160 67532
rect 176016 52352 176068 52358
rect 176016 52294 176068 52300
rect 160744 22840 160796 22846
rect 160744 22782 160796 22788
rect 135260 14748 135312 14754
rect 135260 14690 135312 14696
rect 136456 14748 136508 14754
rect 136456 14690 136508 14696
rect 132958 13016 133014 13025
rect 132958 12951 133014 12960
rect 129372 3528 129424 3534
rect 124128 3470 124180 3476
rect 124862 3496 124918 3505
rect 123392 3460 123444 3466
rect 123392 3402 123444 3408
rect 122288 3324 122340 3330
rect 122288 3266 122340 3272
rect 122748 3324 122800 3330
rect 122748 3266 122800 3272
rect 122300 480 122328 3266
rect 123496 480 123524 3470
rect 124680 3460 124732 3466
rect 124862 3431 124918 3440
rect 125874 3496 125930 3505
rect 129372 3470 129424 3476
rect 130384 3528 130436 3534
rect 130384 3470 130436 3476
rect 125874 3431 125930 3440
rect 124680 3402 124732 3408
rect 124692 480 124720 3402
rect 125888 480 125916 3431
rect 129384 480 129412 3470
rect 132972 480 133000 12951
rect 136468 480 136496 14690
rect 177316 9042 177344 329938
rect 177408 135930 177436 346559
rect 177500 294001 177528 382910
rect 178684 360324 178736 360330
rect 178684 360266 178736 360272
rect 177580 309188 177632 309194
rect 177580 309130 177632 309136
rect 177592 297537 177620 309130
rect 177578 297528 177634 297537
rect 177578 297463 177634 297472
rect 177486 293992 177542 294001
rect 177486 293927 177542 293936
rect 177500 260846 177528 293927
rect 177580 261588 177632 261594
rect 177580 261530 177632 261536
rect 177488 260840 177540 260846
rect 177488 260782 177540 260788
rect 177592 234598 177620 261530
rect 177948 256760 178000 256766
rect 177948 256702 178000 256708
rect 177580 234592 177632 234598
rect 177580 234534 177632 234540
rect 177960 193866 177988 256702
rect 178696 256222 178724 360266
rect 178774 341184 178830 341193
rect 178774 341119 178830 341128
rect 178788 330546 178816 341119
rect 178776 330540 178828 330546
rect 178776 330482 178828 330488
rect 179420 329180 179472 329186
rect 179420 329122 179472 329128
rect 179432 327758 179460 329122
rect 179420 327752 179472 327758
rect 179420 327694 179472 327700
rect 178868 318844 178920 318850
rect 178868 318786 178920 318792
rect 178880 315314 178908 318786
rect 178776 315308 178828 315314
rect 178776 315250 178828 315256
rect 178868 315308 178920 315314
rect 178868 315250 178920 315256
rect 178788 269006 178816 315250
rect 178866 285832 178922 285841
rect 178866 285767 178922 285776
rect 178776 269000 178828 269006
rect 178776 268942 178828 268948
rect 178684 256216 178736 256222
rect 178684 256158 178736 256164
rect 178682 254552 178738 254561
rect 178682 254487 178738 254496
rect 178696 235793 178724 254487
rect 178880 240281 178908 285767
rect 178960 269136 179012 269142
rect 178960 269078 179012 269084
rect 178972 259486 179000 269078
rect 180076 268394 180104 396034
rect 185584 376780 185636 376786
rect 185584 376722 185636 376728
rect 182824 368552 182876 368558
rect 182824 368494 182876 368500
rect 181536 358896 181588 358902
rect 181536 358838 181588 358844
rect 180154 347984 180210 347993
rect 180154 347919 180210 347928
rect 180064 268388 180116 268394
rect 180064 268330 180116 268336
rect 179052 260160 179104 260166
rect 179052 260102 179104 260108
rect 178960 259480 179012 259486
rect 178960 259422 179012 259428
rect 178958 249928 179014 249937
rect 178958 249863 179014 249872
rect 178866 240272 178922 240281
rect 178866 240207 178922 240216
rect 178880 238754 178908 240207
rect 178788 238726 178908 238754
rect 178682 235784 178738 235793
rect 178682 235719 178738 235728
rect 178682 209128 178738 209137
rect 178682 209063 178738 209072
rect 177948 193860 178000 193866
rect 177948 193802 178000 193808
rect 177486 178256 177542 178265
rect 177486 178191 177542 178200
rect 177500 164150 177528 178191
rect 177488 164144 177540 164150
rect 177488 164086 177540 164092
rect 177488 143608 177540 143614
rect 177488 143550 177540 143556
rect 177396 135924 177448 135930
rect 177396 135866 177448 135872
rect 177396 134564 177448 134570
rect 177396 134506 177448 134512
rect 177408 93226 177436 134506
rect 177396 93220 177448 93226
rect 177396 93162 177448 93168
rect 177500 81326 177528 143550
rect 177580 100768 177632 100774
rect 177580 100710 177632 100716
rect 177488 81320 177540 81326
rect 177488 81262 177540 81268
rect 177592 78441 177620 100710
rect 178696 83502 178724 209063
rect 178788 175273 178816 238726
rect 178972 236881 179000 249863
rect 179064 241505 179092 260102
rect 180076 257281 180104 268330
rect 180062 257272 180118 257281
rect 180062 257207 180118 257216
rect 180064 251252 180116 251258
rect 180064 251194 180116 251200
rect 179050 241496 179106 241505
rect 179050 241431 179106 241440
rect 178958 236872 179014 236881
rect 178958 236807 179014 236816
rect 180076 216578 180104 251194
rect 180064 216572 180116 216578
rect 180064 216514 180116 216520
rect 180062 213344 180118 213353
rect 180062 213279 180118 213288
rect 179328 191752 179380 191758
rect 179328 191694 179380 191700
rect 179340 191146 179368 191694
rect 179328 191140 179380 191146
rect 179328 191082 179380 191088
rect 179340 182850 179368 191082
rect 179328 182844 179380 182850
rect 179328 182786 179380 182792
rect 178866 182200 178922 182209
rect 178866 182135 178922 182144
rect 178774 175264 178830 175273
rect 178774 175199 178830 175208
rect 178880 155922 178908 182135
rect 178868 155916 178920 155922
rect 178868 155858 178920 155864
rect 178868 136672 178920 136678
rect 178868 136614 178920 136620
rect 178776 128376 178828 128382
rect 178776 128318 178828 128324
rect 178684 83496 178736 83502
rect 178684 83438 178736 83444
rect 177578 78432 177634 78441
rect 177578 78367 177634 78376
rect 178788 57934 178816 128318
rect 178880 91866 178908 136614
rect 178960 121508 179012 121514
rect 178960 121450 179012 121456
rect 178972 93129 179000 121450
rect 179052 93220 179104 93226
rect 179052 93162 179104 93168
rect 178958 93120 179014 93129
rect 178958 93055 179014 93064
rect 178868 91860 178920 91866
rect 178868 91802 178920 91808
rect 179064 70378 179092 93162
rect 179052 70372 179104 70378
rect 179052 70314 179104 70320
rect 178776 57928 178828 57934
rect 178776 57870 178828 57876
rect 180076 46209 180104 213279
rect 180168 184210 180196 347919
rect 180246 327584 180302 327593
rect 180246 327519 180302 327528
rect 180260 283257 180288 327519
rect 181442 324456 181498 324465
rect 181442 324391 181498 324400
rect 180340 287156 180392 287162
rect 180340 287098 180392 287104
rect 180246 283248 180302 283257
rect 180246 283183 180302 283192
rect 180248 278112 180300 278118
rect 180248 278054 180300 278060
rect 180260 191758 180288 278054
rect 180352 269074 180380 287098
rect 180340 269068 180392 269074
rect 180340 269010 180392 269016
rect 180340 250504 180392 250510
rect 180340 250446 180392 250452
rect 180352 231810 180380 250446
rect 181456 234569 181484 324391
rect 181548 311234 181576 358838
rect 181626 335608 181682 335617
rect 181626 335543 181682 335552
rect 181640 324970 181668 335543
rect 181628 324964 181680 324970
rect 181628 324906 181680 324912
rect 181536 311228 181588 311234
rect 181536 311170 181588 311176
rect 181628 304292 181680 304298
rect 181628 304234 181680 304240
rect 181534 288688 181590 288697
rect 181534 288623 181590 288632
rect 181442 234560 181498 234569
rect 181442 234495 181498 234504
rect 180340 231804 180392 231810
rect 180340 231746 180392 231752
rect 181548 217938 181576 288623
rect 181640 281450 181668 304234
rect 181628 281444 181680 281450
rect 181628 281386 181680 281392
rect 181628 269612 181680 269618
rect 181628 269554 181680 269560
rect 181640 235958 181668 269554
rect 182180 259480 182232 259486
rect 182180 259422 182232 259428
rect 182192 256737 182220 259422
rect 182178 256728 182234 256737
rect 182178 256663 182234 256672
rect 181628 235952 181680 235958
rect 181628 235894 181680 235900
rect 181536 217932 181588 217938
rect 181536 217874 181588 217880
rect 180338 194032 180394 194041
rect 180338 193967 180394 193976
rect 180248 191752 180300 191758
rect 180248 191694 180300 191700
rect 180246 188456 180302 188465
rect 180246 188391 180302 188400
rect 180156 184204 180208 184210
rect 180156 184146 180208 184152
rect 180154 108352 180210 108361
rect 180154 108287 180210 108296
rect 180168 66230 180196 108287
rect 180156 66224 180208 66230
rect 180156 66166 180208 66172
rect 180062 46200 180118 46209
rect 180062 46135 180118 46144
rect 180062 43480 180118 43489
rect 180062 43415 180118 43424
rect 180076 10334 180104 43415
rect 180260 37913 180288 188391
rect 180352 187649 180380 193967
rect 181442 189952 181498 189961
rect 181442 189887 181498 189896
rect 180338 187640 180394 187649
rect 180338 187575 180394 187584
rect 180338 183696 180394 183705
rect 180338 183631 180394 183640
rect 180352 157282 180380 183631
rect 180340 157276 180392 157282
rect 180340 157218 180392 157224
rect 180246 37904 180302 37913
rect 180246 37839 180302 37848
rect 181456 15978 181484 189887
rect 181548 185638 181576 217874
rect 181536 185632 181588 185638
rect 181536 185574 181588 185580
rect 181640 179353 181668 235894
rect 181626 179344 181682 179353
rect 181626 179279 181682 179288
rect 181534 176896 181590 176905
rect 181534 176831 181590 176840
rect 181548 158642 181576 176831
rect 181536 158636 181588 158642
rect 181536 158578 181588 158584
rect 181536 131776 181588 131782
rect 181536 131718 181588 131724
rect 181548 73098 181576 131718
rect 181628 118720 181680 118726
rect 181628 118662 181680 118668
rect 181640 89690 181668 118662
rect 181628 89684 181680 89690
rect 181628 89626 181680 89632
rect 181536 73092 181588 73098
rect 181536 73034 181588 73040
rect 182836 35193 182864 368494
rect 184202 349344 184258 349353
rect 184202 349279 184258 349288
rect 182916 335436 182968 335442
rect 182916 335378 182968 335384
rect 182928 273970 182956 335378
rect 184216 318102 184244 349279
rect 184296 338156 184348 338162
rect 184296 338098 184348 338104
rect 184204 318096 184256 318102
rect 184204 318038 184256 318044
rect 184204 299600 184256 299606
rect 184204 299542 184256 299548
rect 184216 281518 184244 299542
rect 184204 281512 184256 281518
rect 184204 281454 184256 281460
rect 182916 273964 182968 273970
rect 182916 273906 182968 273912
rect 184204 266416 184256 266422
rect 184204 266358 184256 266364
rect 183466 257272 183522 257281
rect 183466 257207 183522 257216
rect 183480 256737 183508 257207
rect 183466 256728 183522 256737
rect 183466 256663 183522 256672
rect 182916 256216 182968 256222
rect 182916 256158 182968 256164
rect 182928 233238 182956 256158
rect 182916 233232 182968 233238
rect 182916 233174 182968 233180
rect 182916 184952 182968 184958
rect 182916 184894 182968 184900
rect 182928 160070 182956 184894
rect 183480 178673 183508 256663
rect 183466 178664 183522 178673
rect 183466 178599 183522 178608
rect 182916 160064 182968 160070
rect 182916 160006 182968 160012
rect 182914 109168 182970 109177
rect 182914 109103 182970 109112
rect 182928 84182 182956 109103
rect 182916 84176 182968 84182
rect 182916 84118 182968 84124
rect 182822 35184 182878 35193
rect 182822 35119 182878 35128
rect 181444 15972 181496 15978
rect 181444 15914 181496 15920
rect 184216 10334 184244 266358
rect 184308 259350 184336 338098
rect 184386 295352 184442 295361
rect 184386 295287 184442 295296
rect 184296 259344 184348 259350
rect 184296 259286 184348 259292
rect 184400 234530 184428 295287
rect 184848 282192 184900 282198
rect 184848 282134 184900 282140
rect 185032 282192 185084 282198
rect 185032 282134 185084 282140
rect 184860 281586 184888 282134
rect 184848 281580 184900 281586
rect 184848 281522 184900 281528
rect 184756 259344 184808 259350
rect 184756 259286 184808 259292
rect 184768 258738 184796 259286
rect 184756 258732 184808 258738
rect 184756 258674 184808 258680
rect 184388 234524 184440 234530
rect 184388 234466 184440 234472
rect 184768 188465 184796 258674
rect 184754 188456 184810 188465
rect 184754 188391 184810 188400
rect 184860 186998 184888 281522
rect 185044 278050 185072 282134
rect 185032 278044 185084 278050
rect 185032 277986 185084 277992
rect 185596 273154 185624 376722
rect 185766 336832 185822 336841
rect 185766 336767 185822 336776
rect 185674 323640 185730 323649
rect 185674 323575 185730 323584
rect 185584 273148 185636 273154
rect 185584 273090 185636 273096
rect 185688 250510 185716 323575
rect 185780 322318 185808 336767
rect 185768 322312 185820 322318
rect 185768 322254 185820 322260
rect 185766 284880 185822 284889
rect 185766 284815 185822 284824
rect 185676 250504 185728 250510
rect 185676 250446 185728 250452
rect 185584 236700 185636 236706
rect 185584 236642 185636 236648
rect 184848 186992 184900 186998
rect 184848 186934 184900 186940
rect 184296 150544 184348 150550
rect 184296 150486 184348 150492
rect 184308 110430 184336 150486
rect 185596 142866 185624 236642
rect 185780 230489 185808 284815
rect 186318 273456 186374 273465
rect 186318 273391 186374 273400
rect 186332 269618 186360 273391
rect 186320 269612 186372 269618
rect 186320 269554 186372 269560
rect 186136 264988 186188 264994
rect 186136 264930 186188 264936
rect 185860 247716 185912 247722
rect 185860 247658 185912 247664
rect 185872 247110 185900 247658
rect 185860 247104 185912 247110
rect 185860 247046 185912 247052
rect 185766 230480 185822 230489
rect 185766 230415 185822 230424
rect 186148 200190 186176 264930
rect 186976 261594 187004 438874
rect 188344 379568 188396 379574
rect 188344 379510 188396 379516
rect 187056 308440 187108 308446
rect 187056 308382 187108 308388
rect 186964 261588 187016 261594
rect 186964 261530 187016 261536
rect 186976 256018 187004 261530
rect 186964 256012 187016 256018
rect 186964 255954 187016 255960
rect 186964 249824 187016 249830
rect 186964 249766 187016 249772
rect 186228 247104 186280 247110
rect 186228 247046 186280 247052
rect 186136 200184 186188 200190
rect 186136 200126 186188 200132
rect 186148 197334 186176 200126
rect 186136 197328 186188 197334
rect 186136 197270 186188 197276
rect 186240 180198 186268 247046
rect 186976 237250 187004 249766
rect 187068 247353 187096 308382
rect 188356 264926 188384 379510
rect 188436 362976 188488 362982
rect 188436 362918 188488 362924
rect 188448 286385 188476 362918
rect 188526 351928 188582 351937
rect 188526 351863 188582 351872
rect 188540 329186 188568 351863
rect 191116 349081 191144 445839
rect 582392 432614 582420 484599
rect 582654 471472 582710 471481
rect 582654 471407 582710 471416
rect 582470 458144 582526 458153
rect 582470 458079 582526 458088
rect 582484 449206 582512 458079
rect 582472 449200 582524 449206
rect 582472 449142 582524 449148
rect 582380 432608 582432 432614
rect 582380 432550 582432 432556
rect 582378 431624 582434 431633
rect 582378 431559 582434 431568
rect 582392 403646 582420 431559
rect 582470 418296 582526 418305
rect 582470 418231 582526 418240
rect 582380 403640 582432 403646
rect 582380 403582 582432 403588
rect 211804 374060 211856 374066
rect 211804 374002 211856 374008
rect 204904 372632 204956 372638
rect 204904 372574 204956 372580
rect 202142 359000 202198 359009
rect 202142 358935 202198 358944
rect 193862 357504 193918 357513
rect 193862 357439 193918 357448
rect 191102 349072 191158 349081
rect 191102 349007 191158 349016
rect 191746 349072 191802 349081
rect 191746 349007 191802 349016
rect 188528 329180 188580 329186
rect 188528 329122 188580 329128
rect 189722 320784 189778 320793
rect 189722 320719 189778 320728
rect 188434 286376 188490 286385
rect 188434 286311 188490 286320
rect 188988 283620 189040 283626
rect 188988 283562 189040 283568
rect 188434 279440 188490 279449
rect 188434 279375 188490 279384
rect 188344 264920 188396 264926
rect 188344 264862 188396 264868
rect 187240 264240 187292 264246
rect 187240 264182 187292 264188
rect 187054 247344 187110 247353
rect 187054 247279 187110 247288
rect 187148 247104 187200 247110
rect 187148 247046 187200 247052
rect 186964 237244 187016 237250
rect 186964 237186 187016 237192
rect 186964 202224 187016 202230
rect 186964 202166 187016 202172
rect 186228 180192 186280 180198
rect 186228 180134 186280 180140
rect 185674 179480 185730 179489
rect 185674 179415 185730 179424
rect 185688 162790 185716 179415
rect 185676 162784 185728 162790
rect 185676 162726 185728 162732
rect 185676 146328 185728 146334
rect 185676 146270 185728 146276
rect 185584 142860 185636 142866
rect 185584 142802 185636 142808
rect 184388 112464 184440 112470
rect 184388 112406 184440 112412
rect 184296 110424 184348 110430
rect 184296 110366 184348 110372
rect 184296 86284 184348 86290
rect 184296 86226 184348 86232
rect 184308 38010 184336 86226
rect 184400 82754 184428 112406
rect 184480 106412 184532 106418
rect 184480 106354 184532 106360
rect 184492 86737 184520 106354
rect 184664 97300 184716 97306
rect 184664 97242 184716 97248
rect 184478 86728 184534 86737
rect 184478 86663 184534 86672
rect 184676 86601 184704 97242
rect 185688 96014 185716 146270
rect 186976 141506 187004 202166
rect 187160 200114 187188 247046
rect 187252 230450 187280 264182
rect 187700 254584 187752 254590
rect 187700 254526 187752 254532
rect 187712 253978 187740 254526
rect 187700 253972 187752 253978
rect 187700 253914 187752 253920
rect 187608 252680 187660 252686
rect 187608 252622 187660 252628
rect 187240 230444 187292 230450
rect 187240 230386 187292 230392
rect 187068 200086 187188 200114
rect 187068 200054 187096 200086
rect 187056 200048 187108 200054
rect 187056 199990 187108 199996
rect 187068 188426 187096 199990
rect 187620 198694 187648 252622
rect 187700 251864 187752 251870
rect 187700 251806 187752 251812
rect 187712 251258 187740 251806
rect 187700 251252 187752 251258
rect 187700 251194 187752 251200
rect 187700 230512 187752 230518
rect 187698 230480 187700 230489
rect 187752 230480 187754 230489
rect 187698 230415 187754 230424
rect 188068 223576 188120 223582
rect 188068 223518 188120 223524
rect 188080 222902 188108 223518
rect 188068 222896 188120 222902
rect 188068 222838 188120 222844
rect 187700 222148 187752 222154
rect 187700 222090 187752 222096
rect 187712 222057 187740 222090
rect 187698 222048 187754 222057
rect 188448 222018 188476 279375
rect 189000 278905 189028 283562
rect 188986 278896 189042 278905
rect 188986 278831 189042 278840
rect 188804 254584 188856 254590
rect 188804 254526 188856 254532
rect 188816 234530 188844 254526
rect 188896 251252 188948 251258
rect 188896 251194 188948 251200
rect 188804 234524 188856 234530
rect 188804 234466 188856 234472
rect 188804 223576 188856 223582
rect 188804 223518 188856 223524
rect 187698 221983 187754 221992
rect 188436 222012 188488 222018
rect 188436 221954 188488 221960
rect 187608 198688 187660 198694
rect 187608 198630 187660 198636
rect 187056 188420 187108 188426
rect 187056 188362 187108 188368
rect 187056 178152 187108 178158
rect 187056 178094 187108 178100
rect 187068 169658 187096 178094
rect 188816 176594 188844 223518
rect 188908 193934 188936 251194
rect 188896 193928 188948 193934
rect 188896 193870 188948 193876
rect 189000 189786 189028 278831
rect 189080 217388 189132 217394
rect 189080 217330 189132 217336
rect 189092 211138 189120 217330
rect 189080 211132 189132 211138
rect 189080 211074 189132 211080
rect 189264 195900 189316 195906
rect 189264 195842 189316 195848
rect 189276 195362 189304 195842
rect 189264 195356 189316 195362
rect 189264 195298 189316 195304
rect 188988 189780 189040 189786
rect 188988 189722 189040 189728
rect 188804 176588 188856 176594
rect 188804 176530 188856 176536
rect 187056 169652 187108 169658
rect 187056 169594 187108 169600
rect 188344 159384 188396 159390
rect 188344 159326 188396 159332
rect 186964 141500 187016 141506
rect 186964 141442 187016 141448
rect 185768 127084 185820 127090
rect 185768 127026 185820 127032
rect 185676 96008 185728 96014
rect 185676 95950 185728 95956
rect 185582 89040 185638 89049
rect 185582 88975 185638 88984
rect 184662 86592 184718 86601
rect 184662 86527 184718 86536
rect 184388 82748 184440 82754
rect 184388 82690 184440 82696
rect 184296 38004 184348 38010
rect 184296 37946 184348 37952
rect 185596 35290 185624 88975
rect 185780 80073 185808 127026
rect 186964 124908 187016 124914
rect 186964 124850 187016 124856
rect 185766 80064 185822 80073
rect 185766 79999 185822 80008
rect 186976 62082 187004 124850
rect 187056 111852 187108 111858
rect 187056 111794 187108 111800
rect 187068 82822 187096 111794
rect 187976 95260 188028 95266
rect 187976 95202 188028 95208
rect 187988 88233 188016 95202
rect 187974 88224 188030 88233
rect 187974 88159 188030 88168
rect 187056 82816 187108 82822
rect 187056 82758 187108 82764
rect 186964 62076 187016 62082
rect 186964 62018 187016 62024
rect 185584 35284 185636 35290
rect 185584 35226 185636 35232
rect 188356 21486 188384 159326
rect 188436 113280 188488 113286
rect 188436 113222 188488 113228
rect 188448 89729 188476 113222
rect 188434 89720 188490 89729
rect 188434 89655 188490 89664
rect 189736 42129 189764 320719
rect 189816 316736 189868 316742
rect 189816 316678 189868 316684
rect 189828 256698 189856 316678
rect 191102 311128 191158 311137
rect 191102 311063 191158 311072
rect 191116 305318 191144 311063
rect 191104 305312 191156 305318
rect 191104 305254 191156 305260
rect 191656 305312 191708 305318
rect 191656 305254 191708 305260
rect 191668 305046 191696 305254
rect 191656 305040 191708 305046
rect 191656 304982 191708 304988
rect 191104 296744 191156 296750
rect 191104 296686 191156 296692
rect 190366 286104 190422 286113
rect 190366 286039 190422 286048
rect 189816 256692 189868 256698
rect 189816 256634 189868 256640
rect 189906 255912 189962 255921
rect 189906 255847 189962 255856
rect 189816 246356 189868 246362
rect 189816 246298 189868 246304
rect 189828 231577 189856 246298
rect 189920 235958 189948 255847
rect 189908 235952 189960 235958
rect 189908 235894 189960 235900
rect 189814 231568 189870 231577
rect 189814 231503 189870 231512
rect 190380 195362 190408 286039
rect 191116 274650 191144 296686
rect 191194 292632 191250 292641
rect 191194 292567 191250 292576
rect 191208 286346 191236 292567
rect 191196 286340 191248 286346
rect 191196 286282 191248 286288
rect 191196 283960 191248 283966
rect 191196 283902 191248 283908
rect 191104 274644 191156 274650
rect 191104 274586 191156 274592
rect 191104 255332 191156 255338
rect 191104 255274 191156 255280
rect 191116 223582 191144 255274
rect 191208 253201 191236 283902
rect 191668 278730 191696 304982
rect 191760 292641 191788 349007
rect 192484 335368 192536 335374
rect 192484 335310 192536 335316
rect 191746 292632 191802 292641
rect 191746 292567 191802 292576
rect 191656 278724 191708 278730
rect 191656 278666 191708 278672
rect 191380 271176 191432 271182
rect 191380 271118 191432 271124
rect 191194 253192 191250 253201
rect 191194 253127 191250 253136
rect 191196 249824 191248 249830
rect 191196 249766 191248 249772
rect 191104 223576 191156 223582
rect 191104 223518 191156 223524
rect 191102 221640 191158 221649
rect 191102 221575 191158 221584
rect 190368 195356 190420 195362
rect 190368 195298 190420 195304
rect 189816 116000 189868 116006
rect 189816 115942 189868 115948
rect 189828 88097 189856 115942
rect 189814 88088 189870 88097
rect 189814 88023 189870 88032
rect 189722 42120 189778 42129
rect 189722 42055 189778 42064
rect 188344 21480 188396 21486
rect 188344 21422 188396 21428
rect 180064 10328 180116 10334
rect 180064 10270 180116 10276
rect 184204 10328 184256 10334
rect 184204 10270 184256 10276
rect 177304 9036 177356 9042
rect 177304 8978 177356 8984
rect 191116 3505 191144 221575
rect 191208 219434 191236 249766
rect 191392 249694 191420 271118
rect 191380 249688 191432 249694
rect 191380 249630 191432 249636
rect 191288 249076 191340 249082
rect 191288 249018 191340 249024
rect 191300 226001 191328 249018
rect 191748 245676 191800 245682
rect 191748 245618 191800 245624
rect 191654 242584 191710 242593
rect 191654 242519 191710 242528
rect 191668 241641 191696 242519
rect 191654 241632 191710 241641
rect 191654 241567 191710 241576
rect 191668 241534 191696 241567
rect 191656 241528 191708 241534
rect 191656 241470 191708 241476
rect 191760 226953 191788 245618
rect 192496 244186 192524 335310
rect 192852 327752 192904 327758
rect 192852 327694 192904 327700
rect 192864 326369 192892 327694
rect 192850 326360 192906 326369
rect 192850 326295 192906 326304
rect 193876 320958 193904 357439
rect 200762 356144 200818 356153
rect 200762 356079 200818 356088
rect 198002 353560 198058 353569
rect 198002 353495 198058 353504
rect 195244 352028 195296 352034
rect 195244 351970 195296 351976
rect 193954 327040 194010 327049
rect 193954 326975 194010 326984
rect 193864 320952 193916 320958
rect 193864 320894 193916 320900
rect 193864 311908 193916 311914
rect 193864 311850 193916 311856
rect 192668 305652 192720 305658
rect 192668 305594 192720 305600
rect 192576 278860 192628 278866
rect 192576 278802 192628 278808
rect 192588 257378 192616 278802
rect 192576 257372 192628 257378
rect 192576 257314 192628 257320
rect 192484 244180 192536 244186
rect 192484 244122 192536 244128
rect 192484 234524 192536 234530
rect 192484 234466 192536 234472
rect 191746 226944 191802 226953
rect 191746 226879 191802 226888
rect 191286 225992 191342 226001
rect 191286 225927 191342 225936
rect 192496 220289 192524 234466
rect 192482 220280 192538 220289
rect 192482 220215 192538 220224
rect 191208 219406 191328 219434
rect 191300 216646 191328 219406
rect 191288 216640 191340 216646
rect 191288 216582 191340 216588
rect 191194 214704 191250 214713
rect 191194 214639 191250 214648
rect 191208 118289 191236 214639
rect 191300 191214 191328 216582
rect 192588 198694 192616 257314
rect 192680 249762 192708 305594
rect 193876 294642 193904 311850
rect 193864 294636 193916 294642
rect 193864 294578 193916 294584
rect 193864 291236 193916 291242
rect 193864 291178 193916 291184
rect 193036 253972 193088 253978
rect 193036 253914 193088 253920
rect 192668 249756 192720 249762
rect 192668 249698 192720 249704
rect 192668 242956 192720 242962
rect 192668 242898 192720 242904
rect 192680 234530 192708 242898
rect 192668 234524 192720 234530
rect 192668 234466 192720 234472
rect 193048 223650 193076 253914
rect 193128 249688 193180 249694
rect 193128 249630 193180 249636
rect 193036 223644 193088 223650
rect 193036 223586 193088 223592
rect 193048 222154 193076 223586
rect 193036 222148 193088 222154
rect 193036 222090 193088 222096
rect 193036 220720 193088 220726
rect 193036 220662 193088 220668
rect 193048 220114 193076 220662
rect 193036 220108 193088 220114
rect 193036 220050 193088 220056
rect 192576 198688 192628 198694
rect 192576 198630 192628 198636
rect 191288 191208 191340 191214
rect 191288 191150 191340 191156
rect 193048 184385 193076 220050
rect 193140 202230 193168 249630
rect 193404 244384 193456 244390
rect 193404 244326 193456 244332
rect 193416 243642 193444 244326
rect 193404 243636 193456 243642
rect 193404 243578 193456 243584
rect 193876 241466 193904 291178
rect 193968 291145 193996 326975
rect 193954 291136 194010 291145
rect 193954 291071 194010 291080
rect 194506 291136 194562 291145
rect 194506 291071 194562 291080
rect 194520 290057 194548 291071
rect 194506 290048 194562 290057
rect 194506 289983 194562 289992
rect 193956 259480 194008 259486
rect 193956 259422 194008 259428
rect 193864 241460 193916 241466
rect 193864 241402 193916 241408
rect 193968 220726 193996 259422
rect 194048 243568 194100 243574
rect 194048 243510 194100 243516
rect 194060 233170 194088 243510
rect 194048 233164 194100 233170
rect 194048 233106 194100 233112
rect 193956 220720 194008 220726
rect 193956 220662 194008 220668
rect 193956 215960 194008 215966
rect 193956 215902 194008 215908
rect 193864 209160 193916 209166
rect 193864 209102 193916 209108
rect 193128 202224 193180 202230
rect 193128 202166 193180 202172
rect 193034 184376 193090 184385
rect 193034 184311 193090 184320
rect 192484 184204 192536 184210
rect 192484 184146 192536 184152
rect 191286 180840 191342 180849
rect 191286 180775 191342 180784
rect 191300 165510 191328 180775
rect 191288 165504 191340 165510
rect 191288 165446 191340 165452
rect 191288 131164 191340 131170
rect 191288 131106 191340 131112
rect 191194 118280 191250 118289
rect 191194 118215 191250 118224
rect 191196 103556 191248 103562
rect 191196 103498 191248 103504
rect 191208 73137 191236 103498
rect 191194 73128 191250 73137
rect 191194 73063 191250 73072
rect 191300 59362 191328 131106
rect 191380 120148 191432 120154
rect 191380 120090 191432 120096
rect 191392 102814 191420 120090
rect 191380 102808 191432 102814
rect 191380 102750 191432 102756
rect 191288 59356 191340 59362
rect 191288 59298 191340 59304
rect 192496 28257 192524 184146
rect 192576 141432 192628 141438
rect 192576 141374 192628 141380
rect 192588 92313 192616 141374
rect 192668 102264 192720 102270
rect 192668 102206 192720 102212
rect 192574 92304 192630 92313
rect 192574 92239 192630 92248
rect 192680 64802 192708 102206
rect 192668 64796 192720 64802
rect 192668 64738 192720 64744
rect 192482 28248 192538 28257
rect 192482 28183 192538 28192
rect 193876 10305 193904 209102
rect 193968 190466 193996 215902
rect 194520 209137 194548 289983
rect 195256 267170 195284 351970
rect 196624 347880 196676 347886
rect 196624 347822 196676 347828
rect 195334 334248 195390 334257
rect 195334 334183 195390 334192
rect 195348 285705 195376 334183
rect 195428 331356 195480 331362
rect 195428 331298 195480 331304
rect 195440 313954 195468 331298
rect 195428 313948 195480 313954
rect 195428 313890 195480 313896
rect 195978 305688 196034 305697
rect 195978 305623 196034 305632
rect 195992 305017 196020 305623
rect 195978 305008 196034 305017
rect 195978 304943 196034 304952
rect 195334 285696 195390 285705
rect 195334 285631 195390 285640
rect 195428 279744 195480 279750
rect 195428 279686 195480 279692
rect 195244 267164 195296 267170
rect 195244 267106 195296 267112
rect 195244 263628 195296 263634
rect 195244 263570 195296 263576
rect 195256 262274 195284 263570
rect 195244 262268 195296 262274
rect 195244 262210 195296 262216
rect 194692 234728 194744 234734
rect 194692 234670 194744 234676
rect 194704 232937 194732 234670
rect 195150 233880 195206 233889
rect 195150 233815 195206 233824
rect 195164 232937 195192 233815
rect 194690 232928 194746 232937
rect 194690 232863 194746 232872
rect 195150 232928 195206 232937
rect 195150 232863 195206 232872
rect 194968 227044 195020 227050
rect 194968 226986 195020 226992
rect 194980 223582 195008 226986
rect 194968 223576 195020 223582
rect 194968 223518 195020 223524
rect 194506 209128 194562 209137
rect 194506 209063 194562 209072
rect 195256 196722 195284 262210
rect 195440 255338 195468 279686
rect 195520 273964 195572 273970
rect 195520 273906 195572 273912
rect 195428 255332 195480 255338
rect 195428 255274 195480 255280
rect 195336 241528 195388 241534
rect 195336 241470 195388 241476
rect 195348 213926 195376 241470
rect 195532 234433 195560 273906
rect 196636 265849 196664 347822
rect 196716 326392 196768 326398
rect 196716 326334 196768 326340
rect 196728 274582 196756 326334
rect 197266 305008 197322 305017
rect 197266 304943 197322 304952
rect 197280 292641 197308 304943
rect 197360 294704 197412 294710
rect 197360 294646 197412 294652
rect 197266 292632 197322 292641
rect 197266 292567 197322 292576
rect 197372 291854 197400 294646
rect 197360 291848 197412 291854
rect 197360 291790 197412 291796
rect 197082 288824 197138 288833
rect 197082 288759 197138 288768
rect 197096 282198 197124 288759
rect 197358 282432 197414 282441
rect 197358 282367 197414 282376
rect 197084 282192 197136 282198
rect 197084 282134 197136 282140
rect 197372 281586 197400 282367
rect 198016 281625 198044 353495
rect 198096 332648 198148 332654
rect 198096 332590 198148 332596
rect 198002 281616 198058 281625
rect 197360 281580 197412 281586
rect 198002 281551 198058 281560
rect 197360 281522 197412 281528
rect 197360 281444 197412 281450
rect 197360 281386 197412 281392
rect 197372 280809 197400 281386
rect 197358 280800 197414 280809
rect 197358 280735 197414 280744
rect 197358 280256 197414 280265
rect 197358 280191 197414 280200
rect 196898 279304 196954 279313
rect 196898 279239 196954 279248
rect 196716 274576 196768 274582
rect 196716 274518 196768 274524
rect 196622 265840 196678 265849
rect 196622 265775 196678 265784
rect 196622 262304 196678 262313
rect 196622 262239 196678 262248
rect 195888 249756 195940 249762
rect 195888 249698 195940 249704
rect 195900 248742 195928 249698
rect 195888 248736 195940 248742
rect 195888 248678 195940 248684
rect 195900 236502 195928 248678
rect 196636 246265 196664 262239
rect 196622 246256 196678 246265
rect 196622 246191 196678 246200
rect 196912 237318 196940 279239
rect 197372 278866 197400 280191
rect 197360 278860 197412 278866
rect 197360 278802 197412 278808
rect 198108 278769 198136 332590
rect 199384 326460 199436 326466
rect 199384 326402 199436 326408
rect 199396 302190 199424 326402
rect 199384 302184 199436 302190
rect 199384 302126 199436 302132
rect 200580 302184 200632 302190
rect 200580 302126 200632 302132
rect 200592 300898 200620 302126
rect 200120 300892 200172 300898
rect 200120 300834 200172 300840
rect 200580 300892 200632 300898
rect 200580 300834 200632 300840
rect 200028 294024 200080 294030
rect 200028 293966 200080 293972
rect 199476 289944 199528 289950
rect 199476 289886 199528 289892
rect 198186 287464 198242 287473
rect 198186 287399 198242 287408
rect 198094 278760 198150 278769
rect 197360 278724 197412 278730
rect 198094 278695 198150 278704
rect 197360 278666 197412 278672
rect 197372 278089 197400 278666
rect 197358 278080 197414 278089
rect 197358 278015 197414 278024
rect 197360 276752 197412 276758
rect 197358 276720 197360 276729
rect 197412 276720 197414 276729
rect 197280 276678 197358 276706
rect 197084 250504 197136 250510
rect 197084 250446 197136 250452
rect 197096 245177 197124 250446
rect 197082 245168 197138 245177
rect 197082 245103 197138 245112
rect 196900 237312 196952 237318
rect 196900 237254 196952 237260
rect 195888 236496 195940 236502
rect 195888 236438 195940 236444
rect 196808 236496 196860 236502
rect 196808 236438 196860 236444
rect 195518 234424 195574 234433
rect 195518 234359 195574 234368
rect 195426 223000 195482 223009
rect 195426 222935 195482 222944
rect 195440 216617 195468 222935
rect 196622 221504 196678 221513
rect 196622 221439 196678 221448
rect 195426 216608 195482 216617
rect 195426 216543 195482 216552
rect 195336 213920 195388 213926
rect 195336 213862 195388 213868
rect 195244 196716 195296 196722
rect 195244 196658 195296 196664
rect 193956 190460 194008 190466
rect 193956 190402 194008 190408
rect 193956 186380 194008 186386
rect 193956 186322 194008 186328
rect 193968 161362 193996 186322
rect 195348 177449 195376 213862
rect 195428 203584 195480 203590
rect 195428 203526 195480 203532
rect 195440 189961 195468 203526
rect 195426 189952 195482 189961
rect 195426 189887 195482 189896
rect 195334 177440 195390 177449
rect 195334 177375 195390 177384
rect 195518 177168 195574 177177
rect 195518 177103 195574 177112
rect 193956 161356 194008 161362
rect 193956 161298 194008 161304
rect 195532 160002 195560 177103
rect 195520 159996 195572 160002
rect 195520 159938 195572 159944
rect 195244 141500 195296 141506
rect 195244 141442 195296 141448
rect 193954 118824 194010 118833
rect 193954 118759 194010 118768
rect 193968 89457 193996 118759
rect 195256 91769 195284 141442
rect 195336 115252 195388 115258
rect 195336 115194 195388 115200
rect 195242 91760 195298 91769
rect 195242 91695 195298 91704
rect 193954 89448 194010 89457
rect 193954 89383 194010 89392
rect 195244 83564 195296 83570
rect 195244 83506 195296 83512
rect 193862 10296 193918 10305
rect 193862 10231 193918 10240
rect 191102 3496 191158 3505
rect 191102 3431 191158 3440
rect 195256 2009 195284 83506
rect 195348 66162 195376 115194
rect 195336 66156 195388 66162
rect 195336 66098 195388 66104
rect 196636 3505 196664 221439
rect 196714 189816 196770 189825
rect 196714 189751 196770 189760
rect 196728 87553 196756 189751
rect 196820 183161 196848 236438
rect 197096 221474 197124 245103
rect 197176 244180 197228 244186
rect 197176 244122 197228 244128
rect 197084 221468 197136 221474
rect 197084 221410 197136 221416
rect 197188 216073 197216 244122
rect 197174 216064 197230 216073
rect 197174 215999 197230 216008
rect 196900 196648 196952 196654
rect 196900 196590 196952 196596
rect 196806 183152 196862 183161
rect 196806 183087 196862 183096
rect 196912 181529 196940 196590
rect 197280 192574 197308 276678
rect 197358 276655 197414 276664
rect 197358 275088 197414 275097
rect 197358 275023 197414 275032
rect 197372 274786 197400 275023
rect 197360 274780 197412 274786
rect 197360 274722 197412 274728
rect 197360 273216 197412 273222
rect 197360 273158 197412 273164
rect 197372 272921 197400 273158
rect 197452 273148 197504 273154
rect 197452 273090 197504 273096
rect 197358 272912 197414 272921
rect 197358 272847 197414 272856
rect 197464 272377 197492 273090
rect 197450 272368 197506 272377
rect 197450 272303 197506 272312
rect 197450 271552 197506 271561
rect 197450 271487 197506 271496
rect 197464 270570 197492 271487
rect 197452 270564 197504 270570
rect 197452 270506 197504 270512
rect 197360 270496 197412 270502
rect 197360 270438 197412 270444
rect 197372 269385 197400 270438
rect 197358 269376 197414 269385
rect 197358 269311 197414 269320
rect 197360 269000 197412 269006
rect 197360 268942 197412 268948
rect 197372 268841 197400 268942
rect 197358 268832 197414 268841
rect 197358 268767 197414 268776
rect 197360 268388 197412 268394
rect 197360 268330 197412 268336
rect 197372 268025 197400 268330
rect 197358 268016 197414 268025
rect 197358 267951 197414 267960
rect 197358 267200 197414 267209
rect 197358 267135 197414 267144
rect 197452 267164 197504 267170
rect 197372 266490 197400 267135
rect 197452 267106 197504 267112
rect 197464 266665 197492 267106
rect 198200 267073 198228 287399
rect 198832 285796 198884 285802
rect 198832 285738 198884 285744
rect 198738 284336 198794 284345
rect 198738 284271 198794 284280
rect 198752 279750 198780 284271
rect 198740 279744 198792 279750
rect 198740 279686 198792 279692
rect 198646 278760 198702 278769
rect 198646 278695 198702 278704
rect 198554 271008 198610 271017
rect 198554 270943 198610 270952
rect 198186 267064 198242 267073
rect 198186 266999 198242 267008
rect 197450 266656 197506 266665
rect 197450 266591 197506 266600
rect 197360 266484 197412 266490
rect 197360 266426 197412 266432
rect 197358 265296 197414 265305
rect 197358 265231 197414 265240
rect 197372 264994 197400 265231
rect 197360 264988 197412 264994
rect 197360 264930 197412 264936
rect 197452 264920 197504 264926
rect 197452 264862 197504 264868
rect 197464 264489 197492 264862
rect 197450 264480 197506 264489
rect 197450 264415 197506 264424
rect 197358 263664 197414 263673
rect 197358 263599 197360 263608
rect 197412 263599 197414 263608
rect 197360 263570 197412 263576
rect 197360 261588 197412 261594
rect 197360 261530 197412 261536
rect 197372 261497 197400 261530
rect 197358 261488 197414 261497
rect 197358 261423 197414 261432
rect 198002 260944 198058 260953
rect 198002 260879 198058 260888
rect 197358 260128 197414 260137
rect 197358 260063 197414 260072
rect 197372 259486 197400 260063
rect 197360 259480 197412 259486
rect 197360 259422 197412 259428
rect 197452 259412 197504 259418
rect 197452 259354 197504 259360
rect 197358 259312 197414 259321
rect 197358 259247 197414 259256
rect 197372 258738 197400 259247
rect 197464 258777 197492 259354
rect 197450 258768 197506 258777
rect 197360 258732 197412 258738
rect 197450 258703 197506 258712
rect 197360 258674 197412 258680
rect 197450 257952 197506 257961
rect 197450 257887 197506 257896
rect 197464 256766 197492 257887
rect 197452 256760 197504 256766
rect 197452 256702 197504 256708
rect 197360 256692 197412 256698
rect 197360 256634 197412 256640
rect 197372 255785 197400 256634
rect 197358 255776 197414 255785
rect 197358 255711 197414 255720
rect 197358 255232 197414 255241
rect 197358 255167 197414 255176
rect 197372 253978 197400 255167
rect 198016 254590 198044 260879
rect 198568 259457 198596 270943
rect 198554 259448 198610 259457
rect 198554 259383 198610 259392
rect 198004 254584 198056 254590
rect 198004 254526 198056 254532
rect 197360 253972 197412 253978
rect 197360 253914 197412 253920
rect 197450 253600 197506 253609
rect 197450 253535 197506 253544
rect 197358 253056 197414 253065
rect 197358 252991 197414 253000
rect 197372 252686 197400 252991
rect 197360 252680 197412 252686
rect 197360 252622 197412 252628
rect 197464 252618 197492 253535
rect 197452 252612 197504 252618
rect 197452 252554 197504 252560
rect 198002 252240 198058 252249
rect 198002 252175 198058 252184
rect 197358 251696 197414 251705
rect 197358 251631 197414 251640
rect 197372 251258 197400 251631
rect 197360 251252 197412 251258
rect 197360 251194 197412 251200
rect 197358 250880 197414 250889
rect 197358 250815 197414 250824
rect 197372 249830 197400 250815
rect 197360 249824 197412 249830
rect 197360 249766 197412 249772
rect 197360 249688 197412 249694
rect 197360 249630 197412 249636
rect 197372 249529 197400 249630
rect 197358 249520 197414 249529
rect 197358 249455 197414 249464
rect 197360 248736 197412 248742
rect 197358 248704 197360 248713
rect 197412 248704 197414 248713
rect 197358 248639 197414 248648
rect 197358 247888 197414 247897
rect 197358 247823 197414 247832
rect 197372 247110 197400 247823
rect 197360 247104 197412 247110
rect 197360 247046 197412 247052
rect 197358 246528 197414 246537
rect 197358 246463 197414 246472
rect 197372 245682 197400 246463
rect 197360 245676 197412 245682
rect 197360 245618 197412 245624
rect 197450 244352 197506 244361
rect 197450 244287 197506 244296
rect 197464 244186 197492 244287
rect 197452 244180 197504 244186
rect 197452 244122 197504 244128
rect 197360 243636 197412 243642
rect 197360 243578 197412 243584
rect 197372 243001 197400 243578
rect 197358 242992 197414 243001
rect 197358 242927 197414 242936
rect 198016 242593 198044 252175
rect 198002 242584 198058 242593
rect 198002 242519 198058 242528
rect 197360 242208 197412 242214
rect 197360 242150 197412 242156
rect 197542 242176 197598 242185
rect 197372 241641 197400 242150
rect 197542 242111 197598 242120
rect 197358 241632 197414 241641
rect 197358 241567 197414 241576
rect 197556 241534 197584 242111
rect 197544 241528 197596 241534
rect 197544 241470 197596 241476
rect 197360 241460 197412 241466
rect 197360 241402 197412 241408
rect 197372 240825 197400 241402
rect 197358 240816 197414 240825
rect 197358 240751 197414 240760
rect 198660 240174 198688 278695
rect 198844 278118 198872 285738
rect 199384 285728 199436 285734
rect 199384 285670 199436 285676
rect 198832 278112 198884 278118
rect 198832 278054 198884 278060
rect 199396 276690 199424 285670
rect 199488 282849 199516 289886
rect 200040 284617 200068 293966
rect 200132 285326 200160 300834
rect 200212 298172 200264 298178
rect 200212 298114 200264 298120
rect 200120 285320 200172 285326
rect 200120 285262 200172 285268
rect 200026 284608 200082 284617
rect 200026 284543 200082 284552
rect 200224 283914 200252 298114
rect 200776 291145 200804 356079
rect 202156 310418 202184 358935
rect 203524 354748 203576 354754
rect 203524 354690 203576 354696
rect 203064 347064 203116 347070
rect 203064 347006 203116 347012
rect 203076 346633 203104 347006
rect 203062 346624 203118 346633
rect 203062 346559 203118 346568
rect 203536 326398 203564 354690
rect 204352 347812 204404 347818
rect 204352 347754 204404 347760
rect 204168 347744 204220 347750
rect 204168 347686 204220 347692
rect 204180 347070 204208 347686
rect 204168 347064 204220 347070
rect 204168 347006 204220 347012
rect 203524 326392 203576 326398
rect 203524 326334 203576 326340
rect 202880 322312 202932 322318
rect 202880 322254 202932 322260
rect 202788 318164 202840 318170
rect 202788 318106 202840 318112
rect 201684 310412 201736 310418
rect 201684 310354 201736 310360
rect 202144 310412 202196 310418
rect 202144 310354 202196 310360
rect 201696 309194 201724 310354
rect 201684 309188 201736 309194
rect 201684 309130 201736 309136
rect 200762 291136 200818 291145
rect 200762 291071 200818 291080
rect 200776 287054 200804 291071
rect 200684 287026 200804 287054
rect 200684 284186 200712 287026
rect 200762 285696 200818 285705
rect 200762 285631 200818 285640
rect 201406 285696 201462 285705
rect 201406 285631 201462 285640
rect 200776 284617 200804 285631
rect 200948 285320 201000 285326
rect 200948 285262 201000 285268
rect 200762 284608 200818 284617
rect 200762 284543 200818 284552
rect 200422 284158 200712 284186
rect 200776 284172 200804 284543
rect 200960 284186 200988 285262
rect 200960 284158 201342 284186
rect 201420 283966 201448 285631
rect 201696 284172 201724 309130
rect 202234 288552 202290 288561
rect 202234 288487 202290 288496
rect 201958 284064 202014 284073
rect 202248 284050 202276 288487
rect 202800 284172 202828 318106
rect 202892 298178 202920 322254
rect 204364 306374 204392 347754
rect 204364 306346 204760 306374
rect 202880 298172 202932 298178
rect 202880 298114 202932 298120
rect 202892 297430 202920 298114
rect 202880 297424 202932 297430
rect 202880 297366 202932 297372
rect 203154 290048 203210 290057
rect 203154 289983 203210 289992
rect 203168 284172 203196 289983
rect 203706 285832 203762 285841
rect 203706 285767 203762 285776
rect 203720 284172 203748 285767
rect 204628 285728 204680 285734
rect 204628 285670 204680 285676
rect 204258 284472 204314 284481
rect 204258 284407 204314 284416
rect 204272 284172 204300 284407
rect 204640 284172 204668 285670
rect 202014 284036 202276 284050
rect 202014 284022 202262 284036
rect 201958 283999 202014 284008
rect 200132 283886 200252 283914
rect 201408 283960 201460 283966
rect 201408 283902 201460 283908
rect 204732 283914 204760 306346
rect 204916 285734 204944 372574
rect 206282 349480 206338 349489
rect 206282 349415 206338 349424
rect 204996 303680 205048 303686
rect 204996 303622 205048 303628
rect 205008 293282 205036 303622
rect 206296 298217 206324 349415
rect 210424 345092 210476 345098
rect 210424 345034 210476 345040
rect 209136 343664 209188 343670
rect 209136 343606 209188 343612
rect 209042 339688 209098 339697
rect 209042 339623 209098 339632
rect 206376 336796 206428 336802
rect 206376 336738 206428 336744
rect 206388 303686 206416 336738
rect 207662 331256 207718 331265
rect 207662 331191 207718 331200
rect 207676 316034 207704 331191
rect 207584 316006 207704 316034
rect 207584 311914 207612 316006
rect 207572 311908 207624 311914
rect 207572 311850 207624 311856
rect 206376 303680 206428 303686
rect 206376 303622 206428 303628
rect 207020 303680 207072 303686
rect 207020 303622 207072 303628
rect 206282 298208 206338 298217
rect 206282 298143 206338 298152
rect 206296 296714 206324 298143
rect 206296 296686 206692 296714
rect 204996 293276 205048 293282
rect 204996 293218 205048 293224
rect 204996 291236 205048 291242
rect 204996 291178 205048 291184
rect 204904 285728 204956 285734
rect 204904 285670 204956 285676
rect 205008 284889 205036 291178
rect 205548 285796 205600 285802
rect 205548 285738 205600 285744
rect 204994 284880 205050 284889
rect 204994 284815 205050 284824
rect 205560 284172 205588 285738
rect 206098 285696 206154 285705
rect 206098 285631 206154 285640
rect 206112 284172 206140 285631
rect 206664 284172 206692 296686
rect 207032 284172 207060 303622
rect 207584 284172 207612 311850
rect 208490 310584 208546 310593
rect 208490 310519 208546 310528
rect 208124 285728 208176 285734
rect 208124 285670 208176 285676
rect 208136 284172 208164 285670
rect 208504 284172 208532 310519
rect 209056 298178 209084 339623
rect 209148 310593 209176 343606
rect 209134 310584 209190 310593
rect 209134 310519 209190 310528
rect 209044 298172 209096 298178
rect 209044 298114 209096 298120
rect 209412 298172 209464 298178
rect 209412 298114 209464 298120
rect 209044 291848 209096 291854
rect 209044 291790 209096 291796
rect 209056 284172 209084 291790
rect 209424 284172 209452 298114
rect 209962 292632 210018 292641
rect 209962 292567 210018 292576
rect 209976 284172 210004 292567
rect 210436 286278 210464 345034
rect 210516 311160 210568 311166
rect 210516 311102 210568 311108
rect 210528 292913 210556 311102
rect 210514 292904 210570 292913
rect 210514 292839 210570 292848
rect 210424 286272 210476 286278
rect 210424 286214 210476 286220
rect 210528 284172 210556 292839
rect 211436 286272 211488 286278
rect 211436 286214 211488 286220
rect 210882 284336 210938 284345
rect 210882 284271 210938 284280
rect 210896 284172 210924 284271
rect 205362 283928 205418 283937
rect 204732 283886 205362 283914
rect 200026 282976 200082 282985
rect 200132 282962 200160 283886
rect 211448 283914 211476 286214
rect 211816 285734 211844 374002
rect 321558 371376 321614 371385
rect 321558 371311 321614 371320
rect 258080 371272 258132 371278
rect 258080 371214 258132 371220
rect 242164 369980 242216 369986
rect 242164 369922 242216 369928
rect 231124 369912 231176 369918
rect 231124 369854 231176 369860
rect 214564 365832 214616 365838
rect 214564 365774 214616 365780
rect 212906 363624 212962 363633
rect 212906 363559 212962 363568
rect 211896 329180 211948 329186
rect 211896 329122 211948 329128
rect 211908 306374 211936 329122
rect 211908 306346 212120 306374
rect 211986 287600 212042 287609
rect 211986 287535 212042 287544
rect 211804 285728 211856 285734
rect 211804 285670 211856 285676
rect 212000 284172 212028 287535
rect 212092 284186 212120 306346
rect 212354 284472 212410 284481
rect 212354 284407 212410 284416
rect 212368 284186 212396 284407
rect 212092 284172 212396 284186
rect 212920 284172 212948 363559
rect 213642 298752 213698 298761
rect 213642 298687 213698 298696
rect 213458 291408 213514 291417
rect 213458 291343 213514 291352
rect 213472 284172 213500 291343
rect 213656 290465 213684 298687
rect 213826 291816 213882 291825
rect 213826 291751 213882 291760
rect 213840 291417 213868 291751
rect 213826 291408 213882 291417
rect 213826 291343 213882 291352
rect 213642 290456 213698 290465
rect 213642 290391 213698 290400
rect 213828 285728 213880 285734
rect 213828 285670 213880 285676
rect 213840 284172 213868 285670
rect 214576 284186 214604 365774
rect 224224 365764 224276 365770
rect 224224 365706 224276 365712
rect 214656 363044 214708 363050
rect 214656 362986 214708 362992
rect 214668 309126 214696 362986
rect 218242 361856 218298 361865
rect 218242 361791 218298 361800
rect 216036 343732 216088 343738
rect 216036 343674 216088 343680
rect 215944 331288 215996 331294
rect 215944 331230 215996 331236
rect 215852 318776 215904 318782
rect 215852 318718 215904 318724
rect 215864 317490 215892 318718
rect 215852 317484 215904 317490
rect 215852 317426 215904 317432
rect 214656 309120 214708 309126
rect 214656 309062 214708 309068
rect 215208 309120 215260 309126
rect 215208 309062 215260 309068
rect 215220 307834 215248 309062
rect 215208 307828 215260 307834
rect 215208 307770 215260 307776
rect 215220 286657 215248 307770
rect 215298 294128 215354 294137
rect 215298 294063 215354 294072
rect 215312 293185 215340 294063
rect 215298 293176 215354 293185
rect 215298 293111 215354 293120
rect 215298 292632 215354 292641
rect 215298 292567 215354 292576
rect 215206 286648 215262 286657
rect 215206 286583 215262 286592
rect 214746 284336 214802 284345
rect 214746 284271 214802 284280
rect 214760 284186 214788 284271
rect 214576 284172 214788 284186
rect 215312 284172 215340 292567
rect 215864 284172 215892 317426
rect 215956 292641 215984 331230
rect 216048 318782 216076 343674
rect 216036 318776 216088 318782
rect 216036 318718 216088 318724
rect 216954 292904 217010 292913
rect 216954 292839 217010 292848
rect 216968 292641 216996 292839
rect 215942 292632 215998 292641
rect 215942 292567 215998 292576
rect 216954 292632 217010 292641
rect 216954 292567 217010 292576
rect 217322 288688 217378 288697
rect 217322 288623 217378 288632
rect 216770 284608 216826 284617
rect 216770 284543 216826 284552
rect 216784 284442 216812 284543
rect 216772 284436 216824 284442
rect 216772 284378 216824 284384
rect 216784 284172 216812 284378
rect 217336 284172 217364 288623
rect 218256 284172 218284 361791
rect 222842 361720 222898 361729
rect 222842 361655 222898 361664
rect 220082 342408 220138 342417
rect 220082 342343 220138 342352
rect 218702 320240 218758 320249
rect 218702 320175 218758 320184
rect 218716 311166 218744 320175
rect 218704 311160 218756 311166
rect 218704 311102 218756 311108
rect 218612 291236 218664 291242
rect 218612 291178 218664 291184
rect 218624 284172 218652 291178
rect 219162 286104 219218 286113
rect 219162 286039 219218 286048
rect 219176 284172 219204 286039
rect 220096 285954 220124 342343
rect 220174 338464 220230 338473
rect 220174 338399 220230 338408
rect 220188 295497 220216 338399
rect 220820 323672 220872 323678
rect 220820 323614 220872 323620
rect 220174 295488 220230 295497
rect 220174 295423 220230 295432
rect 220726 295488 220782 295497
rect 220726 295423 220782 295432
rect 220176 292596 220228 292602
rect 220176 292538 220228 292544
rect 220004 285938 220124 285954
rect 220004 285932 220136 285938
rect 220004 285926 220084 285932
rect 220004 284186 220032 285926
rect 220084 285874 220136 285880
rect 220082 285832 220138 285841
rect 220082 285767 220138 285776
rect 212092 284158 212382 284172
rect 214576 284158 214774 284172
rect 219742 284158 220032 284186
rect 220096 284172 220124 285767
rect 220188 284050 220216 292538
rect 220740 285734 220768 295423
rect 220728 285728 220780 285734
rect 220728 285670 220780 285676
rect 220726 284064 220782 284073
rect 220188 284022 220726 284050
rect 220726 283999 220782 284008
rect 211618 283928 211674 283937
rect 211448 283900 211618 283914
rect 211462 283886 211618 283900
rect 205362 283863 205418 283872
rect 214470 283928 214526 283937
rect 214406 283886 214470 283914
rect 211618 283863 211674 283872
rect 214470 283863 214526 283872
rect 215942 283928 215998 283937
rect 217414 283928 217470 283937
rect 215998 283886 216246 283914
rect 215942 283863 215998 283872
rect 220832 283914 220860 323614
rect 222856 304298 222884 361655
rect 222934 332616 222990 332625
rect 222934 332551 222990 332560
rect 222844 304292 222896 304298
rect 222844 304234 222896 304240
rect 222948 302326 222976 332551
rect 223026 319424 223082 319433
rect 223026 319359 223082 319368
rect 222936 302320 222988 302326
rect 222936 302262 222988 302268
rect 222200 294024 222252 294030
rect 222200 293966 222252 293972
rect 221554 286648 221610 286657
rect 221554 286583 221610 286592
rect 221568 284172 221596 286583
rect 222108 285728 222160 285734
rect 222108 285670 222160 285676
rect 222120 284172 222148 285670
rect 222212 285326 222240 293966
rect 223040 291718 223068 319359
rect 223488 302320 223540 302326
rect 223488 302262 223540 302268
rect 222476 291712 222528 291718
rect 222476 291654 222528 291660
rect 223028 291712 223080 291718
rect 223028 291654 223080 291660
rect 222200 285320 222252 285326
rect 222200 285262 222252 285268
rect 222488 284172 222516 291654
rect 223040 291310 223068 291654
rect 223028 291304 223080 291310
rect 223028 291246 223080 291252
rect 223500 285841 223528 302262
rect 223580 287156 223632 287162
rect 223580 287098 223632 287104
rect 223486 285832 223542 285841
rect 223486 285767 223542 285776
rect 222660 285320 222712 285326
rect 222660 285262 222712 285268
rect 222672 284186 222700 285262
rect 222672 284158 223054 284186
rect 223592 284050 223620 287098
rect 224236 286414 224264 365706
rect 226984 360256 227036 360262
rect 226984 360198 227036 360204
rect 225604 357468 225656 357474
rect 225604 357410 225656 357416
rect 225052 313948 225104 313954
rect 225052 313890 225104 313896
rect 224314 295352 224370 295361
rect 224314 295287 224370 295296
rect 224224 286408 224276 286414
rect 224224 286350 224276 286356
rect 224328 285705 224356 295287
rect 224500 288516 224552 288522
rect 224500 288458 224552 288464
rect 223946 285696 224002 285705
rect 223946 285631 224002 285640
rect 224314 285696 224370 285705
rect 224314 285631 224370 285640
rect 223960 284172 223988 285631
rect 223762 284064 223818 284073
rect 223592 284036 223762 284050
rect 223606 284022 223762 284036
rect 223762 283999 223818 284008
rect 221278 283928 221334 283937
rect 217470 283886 217718 283914
rect 220832 283886 221278 283914
rect 217414 283863 217470 283872
rect 224512 283914 224540 288458
rect 224682 283928 224738 283937
rect 224512 283900 224682 283914
rect 224526 283886 224682 283900
rect 221278 283863 221334 283872
rect 225064 283914 225092 313890
rect 225616 298761 225644 357410
rect 225972 300144 226024 300150
rect 225972 300086 226024 300092
rect 225602 298752 225658 298761
rect 225602 298687 225658 298696
rect 225418 285696 225474 285705
rect 225418 285631 225474 285640
rect 225432 284172 225460 285631
rect 225984 284172 226012 300086
rect 226996 288697 227024 360198
rect 227442 352064 227498 352073
rect 227442 351999 227498 352008
rect 227076 318096 227128 318102
rect 227076 318038 227128 318044
rect 227088 299538 227116 318038
rect 227076 299532 227128 299538
rect 227076 299474 227128 299480
rect 226982 288688 227038 288697
rect 226982 288623 227038 288632
rect 226522 285832 226578 285841
rect 226522 285767 226578 285776
rect 226536 284172 226564 285767
rect 226996 284186 227024 288623
rect 226918 284158 227024 284186
rect 227456 284172 227484 351999
rect 229192 345160 229244 345166
rect 229192 345102 229244 345108
rect 228364 330540 228416 330546
rect 228364 330482 228416 330488
rect 227812 294024 227864 294030
rect 227812 293966 227864 293972
rect 227824 284172 227852 293966
rect 227902 290456 227958 290465
rect 227902 290391 227958 290400
rect 227916 284186 227944 290391
rect 228376 286657 228404 330482
rect 228456 326392 228508 326398
rect 228456 326334 228508 326340
rect 228468 294030 228496 326334
rect 229204 306374 229232 345102
rect 230478 326360 230534 326369
rect 230478 326295 230534 326304
rect 230492 322522 230520 326295
rect 230480 322516 230532 322522
rect 230480 322458 230532 322464
rect 230480 311228 230532 311234
rect 230480 311170 230532 311176
rect 229204 306346 229416 306374
rect 228916 299532 228968 299538
rect 228916 299474 228968 299480
rect 228456 294024 228508 294030
rect 228456 293966 228508 293972
rect 228362 286648 228418 286657
rect 228362 286583 228418 286592
rect 227916 284158 228390 284186
rect 228928 284172 228956 299474
rect 229284 286408 229336 286414
rect 229284 286350 229336 286356
rect 229296 284172 229324 286350
rect 225234 283928 225290 283937
rect 225064 283900 225234 283914
rect 225078 283886 225234 283900
rect 224682 283863 224738 283872
rect 229388 283914 229416 306346
rect 229742 294128 229798 294137
rect 229742 294063 229798 294072
rect 229756 287065 229784 294063
rect 229742 287056 229798 287065
rect 229742 286991 229798 287000
rect 230386 286648 230442 286657
rect 230386 286583 230442 286592
rect 230112 286408 230164 286414
rect 230112 286350 230164 286356
rect 230124 285802 230152 286350
rect 230112 285796 230164 285802
rect 230112 285738 230164 285744
rect 230400 284172 230428 286583
rect 230492 284442 230520 311170
rect 231136 292602 231164 369854
rect 238024 364472 238076 364478
rect 238024 364414 238076 364420
rect 231216 356176 231268 356182
rect 231216 356118 231268 356124
rect 231228 309126 231256 356118
rect 236644 349172 236696 349178
rect 236644 349114 236696 349120
rect 233974 332752 234030 332761
rect 233974 332687 234030 332696
rect 232504 322244 232556 322250
rect 232504 322186 232556 322192
rect 231216 309120 231268 309126
rect 231216 309062 231268 309068
rect 232516 306474 232544 322186
rect 233884 320884 233936 320890
rect 233884 320826 233936 320832
rect 232504 306468 232556 306474
rect 232504 306410 232556 306416
rect 232516 306374 232544 306410
rect 232240 306346 232544 306374
rect 231124 292596 231176 292602
rect 231124 292538 231176 292544
rect 230754 288824 230810 288833
rect 230754 288759 230810 288768
rect 230768 287162 230796 288759
rect 230756 287156 230808 287162
rect 230756 287098 230808 287104
rect 230480 284436 230532 284442
rect 230480 284378 230532 284384
rect 230768 284172 230796 287098
rect 231308 287088 231360 287094
rect 231308 287030 231360 287036
rect 230110 283928 230166 283937
rect 229388 283886 230110 283914
rect 225234 283863 225290 283872
rect 231320 283914 231348 287030
rect 231676 284436 231728 284442
rect 231676 284378 231728 284384
rect 231688 284172 231716 284378
rect 232240 284172 232268 306346
rect 232504 304292 232556 304298
rect 232504 304234 232556 304240
rect 232516 285705 232544 304234
rect 233698 295352 233754 295361
rect 233698 295287 233754 295296
rect 233148 292596 233200 292602
rect 233148 292538 233200 292544
rect 232778 291544 232834 291553
rect 232778 291479 232834 291488
rect 232502 285696 232558 285705
rect 232502 285631 232558 285640
rect 232792 284172 232820 291479
rect 233160 284172 233188 292538
rect 233712 284172 233740 295287
rect 233896 287162 233924 320826
rect 233988 305862 234016 332687
rect 235264 320952 235316 320958
rect 235264 320894 235316 320900
rect 233976 305856 234028 305862
rect 233976 305798 234028 305804
rect 234528 305856 234580 305862
rect 234528 305798 234580 305804
rect 234540 305114 234568 305798
rect 234528 305108 234580 305114
rect 234528 305050 234580 305056
rect 233974 302832 234030 302841
rect 233974 302767 234030 302776
rect 233988 295361 234016 302767
rect 233974 295352 234030 295361
rect 233974 295287 234030 295296
rect 233884 287156 233936 287162
rect 233884 287098 233936 287104
rect 233896 284186 233924 287098
rect 234540 287054 234568 305050
rect 235276 298081 235304 320894
rect 235538 298752 235594 298761
rect 235538 298687 235594 298696
rect 235262 298072 235318 298081
rect 235262 298007 235318 298016
rect 234540 287026 234752 287054
rect 234618 285696 234674 285705
rect 234618 285631 234674 285640
rect 233896 284158 234278 284186
rect 234632 284172 234660 285631
rect 234724 284186 234752 287026
rect 234724 284158 235198 284186
rect 235552 284172 235580 298687
rect 236182 298072 236238 298081
rect 236182 298007 236238 298016
rect 236196 296857 236224 298007
rect 236182 296848 236238 296857
rect 236182 296783 236238 296792
rect 236000 293276 236052 293282
rect 236000 293218 236052 293224
rect 236012 285705 236040 293218
rect 236092 291236 236144 291242
rect 236092 291178 236144 291184
rect 235998 285696 236054 285705
rect 235998 285631 236054 285640
rect 236104 284172 236132 291178
rect 236196 284186 236224 296783
rect 236656 291242 236684 349114
rect 236736 322516 236788 322522
rect 236736 322458 236788 322464
rect 236748 315382 236776 322458
rect 236736 315376 236788 315382
rect 236736 315318 236788 315324
rect 236736 309120 236788 309126
rect 236736 309062 236788 309068
rect 236644 291236 236696 291242
rect 236644 291178 236696 291184
rect 236748 286385 236776 309062
rect 238036 289134 238064 364414
rect 238116 364404 238168 364410
rect 238116 364346 238168 364352
rect 238128 293962 238156 364346
rect 240232 361616 240284 361622
rect 240232 361558 240284 361564
rect 238760 358828 238812 358834
rect 238760 358770 238812 358776
rect 238772 304314 238800 358770
rect 238680 304298 238800 304314
rect 238668 304292 238800 304298
rect 238720 304286 238800 304292
rect 238668 304234 238720 304240
rect 238116 293956 238168 293962
rect 238116 293898 238168 293904
rect 238024 289128 238076 289134
rect 238024 289070 238076 289076
rect 238114 287464 238170 287473
rect 238114 287399 238170 287408
rect 236734 286376 236790 286385
rect 236734 286311 236790 286320
rect 237564 285864 237616 285870
rect 237564 285806 237616 285812
rect 236196 284158 236670 284186
rect 237576 284172 237604 285806
rect 238128 284172 238156 287399
rect 238680 285870 238708 304234
rect 240244 294545 240272 361558
rect 241242 330168 241298 330177
rect 241242 330103 241298 330112
rect 241256 329186 241284 330103
rect 241244 329180 241296 329186
rect 241244 329122 241296 329128
rect 240782 315344 240838 315353
rect 240782 315279 240838 315288
rect 240796 299577 240824 315279
rect 241428 300960 241480 300966
rect 241428 300902 241480 300908
rect 240782 299568 240838 299577
rect 240782 299503 240838 299512
rect 240796 296714 240824 299503
rect 240796 296686 240916 296714
rect 240784 296064 240836 296070
rect 240784 296006 240836 296012
rect 240230 294536 240286 294545
rect 240230 294471 240286 294480
rect 240244 294137 240272 294471
rect 239034 294128 239090 294137
rect 239034 294063 239090 294072
rect 240230 294128 240286 294137
rect 240230 294063 240286 294072
rect 238668 285864 238720 285870
rect 238668 285806 238720 285812
rect 239048 284172 239076 294063
rect 240508 293956 240560 293962
rect 240508 293898 240560 293904
rect 239954 287328 240010 287337
rect 239954 287263 240010 287272
rect 239586 285832 239642 285841
rect 239586 285767 239642 285776
rect 239600 284172 239628 285767
rect 239968 284172 239996 287263
rect 240520 284172 240548 293898
rect 240796 285705 240824 296006
rect 240782 285696 240838 285705
rect 240782 285631 240838 285640
rect 240888 284172 240916 296686
rect 241440 284172 241468 300902
rect 242176 285569 242204 369922
rect 248418 368520 248474 368529
rect 248418 368455 248474 368464
rect 246302 354784 246358 354793
rect 246302 354719 246358 354728
rect 242254 346760 242310 346769
rect 242254 346695 242310 346704
rect 242268 294681 242296 346695
rect 244094 328536 244150 328545
rect 244094 328471 244150 328480
rect 242900 315376 242952 315382
rect 242900 315318 242952 315324
rect 242254 294672 242310 294681
rect 242254 294607 242310 294616
rect 242348 289128 242400 289134
rect 242348 289070 242400 289076
rect 242360 288522 242388 289070
rect 242348 288516 242400 288522
rect 242348 288458 242400 288464
rect 242360 287054 242388 288458
rect 242268 287026 242388 287054
rect 242162 285560 242218 285569
rect 242162 285495 242218 285504
rect 242268 284186 242296 287026
rect 242622 285560 242678 285569
rect 242622 285495 242678 285504
rect 242636 284186 242664 285495
rect 242006 284158 242296 284186
rect 242374 284158 242664 284186
rect 242912 284172 242940 315318
rect 243818 285696 243874 285705
rect 243818 285631 243874 285640
rect 243832 284172 243860 285631
rect 243912 284368 243964 284374
rect 243912 284310 243964 284316
rect 243634 284064 243690 284073
rect 243478 284022 243634 284050
rect 243634 283999 243690 284008
rect 231582 283928 231638 283937
rect 231320 283900 231582 283914
rect 231334 283886 231582 283900
rect 230110 283863 230166 283872
rect 231582 283863 231638 283872
rect 236734 283928 236790 283937
rect 238666 283928 238722 283937
rect 236790 283886 237038 283914
rect 238510 283886 238666 283914
rect 236734 283863 236790 283872
rect 238666 283863 238722 283872
rect 200082 282934 200160 282962
rect 200026 282911 200082 282920
rect 199474 282840 199530 282849
rect 199474 282775 199530 282784
rect 199384 276684 199436 276690
rect 199384 276626 199436 276632
rect 200040 274582 200068 274613
rect 200028 274576 200080 274582
rect 200026 274544 200028 274553
rect 200080 274544 200082 274553
rect 200026 274479 200082 274488
rect 199382 270192 199438 270201
rect 199382 270127 199438 270136
rect 198832 244316 198884 244322
rect 198832 244258 198884 244264
rect 198738 241496 198794 241505
rect 198738 241431 198794 241440
rect 198752 240378 198780 241431
rect 198740 240372 198792 240378
rect 198740 240314 198792 240320
rect 198844 240281 198872 244258
rect 198830 240272 198886 240281
rect 198830 240207 198886 240216
rect 198648 240168 198700 240174
rect 198648 240110 198700 240116
rect 199396 229022 199424 270127
rect 199476 261520 199528 261526
rect 199476 261462 199528 261468
rect 199488 237862 199516 261462
rect 199566 256592 199622 256601
rect 199566 256527 199622 256536
rect 199580 247722 199608 256527
rect 199568 247716 199620 247722
rect 199568 247658 199620 247664
rect 199568 240780 199620 240786
rect 199568 240722 199620 240728
rect 199476 237856 199528 237862
rect 199476 237798 199528 237804
rect 199580 231742 199608 240722
rect 199936 237856 199988 237862
rect 199936 237798 199988 237804
rect 199568 231736 199620 231742
rect 199568 231678 199620 231684
rect 199384 229016 199436 229022
rect 199384 228958 199436 228964
rect 199396 214674 199424 228958
rect 199476 222964 199528 222970
rect 199476 222906 199528 222912
rect 199488 219337 199516 222906
rect 199474 219328 199530 219337
rect 199474 219263 199530 219272
rect 199384 214668 199436 214674
rect 199384 214610 199436 214616
rect 197360 214600 197412 214606
rect 197360 214542 197412 214548
rect 197372 213926 197400 214542
rect 197360 213920 197412 213926
rect 197360 213862 197412 213868
rect 198002 212664 198058 212673
rect 198002 212599 198058 212608
rect 197912 209840 197964 209846
rect 197912 209782 197964 209788
rect 197924 208350 197952 209782
rect 197912 208344 197964 208350
rect 197912 208286 197964 208292
rect 198016 193186 198044 212599
rect 198278 211168 198334 211177
rect 198278 211103 198334 211112
rect 198004 193180 198056 193186
rect 198004 193122 198056 193128
rect 197268 192568 197320 192574
rect 197268 192510 197320 192516
rect 198002 184240 198058 184249
rect 198002 184175 198058 184184
rect 196898 181520 196954 181529
rect 196898 181455 196954 181464
rect 196808 178084 196860 178090
rect 196808 178026 196860 178032
rect 196820 166938 196848 178026
rect 196808 166932 196860 166938
rect 196808 166874 196860 166880
rect 196808 125724 196860 125730
rect 196808 125666 196860 125672
rect 196714 87544 196770 87553
rect 196714 87479 196770 87488
rect 196820 85474 196848 125666
rect 196808 85468 196860 85474
rect 196808 85410 196860 85416
rect 198016 11830 198044 184175
rect 198188 135924 198240 135930
rect 198188 135866 198240 135872
rect 198094 133104 198150 133113
rect 198094 133039 198150 133048
rect 198004 11824 198056 11830
rect 198004 11766 198056 11772
rect 196622 3496 196678 3505
rect 196622 3431 196678 3440
rect 198108 2174 198136 133039
rect 198200 30977 198228 135866
rect 198292 123457 198320 211103
rect 199948 178702 199976 237798
rect 200040 207738 200068 274479
rect 243924 267734 243952 284310
rect 244108 284073 244136 328471
rect 245752 315308 245804 315314
rect 245752 315250 245804 315256
rect 244280 312588 244332 312594
rect 244280 312530 244332 312536
rect 244188 287156 244240 287162
rect 244188 287098 244240 287104
rect 244094 284064 244150 284073
rect 244094 283999 244150 284008
rect 244108 282985 244136 283999
rect 244200 283898 244228 287098
rect 244188 283892 244240 283898
rect 244188 283834 244240 283840
rect 244094 282976 244150 282985
rect 244094 282911 244150 282920
rect 244292 274553 244320 312530
rect 244556 309800 244608 309806
rect 244556 309742 244608 309748
rect 244464 295996 244516 296002
rect 244464 295938 244516 295944
rect 244372 288448 244424 288454
rect 244372 288390 244424 288396
rect 244278 274544 244334 274553
rect 244278 274479 244334 274488
rect 243924 267706 244044 267734
rect 244016 259321 244044 267706
rect 244002 259312 244058 259321
rect 244002 259247 244058 259256
rect 244384 253065 244412 288390
rect 244476 259593 244504 295938
rect 244568 280265 244596 309742
rect 245108 296744 245160 296750
rect 245108 296686 245160 296692
rect 245120 296002 245148 296686
rect 245108 295996 245160 296002
rect 245108 295938 245160 295944
rect 244554 280256 244610 280265
rect 244554 280191 244610 280200
rect 245474 280256 245530 280265
rect 245474 280191 245476 280200
rect 245528 280191 245530 280200
rect 245476 280162 245528 280168
rect 245660 278996 245712 279002
rect 245660 278938 245712 278944
rect 245672 278905 245700 278938
rect 245658 278896 245714 278905
rect 245658 278831 245714 278840
rect 245764 276729 245792 315250
rect 246316 297498 246344 354719
rect 247040 336864 247092 336870
rect 247040 336806 247092 336812
rect 246396 298784 246448 298790
rect 246396 298726 246448 298732
rect 246304 297492 246356 297498
rect 246304 297434 246356 297440
rect 245844 294636 245896 294642
rect 245844 294578 245896 294584
rect 245750 276720 245806 276729
rect 245750 276655 245752 276664
rect 245804 276655 245806 276664
rect 245752 276626 245804 276632
rect 245764 276595 245792 276626
rect 245658 273728 245714 273737
rect 245658 273663 245714 273672
rect 245672 273290 245700 273663
rect 245856 273306 245884 294578
rect 246120 285796 246172 285802
rect 246120 285738 246172 285744
rect 245936 282872 245988 282878
rect 245936 282814 245988 282820
rect 245948 281625 245976 282814
rect 245934 281616 245990 281625
rect 245934 281551 245990 281560
rect 245934 281072 245990 281081
rect 245934 281007 245990 281016
rect 245948 280838 245976 281007
rect 245936 280832 245988 280838
rect 245936 280774 245988 280780
rect 245936 279472 245988 279478
rect 245934 279440 245936 279449
rect 245988 279440 245990 279449
rect 245934 279375 245990 279384
rect 245936 278112 245988 278118
rect 245934 278080 245936 278089
rect 245988 278080 245990 278089
rect 245934 278015 245990 278024
rect 246028 278044 246080 278050
rect 246028 277986 246080 277992
rect 246040 277545 246068 277986
rect 246026 277536 246082 277545
rect 246026 277471 246082 277480
rect 246132 277394 246160 285738
rect 246302 283248 246358 283257
rect 246302 283183 246304 283192
rect 246356 283183 246358 283192
rect 246304 283154 246356 283160
rect 246040 277366 246160 277394
rect 245936 276004 245988 276010
rect 245936 275946 245988 275952
rect 245948 275913 245976 275946
rect 245934 275904 245990 275913
rect 245934 275839 245990 275848
rect 245660 273284 245712 273290
rect 245856 273278 245976 273306
rect 245660 273226 245712 273232
rect 245842 273184 245898 273193
rect 245842 273119 245898 273128
rect 245856 271930 245884 273119
rect 245844 271924 245896 271930
rect 245844 271866 245896 271872
rect 245842 271552 245898 271561
rect 245842 271487 245898 271496
rect 245856 270570 245884 271487
rect 245844 270564 245896 270570
rect 245844 270506 245896 270512
rect 245844 269816 245896 269822
rect 245844 269758 245896 269764
rect 245752 269068 245804 269074
rect 245752 269010 245804 269016
rect 245764 268025 245792 269010
rect 245750 268016 245806 268025
rect 245750 267951 245806 267960
rect 245856 267734 245884 269758
rect 245948 269657 245976 273278
rect 245934 269648 245990 269657
rect 245934 269583 245990 269592
rect 245764 267706 245884 267734
rect 245764 265305 245792 267706
rect 245948 267594 245976 269583
rect 245856 267566 245976 267594
rect 245856 267034 245884 267566
rect 245934 267472 245990 267481
rect 245934 267407 245990 267416
rect 245844 267028 245896 267034
rect 245844 266970 245896 266976
rect 245948 266422 245976 267407
rect 245936 266416 245988 266422
rect 245936 266358 245988 266364
rect 245934 265840 245990 265849
rect 245934 265775 245990 265784
rect 245948 265674 245976 265775
rect 245936 265668 245988 265674
rect 245936 265610 245988 265616
rect 245750 265296 245806 265305
rect 245750 265231 245806 265240
rect 244554 264480 244610 264489
rect 244554 264415 244610 264424
rect 244462 259584 244518 259593
rect 244462 259519 244518 259528
rect 244476 259486 244504 259519
rect 244464 259480 244516 259486
rect 244464 259422 244516 259428
rect 244370 253056 244426 253065
rect 244370 252991 244426 253000
rect 244002 248432 244058 248441
rect 244002 248367 244058 248376
rect 243910 240544 243966 240553
rect 243910 240479 243966 240488
rect 200118 240408 200174 240417
rect 200118 240343 200174 240352
rect 200132 240310 200160 240343
rect 200120 240304 200172 240310
rect 200120 240246 200172 240252
rect 200120 240168 200172 240174
rect 200120 240110 200172 240116
rect 200132 237454 200160 240110
rect 200120 237448 200172 237454
rect 200120 237390 200172 237396
rect 200224 223009 200252 240244
rect 200304 240168 200356 240174
rect 200304 240110 200356 240116
rect 200316 229809 200344 240110
rect 200592 239737 200620 240244
rect 200946 240136 201002 240145
rect 200946 240071 201002 240080
rect 200578 239728 200634 239737
rect 200578 239663 200634 239672
rect 200302 229800 200358 229809
rect 200302 229735 200358 229744
rect 200960 229094 200988 240071
rect 201144 238754 201172 240244
rect 201052 238726 201172 238754
rect 201052 237862 201080 238726
rect 201040 237856 201092 237862
rect 201040 237798 201092 237804
rect 200960 229066 201172 229094
rect 200210 223000 200266 223009
rect 200210 222935 200266 222944
rect 200028 207732 200080 207738
rect 200028 207674 200080 207680
rect 199936 178696 199988 178702
rect 199936 178638 199988 178644
rect 201144 178022 201172 229066
rect 201512 228721 201540 240244
rect 202064 238649 202092 240244
rect 202144 240168 202196 240174
rect 202144 240110 202196 240116
rect 202050 238640 202106 238649
rect 202050 238575 202106 238584
rect 201592 237448 201644 237454
rect 201592 237390 201644 237396
rect 201604 233889 201632 237390
rect 201590 233880 201646 233889
rect 201590 233815 201646 233824
rect 202156 229090 202184 240110
rect 202616 238754 202644 240244
rect 202248 238726 202644 238754
rect 202248 238241 202276 238726
rect 202234 238232 202290 238241
rect 202234 238167 202290 238176
rect 202144 229084 202196 229090
rect 202144 229026 202196 229032
rect 201498 228712 201554 228721
rect 201498 228647 201554 228656
rect 201512 220114 201540 228647
rect 201500 220108 201552 220114
rect 201500 220050 201552 220056
rect 202142 199472 202198 199481
rect 202142 199407 202198 199416
rect 201132 178016 201184 178022
rect 201132 177958 201184 177964
rect 200764 142860 200816 142866
rect 200764 142802 200816 142808
rect 199382 134192 199438 134201
rect 199382 134127 199438 134136
rect 198278 123448 198334 123457
rect 198278 123383 198334 123392
rect 199396 63510 199424 134127
rect 199476 121576 199528 121582
rect 199476 121518 199528 121524
rect 199488 88330 199516 121518
rect 200776 89185 200804 142802
rect 200856 109132 200908 109138
rect 200856 109074 200908 109080
rect 200762 89176 200818 89185
rect 200762 89111 200818 89120
rect 199476 88324 199528 88330
rect 199476 88266 199528 88272
rect 200868 64870 200896 109074
rect 200856 64864 200908 64870
rect 200856 64806 200908 64812
rect 199384 63504 199436 63510
rect 199384 63446 199436 63452
rect 200764 36644 200816 36650
rect 200764 36586 200816 36592
rect 198186 30968 198242 30977
rect 198186 30903 198242 30912
rect 200776 3369 200804 36586
rect 202156 3534 202184 199407
rect 202248 198014 202276 238167
rect 202786 222864 202842 222873
rect 202786 222799 202842 222808
rect 202236 198008 202288 198014
rect 202236 197950 202288 197956
rect 202800 192506 202828 222799
rect 202984 213994 203012 240244
rect 203536 238754 203564 240244
rect 203076 238726 203564 238754
rect 203076 222873 203104 238726
rect 204088 234433 204116 240244
rect 204456 235958 204484 240244
rect 204902 239728 204958 239737
rect 204902 239663 204958 239672
rect 204444 235952 204496 235958
rect 204444 235894 204496 235900
rect 203522 234424 203578 234433
rect 203522 234359 203578 234368
rect 204074 234424 204130 234433
rect 204074 234359 204130 234368
rect 203062 222864 203118 222873
rect 203062 222799 203118 222808
rect 203340 214600 203392 214606
rect 203340 214542 203392 214548
rect 202972 213988 203024 213994
rect 202972 213930 203024 213936
rect 203352 212537 203380 214542
rect 203338 212528 203394 212537
rect 203338 212463 203394 212472
rect 202788 192500 202840 192506
rect 202788 192442 202840 192448
rect 203536 187241 203564 234359
rect 204810 220824 204866 220833
rect 204810 220759 204866 220768
rect 204824 219473 204852 220759
rect 204810 219464 204866 219473
rect 204810 219399 204866 219408
rect 204824 218793 204852 219399
rect 204810 218784 204866 218793
rect 204810 218719 204866 218728
rect 203616 213988 203668 213994
rect 203616 213930 203668 213936
rect 203628 195294 203656 213930
rect 204916 209166 204944 239663
rect 205008 226137 205036 240244
rect 204994 226128 205050 226137
rect 204994 226063 205050 226072
rect 205008 222902 205036 226063
rect 204996 222896 205048 222902
rect 204996 222838 205048 222844
rect 205376 220833 205404 240244
rect 205362 220824 205418 220833
rect 205362 220759 205418 220768
rect 204994 216200 205050 216209
rect 204994 216135 205050 216144
rect 204904 209160 204956 209166
rect 204904 209102 204956 209108
rect 205008 198665 205036 216135
rect 205548 209092 205600 209098
rect 205548 209034 205600 209040
rect 205560 208894 205588 209034
rect 205548 208888 205600 208894
rect 205548 208830 205600 208836
rect 204994 198656 205050 198665
rect 204994 198591 205050 198600
rect 203616 195288 203668 195294
rect 203616 195230 203668 195236
rect 203522 187232 203578 187241
rect 203522 187167 203578 187176
rect 203616 180872 203668 180878
rect 203616 180814 203668 180820
rect 203524 176724 203576 176730
rect 203524 176666 203576 176672
rect 203536 149734 203564 176666
rect 203628 173806 203656 180814
rect 205560 177954 205588 208830
rect 205928 207097 205956 240244
rect 206480 208894 206508 240244
rect 206848 237454 206876 240244
rect 206836 237448 206888 237454
rect 206836 237390 206888 237396
rect 207400 218113 207428 240244
rect 207952 239601 207980 240244
rect 207938 239592 207994 239601
rect 207938 239527 207994 239536
rect 207952 237454 207980 239527
rect 207664 237448 207716 237454
rect 207664 237390 207716 237396
rect 207940 237448 207992 237454
rect 207940 237390 207992 237396
rect 207676 230450 207704 237390
rect 207664 230444 207716 230450
rect 207664 230386 207716 230392
rect 207386 218104 207442 218113
rect 207386 218039 207442 218048
rect 207400 215966 207428 218039
rect 207388 215960 207440 215966
rect 207388 215902 207440 215908
rect 206468 208888 206520 208894
rect 206468 208830 206520 208836
rect 205914 207088 205970 207097
rect 205914 207023 205970 207032
rect 205928 202337 205956 207023
rect 205914 202328 205970 202337
rect 205914 202263 205970 202272
rect 207676 184278 207704 230386
rect 207754 220280 207810 220289
rect 207754 220215 207810 220224
rect 207768 205057 207796 220215
rect 208320 206990 208348 240244
rect 208872 237318 208900 240244
rect 209044 237448 209096 237454
rect 209044 237390 209096 237396
rect 208860 237312 208912 237318
rect 208860 237254 208912 237260
rect 208400 234660 208452 234666
rect 208400 234602 208452 234608
rect 208412 231742 208440 234602
rect 208400 231736 208452 231742
rect 208400 231678 208452 231684
rect 208308 206984 208360 206990
rect 208308 206926 208360 206932
rect 208320 206174 208348 206926
rect 207848 206168 207900 206174
rect 207848 206110 207900 206116
rect 208308 206168 208360 206174
rect 208308 206110 208360 206116
rect 207754 205048 207810 205057
rect 207754 204983 207810 204992
rect 207860 197334 207888 206110
rect 207848 197328 207900 197334
rect 207848 197270 207900 197276
rect 209056 191146 209084 237390
rect 209240 191826 209268 240244
rect 209228 191820 209280 191826
rect 209228 191762 209280 191768
rect 209044 191140 209096 191146
rect 209044 191082 209096 191088
rect 209792 187649 209820 240244
rect 210344 235521 210372 240244
rect 210330 235512 210386 235521
rect 210330 235447 210386 235456
rect 210712 205601 210740 240244
rect 211264 238754 211292 240244
rect 211172 238726 211292 238754
rect 211066 235648 211122 235657
rect 211066 235583 211122 235592
rect 211080 234734 211108 235583
rect 211068 234728 211120 234734
rect 211068 234670 211120 234676
rect 211172 214606 211200 238726
rect 211816 237454 211844 240244
rect 211252 237448 211304 237454
rect 211252 237390 211304 237396
rect 211804 237448 211856 237454
rect 211804 237390 211856 237396
rect 211264 222086 211292 237390
rect 212184 225049 212212 240244
rect 212170 225040 212226 225049
rect 212170 224975 212226 224984
rect 211252 222080 211304 222086
rect 211252 222022 211304 222028
rect 211804 222080 211856 222086
rect 211804 222022 211856 222028
rect 211160 214600 211212 214606
rect 211160 214542 211212 214548
rect 210422 205592 210478 205601
rect 210422 205527 210478 205536
rect 210698 205592 210754 205601
rect 210698 205527 210754 205536
rect 209778 187640 209834 187649
rect 209778 187575 209834 187584
rect 207664 184272 207716 184278
rect 210436 184249 210464 205527
rect 211066 187640 211122 187649
rect 211066 187575 211122 187584
rect 211080 186969 211108 187575
rect 211066 186960 211122 186969
rect 211066 186895 211122 186904
rect 207664 184214 207716 184220
rect 210422 184240 210478 184249
rect 210422 184175 210478 184184
rect 211816 181490 211844 222022
rect 212736 193225 212764 240244
rect 213104 212673 213132 240244
rect 213656 238754 213684 240244
rect 213656 238726 213868 238754
rect 213656 238649 213684 238726
rect 213642 238640 213698 238649
rect 213642 238575 213698 238584
rect 213184 229764 213236 229770
rect 213184 229706 213236 229712
rect 213196 219366 213224 229706
rect 213184 219360 213236 219366
rect 213184 219302 213236 219308
rect 213090 212664 213146 212673
rect 213090 212599 213146 212608
rect 213734 212664 213790 212673
rect 213734 212599 213790 212608
rect 213748 210497 213776 212599
rect 213182 210488 213238 210497
rect 213182 210423 213238 210432
rect 213734 210488 213790 210497
rect 213734 210423 213790 210432
rect 212722 193216 212778 193225
rect 212722 193151 212778 193160
rect 211804 181484 211856 181490
rect 211804 181426 211856 181432
rect 205548 177948 205600 177954
rect 205548 177890 205600 177896
rect 203616 173800 203668 173806
rect 203616 173742 203668 173748
rect 203616 153264 203668 153270
rect 203616 153206 203668 153212
rect 203524 149728 203576 149734
rect 203524 149670 203576 149676
rect 203524 144968 203576 144974
rect 203524 144910 203576 144916
rect 202234 142760 202290 142769
rect 202234 142695 202290 142704
rect 202248 84833 202276 142695
rect 202788 135312 202840 135318
rect 202788 135254 202840 135260
rect 202800 134638 202828 135254
rect 202788 134632 202840 134638
rect 202788 134574 202840 134580
rect 202328 129872 202380 129878
rect 202328 129814 202380 129820
rect 202340 109138 202368 129814
rect 202328 109132 202380 109138
rect 202328 109074 202380 109080
rect 202328 107704 202380 107710
rect 202328 107646 202380 107652
rect 202234 84824 202290 84833
rect 202234 84759 202290 84768
rect 202340 81394 202368 107646
rect 203536 93809 203564 144910
rect 203522 93800 203578 93809
rect 203522 93735 203578 93744
rect 203524 88392 203576 88398
rect 203524 88334 203576 88340
rect 202328 81388 202380 81394
rect 202328 81330 202380 81336
rect 203536 14550 203564 88334
rect 203628 87650 203656 153206
rect 211896 152108 211948 152114
rect 211896 152050 211948 152056
rect 209044 145580 209096 145586
rect 209044 145522 209096 145528
rect 204904 143676 204956 143682
rect 204904 143618 204956 143624
rect 203708 115932 203760 115938
rect 203708 115874 203760 115880
rect 203616 87644 203668 87650
rect 203616 87586 203668 87592
rect 203720 84153 203748 115874
rect 204916 105602 204944 143618
rect 207756 142180 207808 142186
rect 207756 142122 207808 142128
rect 206284 139460 206336 139466
rect 206284 139402 206336 139408
rect 204994 138136 205050 138145
rect 204994 138071 205050 138080
rect 205008 115938 205036 138071
rect 206296 124914 206324 139402
rect 207664 135380 207716 135386
rect 207664 135322 207716 135328
rect 206468 132524 206520 132530
rect 206468 132466 206520 132472
rect 206284 124908 206336 124914
rect 206284 124850 206336 124856
rect 206284 118788 206336 118794
rect 206284 118730 206336 118736
rect 204996 115932 205048 115938
rect 204996 115874 205048 115880
rect 205088 114572 205140 114578
rect 205088 114514 205140 114520
rect 204904 105596 204956 105602
rect 204904 105538 204956 105544
rect 204996 104984 205048 104990
rect 204996 104926 205048 104932
rect 204902 86184 204958 86193
rect 204902 86119 204958 86128
rect 203706 84144 203762 84153
rect 203706 84079 203762 84088
rect 204916 21418 204944 86119
rect 205008 71738 205036 104926
rect 205100 85542 205128 114514
rect 206296 91050 206324 118730
rect 206376 116068 206428 116074
rect 206376 116010 206428 116016
rect 206284 91044 206336 91050
rect 206284 90986 206336 90992
rect 206284 87712 206336 87718
rect 206284 87654 206336 87660
rect 205088 85536 205140 85542
rect 205088 85478 205140 85484
rect 204996 71732 205048 71738
rect 204996 71674 205048 71680
rect 204904 21412 204956 21418
rect 204904 21354 204956 21360
rect 203524 14544 203576 14550
rect 203524 14486 203576 14492
rect 206296 8945 206324 87654
rect 206388 55214 206416 116010
rect 206480 74526 206508 132466
rect 207676 91798 207704 135322
rect 207768 116521 207796 142122
rect 207848 117428 207900 117434
rect 207848 117370 207900 117376
rect 207754 116512 207810 116521
rect 207754 116447 207810 116456
rect 207860 93906 207888 117370
rect 207848 93900 207900 93906
rect 207848 93842 207900 93848
rect 208400 91860 208452 91866
rect 208400 91802 208452 91808
rect 207664 91792 207716 91798
rect 207664 91734 207716 91740
rect 207664 90364 207716 90370
rect 207664 90306 207716 90312
rect 206468 74520 206520 74526
rect 206468 74462 206520 74468
rect 206376 55208 206428 55214
rect 206376 55150 206428 55156
rect 207676 46306 207704 90306
rect 208412 88398 208440 91802
rect 208400 88392 208452 88398
rect 208400 88334 208452 88340
rect 207664 46300 207716 46306
rect 207664 46242 207716 46248
rect 209056 17338 209084 145522
rect 210424 139528 210476 139534
rect 210424 139470 210476 139476
rect 209320 133952 209372 133958
rect 209320 133894 209372 133900
rect 209228 128444 209280 128450
rect 209228 128386 209280 128392
rect 209136 110560 209188 110566
rect 209136 110502 209188 110508
rect 209148 93945 209176 110502
rect 209134 93936 209190 93945
rect 209134 93871 209190 93880
rect 209136 93152 209188 93158
rect 209136 93094 209188 93100
rect 209148 28354 209176 93094
rect 209240 91633 209268 128386
rect 209226 91624 209282 91633
rect 209226 91559 209282 91568
rect 209332 90438 209360 133894
rect 209320 90432 209372 90438
rect 209226 90400 209282 90409
rect 209320 90374 209372 90380
rect 209226 90335 209282 90344
rect 209240 43518 209268 90335
rect 210436 69018 210464 139470
rect 211804 138032 211856 138038
rect 211804 137974 211856 137980
rect 210608 123140 210660 123146
rect 210608 123082 210660 123088
rect 210516 107772 210568 107778
rect 210516 107714 210568 107720
rect 210424 69012 210476 69018
rect 210424 68954 210476 68960
rect 210528 51066 210556 107714
rect 210620 95946 210648 123082
rect 211816 100026 211844 137974
rect 211908 134570 211936 152050
rect 211896 134564 211948 134570
rect 211896 134506 211948 134512
rect 211804 100020 211856 100026
rect 211804 99962 211856 99968
rect 211896 99476 211948 99482
rect 211896 99418 211948 99424
rect 211804 98116 211856 98122
rect 211804 98058 211856 98064
rect 210608 95940 210660 95946
rect 210608 95882 210660 95888
rect 211816 52426 211844 98058
rect 211908 78577 211936 99418
rect 211894 78568 211950 78577
rect 211894 78503 211950 78512
rect 211804 52420 211856 52426
rect 211804 52362 211856 52368
rect 210516 51060 210568 51066
rect 210516 51002 210568 51008
rect 209228 43512 209280 43518
rect 209228 43454 209280 43460
rect 209136 28348 209188 28354
rect 209136 28290 209188 28296
rect 209044 17332 209096 17338
rect 209044 17274 209096 17280
rect 206282 8936 206338 8945
rect 206282 8871 206338 8880
rect 202144 3528 202196 3534
rect 202144 3470 202196 3476
rect 213196 3369 213224 210423
rect 213840 199481 213868 238726
rect 214208 238513 214236 240244
rect 214194 238504 214250 238513
rect 214194 238439 214250 238448
rect 214208 229094 214236 238439
rect 214576 237289 214604 240244
rect 215128 238754 215156 240244
rect 215128 238726 215248 238754
rect 215220 238649 215248 238726
rect 215206 238640 215262 238649
rect 215206 238575 215262 238584
rect 214562 237280 214618 237289
rect 214562 237215 214618 237224
rect 214656 236156 214708 236162
rect 214656 236098 214708 236104
rect 214208 229066 214604 229094
rect 214104 227044 214156 227050
rect 214104 226986 214156 226992
rect 214116 222193 214144 226986
rect 214102 222184 214158 222193
rect 214102 222119 214158 222128
rect 214470 211168 214526 211177
rect 214470 211103 214526 211112
rect 214484 209846 214512 211103
rect 214472 209840 214524 209846
rect 214472 209782 214524 209788
rect 213826 199472 213882 199481
rect 213826 199407 213882 199416
rect 214576 196654 214604 229066
rect 214668 201482 214696 236098
rect 214656 201476 214708 201482
rect 214656 201418 214708 201424
rect 214932 200252 214984 200258
rect 214932 200194 214984 200200
rect 214944 197334 214972 200194
rect 214932 197328 214984 197334
rect 214932 197270 214984 197276
rect 214564 196648 214616 196654
rect 214564 196590 214616 196596
rect 214656 183592 214708 183598
rect 214656 183534 214708 183540
rect 214564 182232 214616 182238
rect 214564 182174 214616 182180
rect 213920 176656 213972 176662
rect 213920 176598 213972 176604
rect 213932 175681 213960 176598
rect 213918 175672 213974 175681
rect 213918 175607 213974 175616
rect 214102 175264 214158 175273
rect 213920 175228 213972 175234
rect 214102 175199 214158 175208
rect 213920 175170 213972 175176
rect 213932 175001 213960 175170
rect 214012 175160 214064 175166
rect 214012 175102 214064 175108
rect 213918 174992 213974 175001
rect 213918 174927 213974 174936
rect 214024 174321 214052 175102
rect 214116 174554 214144 175199
rect 214104 174548 214156 174554
rect 214104 174490 214156 174496
rect 214010 174312 214066 174321
rect 214010 174247 214066 174256
rect 214012 173868 214064 173874
rect 214012 173810 214064 173816
rect 213920 173800 213972 173806
rect 213920 173742 213972 173748
rect 213932 173641 213960 173742
rect 213918 173632 213974 173641
rect 213918 173567 213974 173576
rect 214024 172961 214052 173810
rect 214010 172952 214066 172961
rect 214010 172887 214066 172896
rect 213920 172508 213972 172514
rect 213920 172450 213972 172456
rect 213932 172281 213960 172450
rect 213918 172272 213974 172281
rect 213918 172207 213974 172216
rect 214010 171592 214066 171601
rect 214010 171527 214066 171536
rect 214024 171086 214052 171527
rect 214012 171080 214064 171086
rect 214012 171022 214064 171028
rect 213920 171012 213972 171018
rect 213920 170954 213972 170960
rect 213932 170377 213960 170954
rect 213918 170368 213974 170377
rect 213918 170303 213974 170312
rect 214012 169720 214064 169726
rect 213918 169688 213974 169697
rect 214012 169662 214064 169668
rect 213918 169623 213920 169632
rect 213972 169623 213974 169632
rect 213920 169594 213972 169600
rect 214024 169017 214052 169662
rect 214010 169008 214066 169017
rect 214010 168943 214066 168952
rect 214012 168360 214064 168366
rect 213918 168328 213974 168337
rect 214012 168302 214064 168308
rect 213918 168263 213920 168272
rect 213972 168263 213974 168272
rect 213920 168234 213972 168240
rect 214024 167657 214052 168302
rect 214010 167648 214066 167657
rect 214010 167583 214066 167592
rect 213920 167000 213972 167006
rect 213918 166968 213920 166977
rect 213972 166968 213974 166977
rect 213918 166903 213974 166912
rect 214012 166932 214064 166938
rect 214012 166874 214064 166880
rect 214024 165753 214052 166874
rect 214010 165744 214066 165753
rect 214010 165679 214066 165688
rect 214012 165572 214064 165578
rect 214012 165514 214064 165520
rect 213920 165504 213972 165510
rect 213920 165446 213972 165452
rect 213932 165073 213960 165446
rect 213918 165064 213974 165073
rect 213918 164999 213974 165008
rect 214024 164393 214052 165514
rect 214010 164384 214066 164393
rect 214010 164319 214066 164328
rect 214012 164212 214064 164218
rect 214012 164154 214064 164160
rect 213920 164144 213972 164150
rect 213920 164086 213972 164092
rect 213932 163713 213960 164086
rect 213918 163704 213974 163713
rect 213918 163639 213974 163648
rect 214024 163033 214052 164154
rect 214010 163024 214066 163033
rect 214010 162959 214066 162968
rect 213920 162852 213972 162858
rect 213920 162794 213972 162800
rect 213932 162353 213960 162794
rect 214012 162784 214064 162790
rect 214012 162726 214064 162732
rect 213918 162344 213974 162353
rect 213918 162279 213974 162288
rect 214024 161809 214052 162726
rect 214010 161800 214066 161809
rect 214010 161735 214066 161744
rect 214012 161424 214064 161430
rect 214012 161366 214064 161372
rect 213920 161356 213972 161362
rect 213920 161298 213972 161304
rect 213932 161129 213960 161298
rect 213918 161120 213974 161129
rect 213918 161055 213974 161064
rect 214024 160449 214052 161366
rect 214010 160440 214066 160449
rect 214010 160375 214066 160384
rect 213920 160064 213972 160070
rect 213920 160006 213972 160012
rect 213932 159769 213960 160006
rect 214012 159996 214064 160002
rect 214012 159938 214064 159944
rect 213918 159760 213974 159769
rect 213918 159695 213974 159704
rect 214024 159089 214052 159938
rect 214010 159080 214066 159089
rect 214010 159015 214066 159024
rect 213920 158704 213972 158710
rect 213920 158646 213972 158652
rect 213932 158409 213960 158646
rect 214012 158636 214064 158642
rect 214012 158578 214064 158584
rect 213918 158400 213974 158409
rect 213918 158335 213974 158344
rect 214024 157729 214052 158578
rect 214010 157720 214066 157729
rect 214010 157655 214066 157664
rect 213920 157344 213972 157350
rect 213920 157286 213972 157292
rect 213932 157185 213960 157286
rect 214012 157276 214064 157282
rect 214012 157218 214064 157224
rect 213918 157176 213974 157185
rect 213918 157111 213974 157120
rect 214024 156505 214052 157218
rect 214010 156496 214066 156505
rect 214010 156431 214066 156440
rect 213920 155916 213972 155922
rect 213920 155858 213972 155864
rect 213932 155825 213960 155858
rect 213918 155816 213974 155825
rect 213918 155751 213974 155760
rect 213918 153776 213974 153785
rect 213918 153711 213974 153720
rect 213932 153270 213960 153711
rect 213920 153264 213972 153270
rect 213920 153206 213972 153212
rect 213918 153096 213974 153105
rect 213918 153031 213974 153040
rect 213932 151842 213960 153031
rect 214010 152552 214066 152561
rect 214010 152487 214066 152496
rect 214024 152114 214052 152487
rect 214012 152108 214064 152114
rect 214012 152050 214064 152056
rect 213920 151836 213972 151842
rect 213920 151778 213972 151784
rect 214010 151192 214066 151201
rect 214010 151127 214066 151136
rect 214024 150550 214052 151127
rect 214012 150544 214064 150550
rect 213918 150512 213974 150521
rect 214012 150486 214064 150492
rect 213918 150447 213920 150456
rect 213972 150447 213974 150456
rect 213920 150418 213972 150424
rect 214012 150408 214064 150414
rect 214012 150350 214064 150356
rect 213920 149728 213972 149734
rect 213920 149670 213972 149676
rect 213932 148481 213960 149670
rect 214024 149161 214052 150350
rect 214576 149841 214604 182174
rect 214668 171057 214696 183534
rect 215220 182918 215248 238575
rect 215300 238060 215352 238066
rect 215300 238002 215352 238008
rect 215312 237250 215340 238002
rect 215300 237244 215352 237250
rect 215300 237186 215352 237192
rect 215390 225040 215446 225049
rect 215390 224975 215446 224984
rect 215404 202881 215432 224975
rect 215680 209774 215708 240244
rect 216048 237386 216076 240244
rect 216036 237380 216088 237386
rect 216036 237322 216088 237328
rect 216048 236162 216076 237322
rect 216600 237289 216628 240244
rect 216586 237280 216642 237289
rect 216586 237215 216642 237224
rect 216036 236156 216088 236162
rect 216036 236098 216088 236104
rect 216600 236065 216628 237215
rect 216034 236056 216090 236065
rect 216034 235991 216090 236000
rect 216586 236056 216642 236065
rect 216586 235991 216642 236000
rect 216048 227497 216076 235991
rect 216034 227488 216090 227497
rect 216034 227423 216090 227432
rect 217152 227118 217180 240244
rect 215944 227112 215996 227118
rect 215944 227054 215996 227060
rect 217140 227112 217192 227118
rect 217140 227054 217192 227060
rect 215956 226409 215984 227054
rect 215942 226400 215998 226409
rect 215942 226335 215998 226344
rect 215956 221542 215984 226335
rect 217520 223582 217548 240244
rect 217508 223576 217560 223582
rect 217508 223518 217560 223524
rect 215944 221536 215996 221542
rect 215944 221478 215996 221484
rect 217520 219434 217548 223518
rect 215496 209746 215708 209774
rect 217336 219406 217548 219434
rect 215496 204270 215524 209746
rect 215484 204264 215536 204270
rect 215484 204206 215536 204212
rect 215496 203658 215524 204206
rect 215484 203652 215536 203658
rect 215484 203594 215536 203600
rect 215390 202872 215446 202881
rect 215390 202807 215446 202816
rect 217336 184210 217364 219406
rect 218072 217326 218100 240244
rect 218440 229094 218468 240244
rect 218440 229066 218744 229094
rect 218060 217320 218112 217326
rect 218060 217262 218112 217268
rect 218072 216730 218100 217262
rect 217980 216702 218100 216730
rect 217414 213888 217470 213897
rect 217414 213823 217470 213832
rect 217428 200122 217456 213823
rect 217416 200116 217468 200122
rect 217416 200058 217468 200064
rect 217980 185706 218008 216702
rect 218716 209681 218744 229066
rect 218992 217326 219020 240244
rect 219544 240145 219572 240244
rect 219530 240136 219586 240145
rect 219530 240071 219586 240080
rect 219438 239456 219494 239465
rect 219438 239391 219494 239400
rect 219452 238746 219480 239391
rect 219530 238912 219586 238921
rect 219530 238847 219586 238856
rect 219440 238740 219492 238746
rect 219440 238682 219492 238688
rect 219544 233170 219572 238847
rect 219912 238754 219940 240244
rect 219912 238726 220308 238754
rect 219912 238678 219940 238726
rect 219900 238672 219952 238678
rect 219900 238614 219952 238620
rect 220174 237416 220230 237425
rect 220174 237351 220230 237360
rect 219532 233164 219584 233170
rect 219532 233106 219584 233112
rect 220084 227792 220136 227798
rect 220084 227734 220136 227740
rect 218980 217320 219032 217326
rect 218980 217262 219032 217268
rect 219440 217320 219492 217326
rect 219440 217262 219492 217268
rect 218702 209672 218758 209681
rect 218702 209607 218758 209616
rect 218716 192681 218744 209607
rect 219452 206922 219480 217262
rect 219440 206916 219492 206922
rect 219440 206858 219492 206864
rect 218702 192672 218758 192681
rect 218702 192607 218758 192616
rect 217968 185700 218020 185706
rect 217968 185642 218020 185648
rect 217324 184204 217376 184210
rect 217324 184146 217376 184152
rect 215208 182912 215260 182918
rect 215208 182854 215260 182860
rect 220096 181558 220124 227734
rect 220188 197305 220216 237351
rect 220280 217326 220308 238726
rect 220464 228954 220492 240244
rect 220452 228948 220504 228954
rect 220452 228890 220504 228896
rect 220464 227798 220492 228890
rect 220452 227792 220504 227798
rect 220452 227734 220504 227740
rect 220268 217320 220320 217326
rect 220268 217262 220320 217268
rect 220728 206916 220780 206922
rect 220728 206858 220780 206864
rect 220740 206310 220768 206858
rect 220728 206304 220780 206310
rect 220728 206246 220780 206252
rect 221016 204241 221044 240244
rect 221384 237425 221412 240244
rect 221370 237416 221426 237425
rect 221370 237351 221426 237360
rect 221936 213897 221964 240244
rect 222304 240009 222332 240244
rect 222290 240000 222346 240009
rect 222290 239935 222346 239944
rect 222304 239737 222332 239935
rect 222290 239728 222346 239737
rect 222290 239663 222346 239672
rect 222856 238746 222884 240244
rect 222844 238740 222896 238746
rect 222844 238682 222896 238688
rect 221922 213888 221978 213897
rect 221922 213823 221978 213832
rect 221002 204232 221058 204241
rect 221002 204167 221058 204176
rect 221462 204232 221518 204241
rect 221462 204167 221518 204176
rect 220174 197296 220230 197305
rect 220174 197231 220230 197240
rect 221372 188420 221424 188426
rect 221372 188362 221424 188368
rect 221384 187066 221412 188362
rect 221372 187060 221424 187066
rect 221372 187002 221424 187008
rect 220084 181552 220136 181558
rect 220084 181494 220136 181500
rect 221476 180169 221504 204167
rect 222108 198824 222160 198830
rect 222108 198766 222160 198772
rect 222120 198694 222148 198766
rect 222108 198688 222160 198694
rect 222108 198630 222160 198636
rect 221554 189136 221610 189145
rect 221554 189071 221610 189080
rect 221462 180160 221518 180169
rect 221462 180095 221518 180104
rect 221568 179353 221596 189071
rect 221554 179344 221610 179353
rect 221554 179279 221610 179288
rect 215298 178120 215354 178129
rect 215298 178055 215354 178064
rect 214930 175944 214986 175953
rect 214930 175879 214986 175888
rect 214654 171048 214710 171057
rect 214654 170983 214710 170992
rect 214944 166433 214972 175879
rect 215312 172446 215340 178055
rect 222856 177993 222884 238682
rect 223028 237448 223080 237454
rect 223028 237390 223080 237396
rect 223040 231810 223068 237390
rect 223028 231804 223080 231810
rect 223028 231746 223080 231752
rect 222934 218240 222990 218249
rect 222934 218175 222990 218184
rect 222948 180266 222976 218175
rect 223040 200870 223068 231746
rect 223408 219337 223436 240244
rect 223776 237454 223804 240244
rect 224328 240106 224356 240244
rect 224316 240100 224368 240106
rect 224316 240042 224368 240048
rect 224328 238134 224356 240042
rect 224316 238128 224368 238134
rect 224316 238070 224368 238076
rect 223764 237448 223816 237454
rect 223764 237390 223816 237396
rect 224222 233880 224278 233889
rect 224222 233815 224278 233824
rect 224236 227798 224264 233815
rect 224224 227792 224276 227798
rect 224224 227734 224276 227740
rect 224880 226001 224908 240244
rect 225248 233238 225276 240244
rect 225236 233232 225288 233238
rect 225236 233174 225288 233180
rect 225604 231872 225656 231878
rect 225604 231814 225656 231820
rect 225616 227050 225644 231814
rect 225604 227044 225656 227050
rect 225604 226986 225656 226992
rect 224866 225992 224922 226001
rect 224866 225927 224922 225936
rect 225800 219434 225828 240244
rect 226168 231878 226196 240244
rect 226720 238377 226748 240244
rect 226892 238808 226944 238814
rect 226892 238750 226944 238756
rect 226706 238368 226762 238377
rect 226706 238303 226762 238312
rect 226156 231872 226208 231878
rect 226156 231814 226208 231820
rect 226720 231198 226748 238303
rect 226904 237153 226932 238750
rect 226890 237144 226946 237153
rect 226890 237079 226946 237088
rect 226984 236088 227036 236094
rect 226984 236030 227036 236036
rect 226708 231192 226760 231198
rect 226708 231134 226760 231140
rect 226340 227112 226392 227118
rect 226340 227054 226392 227060
rect 225616 219406 225828 219434
rect 223394 219328 223450 219337
rect 223394 219263 223450 219272
rect 223408 218249 223436 219263
rect 223394 218240 223450 218249
rect 223394 218175 223450 218184
rect 225616 217977 225644 219406
rect 225602 217968 225658 217977
rect 225602 217903 225658 217912
rect 225616 203590 225644 217903
rect 226352 215257 226380 227054
rect 226996 224641 227024 236030
rect 227272 227798 227300 240244
rect 227260 227792 227312 227798
rect 227260 227734 227312 227740
rect 227640 226273 227668 240244
rect 228192 234569 228220 240244
rect 228744 240038 228772 240244
rect 228732 240032 228784 240038
rect 228732 239974 228784 239980
rect 228362 239728 228418 239737
rect 228362 239663 228418 239672
rect 228178 234560 228234 234569
rect 228178 234495 228234 234504
rect 227718 233880 227774 233889
rect 227718 233815 227774 233824
rect 227732 231713 227760 233815
rect 227718 231704 227774 231713
rect 227718 231639 227774 231648
rect 227812 227792 227864 227798
rect 227812 227734 227864 227740
rect 227626 226264 227682 226273
rect 227626 226199 227682 226208
rect 226982 224632 227038 224641
rect 226982 224567 227038 224576
rect 227718 222864 227774 222873
rect 227718 222799 227774 222808
rect 226338 215248 226394 215257
rect 226338 215183 226394 215192
rect 226352 214849 226380 215183
rect 226338 214840 226394 214849
rect 226338 214775 226394 214784
rect 226982 214840 227038 214849
rect 226982 214775 227038 214784
rect 225604 203584 225656 203590
rect 225604 203526 225656 203532
rect 223028 200864 223080 200870
rect 223028 200806 223080 200812
rect 225696 200252 225748 200258
rect 225696 200194 225748 200200
rect 225708 196353 225736 200194
rect 225694 196344 225750 196353
rect 225694 196279 225750 196288
rect 226340 182844 226392 182850
rect 226340 182786 226392 182792
rect 226352 180713 226380 182786
rect 226996 181665 227024 214775
rect 227076 196716 227128 196722
rect 227076 196658 227128 196664
rect 226982 181656 227038 181665
rect 226982 181591 227038 181600
rect 226892 181484 226944 181490
rect 226892 181426 226944 181432
rect 226338 180704 226394 180713
rect 226338 180639 226394 180648
rect 222936 180260 222988 180266
rect 222936 180202 222988 180208
rect 223396 180192 223448 180198
rect 223396 180134 223448 180140
rect 222842 177984 222898 177993
rect 222842 177919 222898 177928
rect 223408 177313 223436 180134
rect 226340 180124 226392 180130
rect 226340 180066 226392 180072
rect 226352 178673 226380 180066
rect 226338 178664 226394 178673
rect 226338 178599 226394 178608
rect 226338 178528 226394 178537
rect 226338 178463 226394 178472
rect 223486 178256 223542 178265
rect 223486 178191 223542 178200
rect 223500 177954 223528 178191
rect 223488 177948 223540 177954
rect 223488 177890 223540 177896
rect 223394 177304 223450 177313
rect 223394 177239 223450 177248
rect 226352 176050 226380 178463
rect 226904 177410 226932 181426
rect 227088 178770 227116 196658
rect 227076 178764 227128 178770
rect 227076 178706 227128 178712
rect 226892 177404 226944 177410
rect 226892 177346 226944 177352
rect 227732 176225 227760 222799
rect 227824 213926 227852 227734
rect 227812 213920 227864 213926
rect 227812 213862 227864 213868
rect 228376 196722 228404 239663
rect 228744 231130 228772 239974
rect 229112 234569 229140 240244
rect 229664 236094 229692 240244
rect 229652 236088 229704 236094
rect 229652 236030 229704 236036
rect 229098 234560 229154 234569
rect 229098 234495 229154 234504
rect 230216 232937 230244 240244
rect 230584 240145 230612 240244
rect 230570 240136 230626 240145
rect 230570 240071 230626 240080
rect 230584 237862 230612 240071
rect 230572 237856 230624 237862
rect 230572 237798 230624 237804
rect 231136 234734 231164 240244
rect 231124 234728 231176 234734
rect 231124 234670 231176 234676
rect 231122 234016 231178 234025
rect 231122 233951 231178 233960
rect 230202 232928 230258 232937
rect 230202 232863 230258 232872
rect 228732 231124 228784 231130
rect 228732 231066 228784 231072
rect 229744 227724 229796 227730
rect 229744 227666 229796 227672
rect 228548 203652 228600 203658
rect 228548 203594 228600 203600
rect 228364 196716 228416 196722
rect 228364 196658 228416 196664
rect 228364 195356 228416 195362
rect 228364 195298 228416 195304
rect 227812 178016 227864 178022
rect 227812 177958 227864 177964
rect 227824 176769 227852 177958
rect 228376 177154 228404 195298
rect 228456 192568 228508 192574
rect 228456 192510 228508 192516
rect 228468 177342 228496 192510
rect 228560 189854 228588 203594
rect 229100 200864 229152 200870
rect 229100 200806 229152 200812
rect 228638 196344 228694 196353
rect 228638 196279 228694 196288
rect 228652 192574 228680 196279
rect 228640 192568 228692 192574
rect 228640 192510 228692 192516
rect 228548 189848 228600 189854
rect 228548 189790 228600 189796
rect 228456 177336 228508 177342
rect 228456 177278 228508 177284
rect 228376 177126 228496 177154
rect 227810 176760 227866 176769
rect 227810 176695 227866 176704
rect 228364 176588 228416 176594
rect 228364 176530 228416 176536
rect 227718 176216 227774 176225
rect 227718 176151 227774 176160
rect 226340 176044 226392 176050
rect 226340 175986 226392 175992
rect 228376 175953 228404 176530
rect 223670 175944 223726 175953
rect 223670 175879 223726 175888
rect 228362 175944 228418 175953
rect 228468 175930 228496 177126
rect 228546 175944 228602 175953
rect 228468 175902 228546 175930
rect 228362 175879 228418 175888
rect 228546 175879 228602 175888
rect 223684 175846 223712 175879
rect 223672 175840 223724 175846
rect 223672 175782 223724 175788
rect 215300 172440 215352 172446
rect 215300 172382 215352 172388
rect 214930 166424 214986 166433
rect 214930 166359 214986 166368
rect 214838 154456 214894 154465
rect 214838 154391 214894 154400
rect 214562 149832 214618 149841
rect 214562 149767 214618 149776
rect 214010 149152 214066 149161
rect 214010 149087 214066 149096
rect 213918 148472 213974 148481
rect 213918 148407 213974 148416
rect 213918 147928 213974 147937
rect 213918 147863 213974 147872
rect 213932 147694 213960 147863
rect 213920 147688 213972 147694
rect 213920 147630 213972 147636
rect 213918 147248 213974 147257
rect 213918 147183 213974 147192
rect 213932 146334 213960 147183
rect 213920 146328 213972 146334
rect 213920 146270 213972 146276
rect 213918 145888 213974 145897
rect 213918 145823 213974 145832
rect 213932 144974 213960 145823
rect 214470 145208 214526 145217
rect 214470 145143 214526 145152
rect 213920 144968 213972 144974
rect 213920 144910 213972 144916
rect 214010 144528 214066 144537
rect 214010 144463 214066 144472
rect 213918 143848 213974 143857
rect 213918 143783 213974 143792
rect 213932 143682 213960 143783
rect 213920 143676 213972 143682
rect 213920 143618 213972 143624
rect 214024 143614 214052 144463
rect 214012 143608 214064 143614
rect 214012 143550 214064 143556
rect 213918 143304 213974 143313
rect 213918 143239 213974 143248
rect 213932 142186 213960 143239
rect 214010 142624 214066 142633
rect 214010 142559 214066 142568
rect 213920 142180 213972 142186
rect 213920 142122 213972 142128
rect 213274 141944 213330 141953
rect 213274 141879 213330 141888
rect 213288 97306 213316 141879
rect 214024 141438 214052 142559
rect 214012 141432 214064 141438
rect 214012 141374 214064 141380
rect 214010 140584 214066 140593
rect 214010 140519 214066 140528
rect 213918 139904 213974 139913
rect 213918 139839 213974 139848
rect 213932 139466 213960 139839
rect 214024 139534 214052 140519
rect 214012 139528 214064 139534
rect 214012 139470 214064 139476
rect 213920 139460 213972 139466
rect 213920 139402 213972 139408
rect 213918 139224 213974 139233
rect 213918 139159 213974 139168
rect 213932 138038 213960 139159
rect 214484 138718 214512 145143
rect 214852 142154 214880 154391
rect 215942 151872 215998 151881
rect 215942 151807 215998 151816
rect 214668 142126 214880 142154
rect 214472 138712 214524 138718
rect 214472 138654 214524 138660
rect 213920 138032 213972 138038
rect 213920 137974 213972 137980
rect 213918 137320 213974 137329
rect 213918 137255 213974 137264
rect 213932 136678 213960 137255
rect 213920 136672 213972 136678
rect 213920 136614 213972 136620
rect 214010 136640 214066 136649
rect 214010 136575 214066 136584
rect 213918 135960 213974 135969
rect 213918 135895 213974 135904
rect 213932 135318 213960 135895
rect 214024 135386 214052 136575
rect 214012 135380 214064 135386
rect 214012 135322 214064 135328
rect 213920 135312 213972 135318
rect 213920 135254 213972 135260
rect 213920 133952 213972 133958
rect 213918 133920 213920 133929
rect 213972 133920 213974 133929
rect 213918 133855 213974 133864
rect 213918 132696 213974 132705
rect 213918 132631 213974 132640
rect 213932 132530 213960 132631
rect 213920 132524 213972 132530
rect 213920 132466 213972 132472
rect 213918 132016 213974 132025
rect 213918 131951 213974 131960
rect 213932 131170 213960 131951
rect 214668 131782 214696 142126
rect 214746 138000 214802 138009
rect 214746 137935 214802 137944
rect 214760 132494 214788 137935
rect 215956 137290 215984 151807
rect 229112 146849 229140 200806
rect 229192 185700 229244 185706
rect 229192 185642 229244 185648
rect 229204 176905 229232 185642
rect 229756 182170 229784 227666
rect 231136 225622 231164 233951
rect 231504 231849 231532 240244
rect 232056 238754 232084 240244
rect 231964 238726 232084 238754
rect 231768 237856 231820 237862
rect 231768 237798 231820 237804
rect 231490 231840 231546 231849
rect 231490 231775 231546 231784
rect 230388 225616 230440 225622
rect 230388 225558 230440 225564
rect 231124 225616 231176 225622
rect 231124 225558 231176 225564
rect 230400 185910 230428 225558
rect 230572 214668 230624 214674
rect 230572 214610 230624 214616
rect 230480 207732 230532 207738
rect 230480 207674 230532 207680
rect 230388 185904 230440 185910
rect 230388 185846 230440 185852
rect 229744 182164 229796 182170
rect 229744 182106 229796 182112
rect 229282 181384 229338 181393
rect 229282 181319 229338 181328
rect 229296 179994 229324 181319
rect 229284 179988 229336 179994
rect 229284 179930 229336 179936
rect 229374 177984 229430 177993
rect 229374 177919 229430 177928
rect 229190 176896 229246 176905
rect 229190 176831 229246 176840
rect 229190 176624 229246 176633
rect 229190 176559 229246 176568
rect 229204 173369 229232 176559
rect 229282 174584 229338 174593
rect 229282 174519 229284 174528
rect 229336 174519 229338 174528
rect 229284 174490 229336 174496
rect 229190 173360 229246 173369
rect 229190 173295 229246 173304
rect 229388 150657 229416 177919
rect 229744 174820 229796 174826
rect 229744 174762 229796 174768
rect 229756 158137 229784 174762
rect 230018 164928 230074 164937
rect 230018 164863 230074 164872
rect 229742 158128 229798 158137
rect 229742 158063 229798 158072
rect 229742 153776 229798 153785
rect 229742 153711 229798 153720
rect 229374 150648 229430 150657
rect 229374 150583 229430 150592
rect 229098 146840 229154 146849
rect 229098 146775 229154 146784
rect 216034 146568 216090 146577
rect 216034 146503 216090 146512
rect 215944 137284 215996 137290
rect 215944 137226 215996 137232
rect 214760 132466 214880 132494
rect 214656 131776 214708 131782
rect 214656 131718 214708 131724
rect 214562 131336 214618 131345
rect 214562 131271 214618 131280
rect 213920 131164 213972 131170
rect 213920 131106 213972 131112
rect 214010 130656 214066 130665
rect 214010 130591 214066 130600
rect 213918 129976 213974 129985
rect 213918 129911 213974 129920
rect 213932 129810 213960 129911
rect 214024 129878 214052 130591
rect 214012 129872 214064 129878
rect 214012 129814 214064 129820
rect 213920 129804 213972 129810
rect 213920 129746 213972 129752
rect 214010 129296 214066 129305
rect 214010 129231 214066 129240
rect 213918 128752 213974 128761
rect 213918 128687 213974 128696
rect 213932 128382 213960 128687
rect 214024 128450 214052 129231
rect 214012 128444 214064 128450
rect 214012 128386 214064 128392
rect 213920 128376 213972 128382
rect 213920 128318 213972 128324
rect 214010 128072 214066 128081
rect 214010 128007 214066 128016
rect 213918 127392 213974 127401
rect 213918 127327 213974 127336
rect 213932 127090 213960 127327
rect 213920 127084 213972 127090
rect 213920 127026 213972 127032
rect 214024 127022 214052 128007
rect 214012 127016 214064 127022
rect 214012 126958 214064 126964
rect 214010 126712 214066 126721
rect 214010 126647 214066 126656
rect 213918 126032 213974 126041
rect 213918 125967 213974 125976
rect 213932 125662 213960 125967
rect 214024 125730 214052 126647
rect 214012 125724 214064 125730
rect 214012 125666 214064 125672
rect 213920 125656 213972 125662
rect 213920 125598 213972 125604
rect 213918 125352 213974 125361
rect 213918 125287 213974 125296
rect 213932 124234 213960 125287
rect 213920 124228 213972 124234
rect 213920 124170 213972 124176
rect 213918 124128 213974 124137
rect 213918 124063 213974 124072
rect 213366 123448 213422 123457
rect 213366 123383 213422 123392
rect 213276 97300 213328 97306
rect 213276 97242 213328 97248
rect 213380 95198 213408 123383
rect 213932 122874 213960 124063
rect 214010 123448 214066 123457
rect 214010 123383 214066 123392
rect 214024 123146 214052 123383
rect 214012 123140 214064 123146
rect 214012 123082 214064 123088
rect 213920 122868 213972 122874
rect 213920 122810 213972 122816
rect 214010 122768 214066 122777
rect 214010 122703 214066 122712
rect 213918 122088 213974 122097
rect 213918 122023 213974 122032
rect 213932 121514 213960 122023
rect 214024 121582 214052 122703
rect 214012 121576 214064 121582
rect 214012 121518 214064 121524
rect 213920 121508 213972 121514
rect 213920 121450 213972 121456
rect 213918 121408 213974 121417
rect 213918 121343 213974 121352
rect 213932 120154 213960 121343
rect 213920 120148 213972 120154
rect 213920 120090 213972 120096
rect 214010 120048 214066 120057
rect 214010 119983 214066 119992
rect 213918 119504 213974 119513
rect 213918 119439 213974 119448
rect 213932 118794 213960 119439
rect 213920 118788 213972 118794
rect 213920 118730 213972 118736
rect 214024 118726 214052 119983
rect 214012 118720 214064 118726
rect 214012 118662 214064 118668
rect 214010 118144 214066 118153
rect 214010 118079 214066 118088
rect 213918 117464 213974 117473
rect 213918 117399 213920 117408
rect 213972 117399 213974 117408
rect 213920 117370 213972 117376
rect 214024 117366 214052 118079
rect 214012 117360 214064 117366
rect 214012 117302 214064 117308
rect 214010 116784 214066 116793
rect 214010 116719 214066 116728
rect 213918 116104 213974 116113
rect 214024 116074 214052 116719
rect 213918 116039 213974 116048
rect 214012 116068 214064 116074
rect 213932 116006 213960 116039
rect 214012 116010 214064 116016
rect 213920 116000 213972 116006
rect 213920 115942 213972 115948
rect 213918 114880 213974 114889
rect 213918 114815 213974 114824
rect 213932 114578 213960 114815
rect 213920 114572 213972 114578
rect 213920 114514 213972 114520
rect 214010 114200 214066 114209
rect 214010 114135 214066 114144
rect 213918 113520 213974 113529
rect 213918 113455 213974 113464
rect 213932 113218 213960 113455
rect 214024 113286 214052 114135
rect 214012 113280 214064 113286
rect 214012 113222 214064 113228
rect 213920 113212 213972 113218
rect 213920 113154 213972 113160
rect 213918 112160 213974 112169
rect 213918 112095 213974 112104
rect 213932 111858 213960 112095
rect 213920 111852 213972 111858
rect 213920 111794 213972 111800
rect 214010 111480 214066 111489
rect 214010 111415 214066 111424
rect 213918 110800 213974 110809
rect 213918 110735 213974 110744
rect 213932 110566 213960 110735
rect 213920 110560 213972 110566
rect 213920 110502 213972 110508
rect 214024 110498 214052 111415
rect 214012 110492 214064 110498
rect 214012 110434 214064 110440
rect 213918 110256 213974 110265
rect 213918 110191 213974 110200
rect 213932 109070 213960 110191
rect 213920 109064 213972 109070
rect 213920 109006 213972 109012
rect 214010 108896 214066 108905
rect 214010 108831 214066 108840
rect 213918 108216 213974 108225
rect 213918 108151 213974 108160
rect 213932 107710 213960 108151
rect 214024 107778 214052 108831
rect 214576 108361 214604 131271
rect 214852 120766 214880 132466
rect 214930 124672 214986 124681
rect 214930 124607 214986 124616
rect 214840 120760 214892 120766
rect 214840 120702 214892 120708
rect 214838 115424 214894 115433
rect 214838 115359 214894 115368
rect 214746 112840 214802 112849
rect 214746 112775 214802 112784
rect 214562 108352 214618 108361
rect 214562 108287 214618 108296
rect 214012 107772 214064 107778
rect 214012 107714 214064 107720
rect 213920 107704 213972 107710
rect 213920 107646 213972 107652
rect 214010 107536 214066 107545
rect 214010 107471 214066 107480
rect 213918 106856 213974 106865
rect 213918 106791 213974 106800
rect 213932 106418 213960 106791
rect 213920 106412 213972 106418
rect 213920 106354 213972 106360
rect 214024 106350 214052 107471
rect 214012 106344 214064 106350
rect 214012 106286 214064 106292
rect 214010 106176 214066 106185
rect 214010 106111 214066 106120
rect 213920 104984 213972 104990
rect 213918 104952 213920 104961
rect 213972 104952 213974 104961
rect 214024 104922 214052 106111
rect 214378 105632 214434 105641
rect 214378 105567 214434 105576
rect 213918 104887 213974 104896
rect 214012 104916 214064 104922
rect 214012 104858 214064 104864
rect 213918 103592 213974 103601
rect 213918 103527 213920 103536
rect 213972 103527 213974 103536
rect 213920 103498 213972 103504
rect 214010 102912 214066 102921
rect 214010 102847 214066 102856
rect 213920 102264 213972 102270
rect 213918 102232 213920 102241
rect 213972 102232 213974 102241
rect 214024 102202 214052 102847
rect 213918 102167 213974 102176
rect 214012 102196 214064 102202
rect 214012 102138 214064 102144
rect 213918 101552 213974 101561
rect 213918 101487 213974 101496
rect 213932 100774 213960 101487
rect 214392 101425 214420 105567
rect 214378 101416 214434 101425
rect 214378 101351 214434 101360
rect 213920 100768 213972 100774
rect 213920 100710 213972 100716
rect 214010 100328 214066 100337
rect 214010 100263 214066 100272
rect 213918 99648 213974 99657
rect 213918 99583 213974 99592
rect 213932 99414 213960 99583
rect 214024 99482 214052 100263
rect 214012 99476 214064 99482
rect 214012 99418 214064 99424
rect 213920 99408 213972 99414
rect 213920 99350 213972 99356
rect 214010 98968 214066 98977
rect 214010 98903 214066 98912
rect 213918 98288 213974 98297
rect 213918 98223 213974 98232
rect 213932 98054 213960 98223
rect 214024 98122 214052 98903
rect 214760 98682 214788 112775
rect 214852 112470 214880 115359
rect 214944 115258 214972 124607
rect 214932 115252 214984 115258
rect 214932 115194 214984 115200
rect 214840 112464 214892 112470
rect 214840 112406 214892 112412
rect 214838 101008 214894 101017
rect 214838 100943 214894 100952
rect 214576 98654 214788 98682
rect 214012 98116 214064 98122
rect 214012 98058 214064 98064
rect 213920 98048 213972 98054
rect 213920 97990 213972 97996
rect 213458 97608 213514 97617
rect 213458 97543 213514 97552
rect 213368 95192 213420 95198
rect 213368 95134 213420 95140
rect 213276 89004 213328 89010
rect 213276 88946 213328 88952
rect 213288 42158 213316 88946
rect 213472 85513 213500 97543
rect 213918 96384 213974 96393
rect 213918 96319 213974 96328
rect 213932 95266 213960 96319
rect 213920 95260 213972 95266
rect 213920 95202 213972 95208
rect 214576 93226 214604 98654
rect 214852 97458 214880 100943
rect 214668 97430 214880 97458
rect 214564 93220 214616 93226
rect 214564 93162 214616 93168
rect 214564 91792 214616 91798
rect 214564 91734 214616 91740
rect 213458 85504 213514 85513
rect 213458 85439 213514 85448
rect 213276 42152 213328 42158
rect 213276 42094 213328 42100
rect 214576 3466 214604 91734
rect 214668 53786 214696 97430
rect 214838 96928 214894 96937
rect 214838 96863 214894 96872
rect 214748 87644 214800 87650
rect 214748 87586 214800 87592
rect 214760 67153 214788 87586
rect 214852 86873 214880 96863
rect 214838 86864 214894 86873
rect 214838 86799 214894 86808
rect 215944 84924 215996 84930
rect 215944 84866 215996 84872
rect 214746 67144 214802 67153
rect 214746 67079 214802 67088
rect 214656 53780 214708 53786
rect 214656 53722 214708 53728
rect 215956 11762 215984 84866
rect 216048 80034 216076 146503
rect 229756 141137 229784 153711
rect 229926 148336 229982 148345
rect 229926 148271 229982 148280
rect 229742 141128 229798 141137
rect 229742 141063 229798 141072
rect 229742 137184 229798 137193
rect 229742 137119 229798 137128
rect 216126 120728 216182 120737
rect 216126 120663 216182 120672
rect 216036 80028 216088 80034
rect 216036 79970 216088 79976
rect 216140 56574 216168 120663
rect 217230 118416 217286 118425
rect 217230 118351 217286 118360
rect 216128 56568 216180 56574
rect 216128 56510 216180 56516
rect 217244 43518 217272 118351
rect 229098 97880 229154 97889
rect 229020 97838 229098 97866
rect 229020 96694 229048 97838
rect 229098 97815 229154 97824
rect 229008 96688 229060 96694
rect 229008 96630 229060 96636
rect 223672 96076 223724 96082
rect 223672 96018 223724 96024
rect 223684 95985 223712 96018
rect 223670 95976 223726 95985
rect 223670 95911 223726 95920
rect 225604 95328 225656 95334
rect 225604 95270 225656 95276
rect 229098 95296 229154 95305
rect 222936 94512 222988 94518
rect 222936 94454 222988 94460
rect 222844 92540 222896 92546
rect 222844 92482 222896 92488
rect 218704 90432 218756 90438
rect 218704 90374 218756 90380
rect 217232 43512 217284 43518
rect 217232 43454 217284 43460
rect 218716 31142 218744 90374
rect 221464 89072 221516 89078
rect 221464 89014 221516 89020
rect 220084 86352 220136 86358
rect 220084 86294 220136 86300
rect 218704 31136 218756 31142
rect 218704 31078 218756 31084
rect 215944 11756 215996 11762
rect 215944 11698 215996 11704
rect 220096 10402 220124 86294
rect 221476 26926 221504 89014
rect 221464 26920 221516 26926
rect 221464 26862 221516 26868
rect 220084 10396 220136 10402
rect 220084 10338 220136 10344
rect 214564 3460 214616 3466
rect 214564 3402 214616 3408
rect 200762 3360 200818 3369
rect 200762 3295 200818 3304
rect 213182 3360 213238 3369
rect 213182 3295 213238 3304
rect 198096 2168 198148 2174
rect 198096 2110 198148 2116
rect 222856 2106 222884 92482
rect 222948 18698 222976 94454
rect 224222 89176 224278 89185
rect 224222 89111 224278 89120
rect 222936 18692 222988 18698
rect 222936 18634 222988 18640
rect 224236 7614 224264 89111
rect 225616 64297 225644 95270
rect 227076 95260 227128 95266
rect 229098 95231 229100 95240
rect 227076 95202 227128 95208
rect 229152 95231 229154 95240
rect 229100 95202 229152 95208
rect 226984 84856 227036 84862
rect 226984 84798 227036 84804
rect 225602 64288 225658 64297
rect 225602 64223 225658 64232
rect 226996 14482 227024 84798
rect 227088 43489 227116 95202
rect 228362 93120 228418 93129
rect 228362 93055 228418 93064
rect 227074 43480 227130 43489
rect 227074 43415 227130 43424
rect 226984 14476 227036 14482
rect 226984 14418 227036 14424
rect 224224 7608 224276 7614
rect 224224 7550 224276 7556
rect 228376 6186 228404 93055
rect 228456 64184 228508 64190
rect 228456 64126 228508 64132
rect 228364 6180 228416 6186
rect 228364 6122 228416 6128
rect 228468 4826 228496 64126
rect 229756 60110 229784 137119
rect 229834 132016 229890 132025
rect 229834 131951 229890 131960
rect 229848 87718 229876 131951
rect 229940 105641 229968 148271
rect 230032 137329 230060 164863
rect 230492 152402 230520 207674
rect 230584 166326 230612 214610
rect 230756 182164 230808 182170
rect 230756 182106 230808 182112
rect 230768 173777 230796 182106
rect 231780 182073 231808 237798
rect 231964 229770 231992 238726
rect 232608 235657 232636 240244
rect 232594 235648 232650 235657
rect 232594 235583 232650 235592
rect 232044 234728 232096 234734
rect 232044 234670 232096 234676
rect 231952 229764 232004 229770
rect 231952 229706 232004 229712
rect 232056 219434 232084 234670
rect 232976 228857 233004 240244
rect 233528 228993 233556 240244
rect 234080 237561 234108 240244
rect 234066 237552 234122 237561
rect 234066 237487 234122 237496
rect 234080 230382 234108 237487
rect 234068 230376 234120 230382
rect 234068 230318 234120 230324
rect 233514 228984 233570 228993
rect 233514 228919 233570 228928
rect 232962 228848 233018 228857
rect 232962 228783 233018 228792
rect 233882 228304 233938 228313
rect 233882 228239 233938 228248
rect 231872 219406 232084 219434
rect 231872 217394 231900 219406
rect 231860 217388 231912 217394
rect 231860 217330 231912 217336
rect 231872 216753 231900 217330
rect 231858 216744 231914 216753
rect 231858 216679 231914 216688
rect 233516 212492 233568 212498
rect 233516 212434 233568 212440
rect 233330 205728 233386 205737
rect 233330 205663 233386 205672
rect 232042 196752 232098 196761
rect 232042 196687 232098 196696
rect 231952 189780 232004 189786
rect 231952 189722 232004 189728
rect 231860 185904 231912 185910
rect 231860 185846 231912 185852
rect 231766 182064 231822 182073
rect 231766 181999 231822 182008
rect 231766 178256 231822 178265
rect 231766 178191 231822 178200
rect 231490 176624 231546 176633
rect 231490 176559 231546 176568
rect 230940 175160 230992 175166
rect 230940 175102 230992 175108
rect 230846 173904 230902 173913
rect 230846 173839 230902 173848
rect 230754 173768 230810 173777
rect 230754 173703 230810 173712
rect 230664 170808 230716 170814
rect 230664 170750 230716 170756
rect 230676 170513 230704 170750
rect 230662 170504 230718 170513
rect 230662 170439 230718 170448
rect 230572 166320 230624 166326
rect 230572 166262 230624 166268
rect 230860 161474 230888 173839
rect 230952 169561 230980 175102
rect 231504 174729 231532 176559
rect 231780 175982 231808 178191
rect 231768 175976 231820 175982
rect 231768 175918 231820 175924
rect 231766 175264 231822 175273
rect 231766 175199 231768 175208
rect 231820 175199 231822 175208
rect 231768 175170 231820 175176
rect 231490 174720 231546 174729
rect 231490 174655 231546 174664
rect 231584 173868 231636 173874
rect 231584 173810 231636 173816
rect 231596 172825 231624 173810
rect 231582 172816 231638 172825
rect 231582 172751 231638 172760
rect 231124 172236 231176 172242
rect 231124 172178 231176 172184
rect 231136 171465 231164 172178
rect 231768 171896 231820 171902
rect 231766 171864 231768 171873
rect 231820 171864 231822 171873
rect 231766 171799 231822 171808
rect 231122 171456 231178 171465
rect 231122 171391 231178 171400
rect 231216 170060 231268 170066
rect 231216 170002 231268 170008
rect 231228 169969 231256 170002
rect 231214 169960 231270 169969
rect 231214 169895 231270 169904
rect 230938 169552 230994 169561
rect 230938 169487 230994 169496
rect 231676 169448 231728 169454
rect 231676 169390 231728 169396
rect 231688 169017 231716 169390
rect 231674 169008 231730 169017
rect 231674 168943 231730 168952
rect 230940 168292 230992 168298
rect 230940 168234 230992 168240
rect 230952 167657 230980 168234
rect 230938 167648 230994 167657
rect 230938 167583 230994 167592
rect 231676 167476 231728 167482
rect 231676 167418 231728 167424
rect 231688 167113 231716 167418
rect 231674 167104 231730 167113
rect 231674 167039 231730 167048
rect 231308 167000 231360 167006
rect 231308 166942 231360 166948
rect 230940 166320 230992 166326
rect 230940 166262 230992 166268
rect 230676 161446 230888 161474
rect 230676 152561 230704 161446
rect 230952 158681 230980 166262
rect 231320 166161 231348 166942
rect 231676 166320 231728 166326
rect 231676 166262 231728 166268
rect 231306 166152 231362 166161
rect 231306 166087 231362 166096
rect 231688 165753 231716 166262
rect 231674 165744 231730 165753
rect 231674 165679 231730 165688
rect 231124 165572 231176 165578
rect 231124 165514 231176 165520
rect 231136 164393 231164 165514
rect 231122 164384 231178 164393
rect 231122 164319 231178 164328
rect 231584 164212 231636 164218
rect 231584 164154 231636 164160
rect 231492 164008 231544 164014
rect 231492 163950 231544 163956
rect 231504 163849 231532 163950
rect 231490 163840 231546 163849
rect 231490 163775 231546 163784
rect 231596 162897 231624 164154
rect 231582 162888 231638 162897
rect 231582 162823 231638 162832
rect 231768 162852 231820 162858
rect 231768 162794 231820 162800
rect 231780 161945 231808 162794
rect 231766 161936 231822 161945
rect 231766 161871 231822 161880
rect 231768 161424 231820 161430
rect 231768 161366 231820 161372
rect 231308 161016 231360 161022
rect 231780 160993 231808 161366
rect 231308 160958 231360 160964
rect 231766 160984 231822 160993
rect 231320 160585 231348 160958
rect 231766 160919 231822 160928
rect 231582 160712 231638 160721
rect 231582 160647 231638 160656
rect 231306 160576 231362 160585
rect 231306 160511 231362 160520
rect 231596 159089 231624 160647
rect 231768 160064 231820 160070
rect 231766 160032 231768 160041
rect 231820 160032 231822 160041
rect 231676 159996 231728 160002
rect 231766 159967 231822 159976
rect 231676 159938 231728 159944
rect 231688 159633 231716 159938
rect 231674 159624 231730 159633
rect 231674 159559 231730 159568
rect 231582 159080 231638 159089
rect 231582 159015 231638 159024
rect 230938 158672 230994 158681
rect 230938 158607 230994 158616
rect 231492 158160 231544 158166
rect 231492 158102 231544 158108
rect 231504 157729 231532 158102
rect 231490 157720 231546 157729
rect 231490 157655 231546 157664
rect 231122 157448 231178 157457
rect 231122 157383 231178 157392
rect 230756 155848 230808 155854
rect 230756 155790 230808 155796
rect 230768 155281 230796 155790
rect 230754 155272 230810 155281
rect 230754 155207 230810 155216
rect 230662 152552 230718 152561
rect 230662 152487 230718 152496
rect 230492 152374 230888 152402
rect 230756 151836 230808 151842
rect 230756 151778 230808 151784
rect 230768 148753 230796 151778
rect 230754 148744 230810 148753
rect 230754 148679 230810 148688
rect 230860 147801 230888 152374
rect 231136 151609 231164 157383
rect 231768 157344 231820 157350
rect 231768 157286 231820 157292
rect 231780 156777 231808 157286
rect 231766 156768 231822 156777
rect 231766 156703 231822 156712
rect 231492 156664 231544 156670
rect 231492 156606 231544 156612
rect 231504 155825 231532 156606
rect 231490 155816 231546 155825
rect 231490 155751 231546 155760
rect 231768 155440 231820 155446
rect 231768 155382 231820 155388
rect 231584 154556 231636 154562
rect 231584 154498 231636 154504
rect 231596 153377 231624 154498
rect 231676 154352 231728 154358
rect 231674 154320 231676 154329
rect 231728 154320 231730 154329
rect 231674 154255 231730 154264
rect 231780 153921 231808 155382
rect 231766 153912 231822 153921
rect 231766 153847 231822 153856
rect 231582 153368 231638 153377
rect 231582 153303 231638 153312
rect 231766 153096 231822 153105
rect 231766 153031 231822 153040
rect 231780 152017 231808 153031
rect 231872 152969 231900 185846
rect 231964 164801 231992 189722
rect 232056 174826 232084 196687
rect 232136 187060 232188 187066
rect 232136 187002 232188 187008
rect 232044 174820 232096 174826
rect 232044 174762 232096 174768
rect 232042 174584 232098 174593
rect 232042 174519 232098 174528
rect 231950 164792 232006 164801
rect 231950 164727 232006 164736
rect 232056 163441 232084 174519
rect 232148 170814 232176 187002
rect 233240 177336 233292 177342
rect 233240 177278 233292 177284
rect 232136 170808 232188 170814
rect 232136 170750 232188 170756
rect 233252 170066 233280 177278
rect 233344 172242 233372 205663
rect 233422 183016 233478 183025
rect 233422 182951 233478 182960
rect 233332 172236 233384 172242
rect 233332 172178 233384 172184
rect 233240 170060 233292 170066
rect 233240 170002 233292 170008
rect 232136 169788 232188 169794
rect 232136 169730 232188 169736
rect 232148 166326 232176 169730
rect 233436 168298 233464 182951
rect 233424 168292 233476 168298
rect 233424 168234 233476 168240
rect 232136 166320 232188 166326
rect 232136 166262 232188 166268
rect 232780 165640 232832 165646
rect 232502 165608 232558 165617
rect 232780 165582 232832 165588
rect 232502 165543 232558 165552
rect 232042 163432 232098 163441
rect 232042 163367 232098 163376
rect 232516 155854 232544 165543
rect 232596 162172 232648 162178
rect 232596 162114 232648 162120
rect 232504 155848 232556 155854
rect 232504 155790 232556 155796
rect 231858 152960 231914 152969
rect 231858 152895 231914 152904
rect 231766 152008 231822 152017
rect 231766 151943 231822 151952
rect 231768 151768 231820 151774
rect 231768 151710 231820 151716
rect 231122 151600 231178 151609
rect 231122 151535 231178 151544
rect 231780 151065 231808 151710
rect 231766 151056 231822 151065
rect 231766 150991 231822 151000
rect 231674 150920 231730 150929
rect 231674 150855 231730 150864
rect 231492 150340 231544 150346
rect 231492 150282 231544 150288
rect 231504 149161 231532 150282
rect 231490 149152 231546 149161
rect 231490 149087 231546 149096
rect 231308 148368 231360 148374
rect 231308 148310 231360 148316
rect 230846 147792 230902 147801
rect 230846 147727 230902 147736
rect 231124 147008 231176 147014
rect 231124 146950 231176 146956
rect 230756 146192 230808 146198
rect 230756 146134 230808 146140
rect 230768 145897 230796 146134
rect 230754 145888 230810 145897
rect 230754 145823 230810 145832
rect 230754 144664 230810 144673
rect 230754 144599 230810 144608
rect 230296 144220 230348 144226
rect 230296 144162 230348 144168
rect 230308 143449 230336 144162
rect 230768 143993 230796 144599
rect 230754 143984 230810 143993
rect 230754 143919 230810 143928
rect 230294 143440 230350 143449
rect 230294 143375 230350 143384
rect 230664 142860 230716 142866
rect 230664 142802 230716 142808
rect 230676 140729 230704 142802
rect 230940 141432 230992 141438
rect 230940 141374 230992 141380
rect 230662 140720 230718 140729
rect 230662 140655 230718 140664
rect 230018 137320 230074 137329
rect 230018 137255 230074 137264
rect 230952 135425 230980 141374
rect 230938 135416 230994 135425
rect 230938 135351 230994 135360
rect 230572 133612 230624 133618
rect 230572 133554 230624 133560
rect 230584 129849 230612 133554
rect 231136 131209 231164 146950
rect 231320 144401 231348 148310
rect 231688 147257 231716 150855
rect 231768 150408 231820 150414
rect 231768 150350 231820 150356
rect 231780 150113 231808 150350
rect 231766 150104 231822 150113
rect 231766 150039 231822 150048
rect 231768 149048 231820 149054
rect 231768 148990 231820 148996
rect 231780 148209 231808 148990
rect 231766 148200 231822 148209
rect 231766 148135 231822 148144
rect 231674 147248 231730 147257
rect 231674 147183 231730 147192
rect 231398 146976 231454 146985
rect 231398 146911 231454 146920
rect 231306 144392 231362 144401
rect 231306 144327 231362 144336
rect 231412 142154 231440 146911
rect 231766 146296 231822 146305
rect 231766 146231 231822 146240
rect 231780 144809 231808 146231
rect 232608 146198 232636 162114
rect 232686 155000 232742 155009
rect 232686 154935 232742 154944
rect 232596 146192 232648 146198
rect 232596 146134 232648 146140
rect 232504 144968 232556 144974
rect 232504 144910 232556 144916
rect 231766 144800 231822 144809
rect 231766 144735 231822 144744
rect 231768 143540 231820 143546
rect 231768 143482 231820 143488
rect 231780 143041 231808 143482
rect 231766 143032 231822 143041
rect 231766 142967 231822 142976
rect 231320 142126 231440 142154
rect 231320 141681 231348 142126
rect 231306 141672 231362 141681
rect 231306 141607 231362 141616
rect 231216 141500 231268 141506
rect 231216 141442 231268 141448
rect 231122 131200 231178 131209
rect 230940 131164 230992 131170
rect 231122 131135 231178 131144
rect 230940 131106 230992 131112
rect 230570 129840 230626 129849
rect 230570 129775 230626 129784
rect 230756 129600 230808 129606
rect 230756 129542 230808 129548
rect 230768 128897 230796 129542
rect 230754 128888 230810 128897
rect 230754 128823 230810 128832
rect 230952 126449 230980 131106
rect 231228 130665 231256 141442
rect 231308 140752 231360 140758
rect 231308 140694 231360 140700
rect 231320 139777 231348 140694
rect 231306 139768 231362 139777
rect 231306 139703 231362 139712
rect 231768 139392 231820 139398
rect 231768 139334 231820 139340
rect 231780 138281 231808 139334
rect 231766 138272 231822 138281
rect 231766 138207 231822 138216
rect 231584 137964 231636 137970
rect 231584 137906 231636 137912
rect 231596 136921 231624 137906
rect 231676 137624 231728 137630
rect 231676 137566 231728 137572
rect 231582 136912 231638 136921
rect 231582 136847 231638 136856
rect 231400 136604 231452 136610
rect 231400 136546 231452 136552
rect 231308 135992 231360 135998
rect 231412 135969 231440 136546
rect 231308 135934 231360 135940
rect 231398 135960 231454 135969
rect 231214 130656 231270 130665
rect 231214 130591 231270 130600
rect 231320 129146 231348 135934
rect 231398 135895 231454 135904
rect 231492 135176 231544 135182
rect 231492 135118 231544 135124
rect 231504 134065 231532 135118
rect 231688 134473 231716 137566
rect 231768 135244 231820 135250
rect 231768 135186 231820 135192
rect 231780 135017 231808 135186
rect 231766 135008 231822 135017
rect 231766 134943 231822 134952
rect 231674 134464 231730 134473
rect 231674 134399 231730 134408
rect 231490 134056 231546 134065
rect 231490 133991 231546 134000
rect 231676 133272 231728 133278
rect 231676 133214 231728 133220
rect 231688 132569 231716 133214
rect 231674 132560 231730 132569
rect 231674 132495 231730 132504
rect 231768 132456 231820 132462
rect 231768 132398 231820 132404
rect 231780 132161 231808 132398
rect 231766 132152 231822 132161
rect 231766 132087 231822 132096
rect 231768 131096 231820 131102
rect 231768 131038 231820 131044
rect 231780 130257 231808 131038
rect 231766 130248 231822 130257
rect 231766 130183 231822 130192
rect 231768 129736 231820 129742
rect 231768 129678 231820 129684
rect 231780 129305 231808 129678
rect 231766 129296 231822 129305
rect 231766 129231 231822 129240
rect 231228 129118 231348 129146
rect 231124 127764 231176 127770
rect 231124 127706 231176 127712
rect 231136 127401 231164 127706
rect 231122 127392 231178 127401
rect 231122 127327 231178 127336
rect 230938 126440 230994 126449
rect 230938 126375 230994 126384
rect 231228 126041 231256 129118
rect 231306 129024 231362 129033
rect 231306 128959 231362 128968
rect 231214 126032 231270 126041
rect 231214 125967 231270 125976
rect 230480 125588 230532 125594
rect 230480 125530 230532 125536
rect 230492 124545 230520 125530
rect 231320 125497 231348 128959
rect 231768 128308 231820 128314
rect 231768 128250 231820 128256
rect 231780 127945 231808 128250
rect 231766 127936 231822 127945
rect 231766 127871 231822 127880
rect 231766 126984 231822 126993
rect 231766 126919 231768 126928
rect 231820 126919 231822 126928
rect 231768 126890 231820 126896
rect 231400 126268 231452 126274
rect 231400 126210 231452 126216
rect 231306 125488 231362 125497
rect 231306 125423 231362 125432
rect 230664 124908 230716 124914
rect 230664 124850 230716 124856
rect 230478 124536 230534 124545
rect 230478 124471 230534 124480
rect 230018 121816 230074 121825
rect 230018 121751 230074 121760
rect 229926 105632 229982 105641
rect 229926 105567 229982 105576
rect 230032 92546 230060 121751
rect 230676 120329 230704 124850
rect 231122 124808 231178 124817
rect 231122 124743 231178 124752
rect 230662 120320 230718 120329
rect 230662 120255 230718 120264
rect 230940 118720 230992 118726
rect 230940 118662 230992 118668
rect 230952 118017 230980 118662
rect 230938 118008 230994 118017
rect 230756 117972 230808 117978
rect 230938 117943 230994 117952
rect 230756 117914 230808 117920
rect 230768 116113 230796 117914
rect 230754 116104 230810 116113
rect 230754 116039 230810 116048
rect 230940 115864 230992 115870
rect 230940 115806 230992 115812
rect 230952 114617 230980 115806
rect 230938 114608 230994 114617
rect 230938 114543 230994 114552
rect 230572 114164 230624 114170
rect 230572 114106 230624 114112
rect 230584 113665 230612 114106
rect 230570 113656 230626 113665
rect 230570 113591 230626 113600
rect 230756 105596 230808 105602
rect 230756 105538 230808 105544
rect 230572 102876 230624 102882
rect 230572 102818 230624 102824
rect 230584 102785 230612 102818
rect 230570 102776 230626 102785
rect 230570 102711 230626 102720
rect 230768 96665 230796 105538
rect 231136 104689 231164 124743
rect 231412 124522 231440 126210
rect 231228 124494 231440 124522
rect 231228 120737 231256 124494
rect 231768 124160 231820 124166
rect 231766 124128 231768 124137
rect 231820 124128 231822 124137
rect 231400 124092 231452 124098
rect 231766 124063 231822 124072
rect 231400 124034 231452 124040
rect 231412 123185 231440 124034
rect 231398 123176 231454 123185
rect 231398 123111 231454 123120
rect 231768 122800 231820 122806
rect 231768 122742 231820 122748
rect 231492 122732 231544 122738
rect 231492 122674 231544 122680
rect 231504 121689 231532 122674
rect 231780 122233 231808 122742
rect 231766 122224 231822 122233
rect 231766 122159 231822 122168
rect 231490 121680 231546 121689
rect 231490 121615 231546 121624
rect 231768 121440 231820 121446
rect 231768 121382 231820 121388
rect 231780 121281 231808 121382
rect 231766 121272 231822 121281
rect 231766 121207 231822 121216
rect 231214 120728 231270 120737
rect 231214 120663 231270 120672
rect 231400 120148 231452 120154
rect 231400 120090 231452 120096
rect 231308 113076 231360 113082
rect 231308 113018 231360 113024
rect 231320 112305 231348 113018
rect 231306 112296 231362 112305
rect 231306 112231 231362 112240
rect 231412 111353 231440 120090
rect 231492 120080 231544 120086
rect 231492 120022 231544 120028
rect 231766 120048 231822 120057
rect 231504 118969 231532 120022
rect 231766 119983 231822 119992
rect 231780 119377 231808 119983
rect 231766 119368 231822 119377
rect 231766 119303 231822 119312
rect 231490 118960 231546 118969
rect 231490 118895 231546 118904
rect 231584 118652 231636 118658
rect 231584 118594 231636 118600
rect 231596 117473 231624 118594
rect 231674 118008 231730 118017
rect 231674 117943 231730 117952
rect 231582 117464 231638 117473
rect 231582 117399 231638 117408
rect 231492 117224 231544 117230
rect 231492 117166 231544 117172
rect 231504 116521 231532 117166
rect 231490 116512 231546 116521
rect 231490 116447 231546 116456
rect 231492 115932 231544 115938
rect 231492 115874 231544 115880
rect 231504 115161 231532 115874
rect 231490 115152 231546 115161
rect 231490 115087 231546 115096
rect 231688 115002 231716 117943
rect 231768 117292 231820 117298
rect 231768 117234 231820 117240
rect 231780 117065 231808 117234
rect 231766 117056 231822 117065
rect 231766 116991 231822 117000
rect 231504 114974 231716 115002
rect 231398 111344 231454 111353
rect 231398 111279 231454 111288
rect 231306 111072 231362 111081
rect 231306 111007 231362 111016
rect 231216 110356 231268 110362
rect 231216 110298 231268 110304
rect 231228 109857 231256 110298
rect 231214 109848 231270 109857
rect 231214 109783 231270 109792
rect 231216 107636 231268 107642
rect 231216 107578 231268 107584
rect 231228 107137 231256 107578
rect 231214 107128 231270 107137
rect 231214 107063 231270 107072
rect 231320 106978 231348 111007
rect 231400 108996 231452 109002
rect 231400 108938 231452 108944
rect 231412 107953 231440 108938
rect 231398 107944 231454 107953
rect 231398 107879 231454 107888
rect 231228 106950 231348 106978
rect 231122 104680 231178 104689
rect 231122 104615 231178 104624
rect 231228 101833 231256 106950
rect 231308 104848 231360 104854
rect 231308 104790 231360 104796
rect 231320 104281 231348 104790
rect 231306 104272 231362 104281
rect 231306 104207 231362 104216
rect 231308 103964 231360 103970
rect 231308 103906 231360 103912
rect 231320 103737 231348 103906
rect 231306 103728 231362 103737
rect 231306 103663 231362 103672
rect 231504 103329 231532 114974
rect 231676 114504 231728 114510
rect 231676 114446 231728 114452
rect 231688 113257 231716 114446
rect 231674 113248 231730 113257
rect 231674 113183 231730 113192
rect 231768 113144 231820 113150
rect 231768 113086 231820 113092
rect 231780 112713 231808 113086
rect 231766 112704 231822 112713
rect 231766 112639 231822 112648
rect 231768 111784 231820 111790
rect 231674 111752 231730 111761
rect 231768 111726 231820 111732
rect 231674 111687 231676 111696
rect 231728 111687 231730 111696
rect 231676 111658 231728 111664
rect 231780 110809 231808 111726
rect 231766 110800 231822 110809
rect 231766 110735 231822 110744
rect 231768 110424 231820 110430
rect 231768 110366 231820 110372
rect 231780 109449 231808 110366
rect 231766 109440 231822 109449
rect 231766 109375 231822 109384
rect 231768 108928 231820 108934
rect 231768 108870 231820 108876
rect 231780 108497 231808 108870
rect 231766 108488 231822 108497
rect 231766 108423 231822 108432
rect 231768 107568 231820 107574
rect 231768 107510 231820 107516
rect 231780 106593 231808 107510
rect 231766 106584 231822 106593
rect 231766 106519 231822 106528
rect 231768 106276 231820 106282
rect 231768 106218 231820 106224
rect 231780 105233 231808 106218
rect 231766 105224 231822 105233
rect 231766 105159 231822 105168
rect 231584 103420 231636 103426
rect 231584 103362 231636 103368
rect 231490 103320 231546 103329
rect 231490 103255 231546 103264
rect 231306 102912 231362 102921
rect 231306 102847 231362 102856
rect 231214 101824 231270 101833
rect 231214 101759 231270 101768
rect 231216 99272 231268 99278
rect 231216 99214 231268 99220
rect 231228 98977 231256 99214
rect 231214 98968 231270 98977
rect 231214 98903 231270 98912
rect 231122 98832 231178 98841
rect 231122 98767 231178 98776
rect 230754 96656 230810 96665
rect 230754 96591 230810 96600
rect 230478 96248 230534 96257
rect 230478 96183 230534 96192
rect 230492 95538 230520 96183
rect 230480 95532 230532 95538
rect 230480 95474 230532 95480
rect 230020 92540 230072 92546
rect 230020 92482 230072 92488
rect 229836 87712 229888 87718
rect 229836 87654 229888 87660
rect 229744 60104 229796 60110
rect 229744 60046 229796 60052
rect 231136 13190 231164 98767
rect 231216 97912 231268 97918
rect 231216 97854 231268 97860
rect 231228 97617 231256 97854
rect 231214 97608 231270 97617
rect 231214 97543 231270 97552
rect 231214 96520 231270 96529
rect 231214 96455 231270 96464
rect 231228 28286 231256 96455
rect 231320 84930 231348 102847
rect 231596 102377 231624 103362
rect 232516 102882 232544 144910
rect 232596 131232 232648 131238
rect 232596 131174 232648 131180
rect 232504 102876 232556 102882
rect 232504 102818 232556 102824
rect 231582 102368 231638 102377
rect 231582 102303 231638 102312
rect 231676 102128 231728 102134
rect 231676 102070 231728 102076
rect 231400 102060 231452 102066
rect 231400 102002 231452 102008
rect 231412 101425 231440 102002
rect 231398 101416 231454 101425
rect 231398 101351 231454 101360
rect 231582 101416 231638 101425
rect 231582 101351 231638 101360
rect 231596 99521 231624 101351
rect 231688 100881 231716 102070
rect 231674 100872 231730 100881
rect 231674 100807 231730 100816
rect 231768 100700 231820 100706
rect 231768 100642 231820 100648
rect 231676 100632 231728 100638
rect 231676 100574 231728 100580
rect 231688 99929 231716 100574
rect 231780 100473 231808 100642
rect 231766 100464 231822 100473
rect 231766 100399 231822 100408
rect 231674 99920 231730 99929
rect 231674 99855 231730 99864
rect 231582 99512 231638 99521
rect 231582 99447 231638 99456
rect 231400 99340 231452 99346
rect 231400 99282 231452 99288
rect 231412 98569 231440 99282
rect 231398 98560 231454 98569
rect 231398 98495 231454 98504
rect 232504 95532 232556 95538
rect 232504 95474 232556 95480
rect 231308 84924 231360 84930
rect 231308 84866 231360 84872
rect 231216 28280 231268 28286
rect 231216 28222 231268 28228
rect 231124 13184 231176 13190
rect 231124 13126 231176 13132
rect 228456 4820 228508 4826
rect 228456 4762 228508 4768
rect 232516 4214 232544 95474
rect 232608 53145 232636 131174
rect 232700 114170 232728 154935
rect 232792 131170 232820 165582
rect 233528 161022 233556 212434
rect 233896 206961 233924 228239
rect 234448 212498 234476 240244
rect 235000 233209 235028 240244
rect 235262 237416 235318 237425
rect 235262 237351 235318 237360
rect 234986 233200 235042 233209
rect 234986 233135 235042 233144
rect 234618 225176 234674 225185
rect 234618 225111 234674 225120
rect 234436 212492 234488 212498
rect 234436 212434 234488 212440
rect 233882 206952 233938 206961
rect 233882 206887 233938 206896
rect 233896 205737 233924 206887
rect 233882 205728 233938 205737
rect 233882 205663 233938 205672
rect 233882 194168 233938 194177
rect 233882 194103 233938 194112
rect 233896 183025 233924 194103
rect 233976 191208 234028 191214
rect 233976 191150 234028 191156
rect 233882 183016 233938 183025
rect 233882 182951 233938 182960
rect 233988 181626 234016 191150
rect 233976 181620 234028 181626
rect 233976 181562 234028 181568
rect 233882 180024 233938 180033
rect 233882 179959 233938 179968
rect 233896 177342 233924 179959
rect 233884 177336 233936 177342
rect 233884 177278 233936 177284
rect 233884 176044 233936 176050
rect 233884 175986 233936 175992
rect 233516 161016 233568 161022
rect 233516 160958 233568 160964
rect 233896 158166 233924 175986
rect 233976 168428 234028 168434
rect 233976 168370 234028 168376
rect 233884 158160 233936 158166
rect 233884 158102 233936 158108
rect 233884 158024 233936 158030
rect 233884 157966 233936 157972
rect 233896 154873 233924 157966
rect 233882 154864 233938 154873
rect 233882 154799 233938 154808
rect 232872 146940 232924 146946
rect 232872 146882 232924 146888
rect 232884 133521 232912 146882
rect 233988 133618 234016 168370
rect 234066 166968 234122 166977
rect 234066 166903 234122 166912
rect 234080 154358 234108 166903
rect 234632 157185 234660 225111
rect 235276 220794 235304 237351
rect 235368 235958 235396 240244
rect 235920 238649 235948 240244
rect 236472 240145 236500 240244
rect 236458 240136 236514 240145
rect 236458 240071 236514 240080
rect 235906 238640 235962 238649
rect 235906 238575 235962 238584
rect 236644 238128 236696 238134
rect 236644 238070 236696 238076
rect 235356 235952 235408 235958
rect 235356 235894 235408 235900
rect 235264 220788 235316 220794
rect 235264 220730 235316 220736
rect 235276 207738 235304 220730
rect 236656 209098 236684 238070
rect 236840 226370 236868 240244
rect 237392 237425 237420 240244
rect 237944 240145 237972 240244
rect 237930 240136 237986 240145
rect 237930 240071 237986 240080
rect 237944 238754 237972 240071
rect 237944 238726 238064 238754
rect 237378 237416 237434 237425
rect 237378 237351 237434 237360
rect 236828 226364 236880 226370
rect 236828 226306 236880 226312
rect 236644 209092 236696 209098
rect 236644 209034 236696 209040
rect 235446 207904 235502 207913
rect 235446 207839 235502 207848
rect 235264 207732 235316 207738
rect 235264 207674 235316 207680
rect 235356 192568 235408 192574
rect 235356 192510 235408 192516
rect 234712 182912 234764 182918
rect 234712 182854 234764 182860
rect 234724 165578 234752 182854
rect 234896 181552 234948 181558
rect 234896 181494 234948 181500
rect 234804 178764 234856 178770
rect 234804 178706 234856 178712
rect 234816 167006 234844 178706
rect 234908 169454 234936 181494
rect 235368 181393 235396 192510
rect 235460 181490 235488 207839
rect 236276 207664 236328 207670
rect 236276 207606 236328 207612
rect 236182 181656 236238 181665
rect 236182 181591 236238 181600
rect 235448 181484 235500 181490
rect 235448 181426 235500 181432
rect 235354 181384 235410 181393
rect 235354 181319 235410 181328
rect 236090 178392 236146 178401
rect 236090 178327 236146 178336
rect 235998 170368 236054 170377
rect 235998 170303 236054 170312
rect 234896 169448 234948 169454
rect 234896 169390 234948 169396
rect 235264 167068 235316 167074
rect 235264 167010 235316 167016
rect 234804 167000 234856 167006
rect 234804 166942 234856 166948
rect 234712 165572 234764 165578
rect 234712 165514 234764 165520
rect 234618 157176 234674 157185
rect 234618 157111 234674 157120
rect 234068 154352 234120 154358
rect 234068 154294 234120 154300
rect 234160 153876 234212 153882
rect 234160 153818 234212 153824
rect 234068 145036 234120 145042
rect 234068 144978 234120 144984
rect 233976 133612 234028 133618
rect 233976 133554 234028 133560
rect 232870 133512 232926 133521
rect 232870 133447 232926 133456
rect 233884 132524 233936 132530
rect 233884 132466 233936 132472
rect 232780 131164 232832 131170
rect 232780 131106 232832 131112
rect 232778 116512 232834 116521
rect 232778 116447 232834 116456
rect 232688 114164 232740 114170
rect 232688 114106 232740 114112
rect 232686 98696 232742 98705
rect 232686 98631 232742 98640
rect 232594 53136 232650 53145
rect 232594 53071 232650 53080
rect 232700 22778 232728 98631
rect 232792 97986 232820 116447
rect 232870 102776 232926 102785
rect 232870 102711 232926 102720
rect 232780 97980 232832 97986
rect 232780 97922 232832 97928
rect 232884 83570 232912 102711
rect 232872 83564 232924 83570
rect 232872 83506 232924 83512
rect 232688 22772 232740 22778
rect 232688 22714 232740 22720
rect 233896 6254 233924 132466
rect 234080 103970 234108 144978
rect 234172 125594 234200 153818
rect 234344 140072 234396 140078
rect 234344 140014 234396 140020
rect 234160 125588 234212 125594
rect 234160 125530 234212 125536
rect 234250 123448 234306 123457
rect 234250 123383 234306 123392
rect 234160 113212 234212 113218
rect 234160 113154 234212 113160
rect 234068 103964 234120 103970
rect 234068 103906 234120 103912
rect 233976 103556 234028 103562
rect 233976 103498 234028 103504
rect 233988 29714 234016 103498
rect 234172 75177 234200 113154
rect 234264 94518 234292 123383
rect 234356 118726 234384 140014
rect 235276 127770 235304 167010
rect 236012 164014 236040 170303
rect 236000 164008 236052 164014
rect 236000 163950 236052 163956
rect 235538 163160 235594 163169
rect 235538 163095 235594 163104
rect 235446 153232 235502 153241
rect 235446 153167 235502 153176
rect 235356 129804 235408 129810
rect 235356 129746 235408 129752
rect 235264 127764 235316 127770
rect 235264 127706 235316 127712
rect 235264 124228 235316 124234
rect 235264 124170 235316 124176
rect 234344 118720 234396 118726
rect 234344 118662 234396 118668
rect 234252 94512 234304 94518
rect 234252 94454 234304 94460
rect 234158 75168 234214 75177
rect 234158 75103 234214 75112
rect 233976 29708 234028 29714
rect 233976 29650 234028 29656
rect 235276 25566 235304 124170
rect 235368 40730 235396 129746
rect 235460 111722 235488 153167
rect 235552 122641 235580 163095
rect 236104 140758 236132 178327
rect 236196 169794 236224 181591
rect 236184 169788 236236 169794
rect 236184 169730 236236 169736
rect 236288 167482 236316 207606
rect 237380 202156 237432 202162
rect 237380 202098 237432 202104
rect 236368 172508 236420 172514
rect 236368 172450 236420 172456
rect 236276 167476 236328 167482
rect 236276 167418 236328 167424
rect 236380 166705 236408 172450
rect 237392 171902 237420 202098
rect 237472 179988 237524 179994
rect 237472 179930 237524 179936
rect 237380 171896 237432 171902
rect 237380 171838 237432 171844
rect 236366 166696 236422 166705
rect 236366 166631 236422 166640
rect 236920 164892 236972 164898
rect 236920 164834 236972 164840
rect 236644 164280 236696 164286
rect 236644 164222 236696 164228
rect 236092 140752 236144 140758
rect 236092 140694 236144 140700
rect 236656 125089 236684 164222
rect 236826 157584 236882 157593
rect 236826 157519 236882 157528
rect 236734 136912 236790 136921
rect 236734 136847 236790 136856
rect 236642 125080 236698 125089
rect 236642 125015 236698 125024
rect 235538 122632 235594 122641
rect 235538 122567 235594 122576
rect 235538 120728 235594 120737
rect 235538 120663 235594 120672
rect 235448 111716 235500 111722
rect 235448 111658 235500 111664
rect 235552 86290 235580 120663
rect 236642 120184 236698 120193
rect 236642 120119 236698 120128
rect 235540 86284 235592 86290
rect 235540 86226 235592 86232
rect 235356 40724 235408 40730
rect 235356 40666 235408 40672
rect 235264 25560 235316 25566
rect 235264 25502 235316 25508
rect 233884 6248 233936 6254
rect 233884 6190 233936 6196
rect 236656 4865 236684 120119
rect 236748 57254 236776 136847
rect 236840 117230 236868 157519
rect 236932 129606 236960 164834
rect 237484 155446 237512 179930
rect 238036 172514 238064 238726
rect 238312 225622 238340 240244
rect 238864 233073 238892 240244
rect 239232 240009 239260 240244
rect 239218 240000 239274 240009
rect 239218 239935 239274 239944
rect 238944 238808 238996 238814
rect 238942 238776 238944 238785
rect 238996 238776 238998 238785
rect 238942 238711 238998 238720
rect 238850 233064 238906 233073
rect 238850 232999 238906 233008
rect 238300 225616 238352 225622
rect 238300 225558 238352 225564
rect 239784 224777 239812 240244
rect 240048 240032 240100 240038
rect 240048 239974 240100 239980
rect 240060 238814 240088 239974
rect 240048 238808 240100 238814
rect 240048 238750 240100 238756
rect 240336 234666 240364 240244
rect 240704 237017 240732 240244
rect 240876 240100 240928 240106
rect 240876 240042 240928 240048
rect 240690 237008 240746 237017
rect 240690 236943 240746 236952
rect 240324 234660 240376 234666
rect 240324 234602 240376 234608
rect 240784 234660 240836 234666
rect 240784 234602 240836 234608
rect 239770 224768 239826 224777
rect 239770 224703 239826 224712
rect 239404 209840 239456 209846
rect 239404 209782 239456 209788
rect 239416 199617 239444 209782
rect 240140 205624 240192 205630
rect 240140 205566 240192 205572
rect 239402 199608 239458 199617
rect 239402 199543 239458 199552
rect 238116 198824 238168 198830
rect 238116 198766 238168 198772
rect 238128 180130 238156 198766
rect 238850 187232 238906 187241
rect 238850 187167 238906 187176
rect 238760 184272 238812 184278
rect 238760 184214 238812 184220
rect 238116 180124 238168 180130
rect 238116 180066 238168 180072
rect 238298 174040 238354 174049
rect 238298 173975 238354 173984
rect 238024 172508 238076 172514
rect 238024 172450 238076 172456
rect 238116 171148 238168 171154
rect 238116 171090 238168 171096
rect 237472 155440 237524 155446
rect 237472 155382 237524 155388
rect 238024 151836 238076 151842
rect 238024 151778 238076 151784
rect 236920 129600 236972 129606
rect 236920 129542 236972 129548
rect 237012 128376 237064 128382
rect 237012 128318 237064 128324
rect 236828 117224 236880 117230
rect 236828 117166 236880 117172
rect 237024 98705 237052 128318
rect 238036 120154 238064 151778
rect 238128 133278 238156 171090
rect 238208 154624 238260 154630
rect 238208 154566 238260 154572
rect 238116 133272 238168 133278
rect 238116 133214 238168 133220
rect 238114 130112 238170 130121
rect 238114 130047 238170 130056
rect 238024 120148 238076 120154
rect 238024 120090 238076 120096
rect 238022 116920 238078 116929
rect 238022 116855 238078 116864
rect 237010 98696 237066 98705
rect 237010 98631 237066 98640
rect 236736 57248 236788 57254
rect 236736 57190 236788 57196
rect 238036 50289 238064 116855
rect 238128 76537 238156 130047
rect 238220 115870 238248 154566
rect 238312 137630 238340 173975
rect 238392 168564 238444 168570
rect 238392 168506 238444 168512
rect 238404 151910 238432 168506
rect 238392 151904 238444 151910
rect 238392 151846 238444 151852
rect 238772 144945 238800 184214
rect 238864 168570 238892 187167
rect 238944 177404 238996 177410
rect 238944 177346 238996 177352
rect 238852 168564 238904 168570
rect 238852 168506 238904 168512
rect 238956 165617 238984 177346
rect 240152 175234 240180 205566
rect 240796 185638 240824 234602
rect 240888 205630 240916 240042
rect 241256 234530 241284 240244
rect 241808 238649 241836 240244
rect 242176 238746 242204 240244
rect 242256 240168 242308 240174
rect 242256 240110 242308 240116
rect 242164 238740 242216 238746
rect 242164 238682 242216 238688
rect 241794 238640 241850 238649
rect 241794 238575 241850 238584
rect 241808 237561 241836 238575
rect 241794 237552 241850 237561
rect 241794 237487 241850 237496
rect 240968 234524 241020 234530
rect 240968 234466 241020 234472
rect 241244 234524 241296 234530
rect 241244 234466 241296 234472
rect 240980 213246 241008 234466
rect 240968 213240 241020 213246
rect 240968 213182 241020 213188
rect 241518 209128 241574 209137
rect 241518 209063 241574 209072
rect 240876 205624 240928 205630
rect 240876 205566 240928 205572
rect 240232 185632 240284 185638
rect 240232 185574 240284 185580
rect 240784 185632 240836 185638
rect 240784 185574 240836 185580
rect 240140 175228 240192 175234
rect 240140 175170 240192 175176
rect 239402 167104 239458 167113
rect 239402 167039 239458 167048
rect 238942 165608 238998 165617
rect 238942 165543 238998 165552
rect 238758 144936 238814 144945
rect 238758 144871 238814 144880
rect 238300 137624 238352 137630
rect 238300 137566 238352 137572
rect 239416 126954 239444 167039
rect 239680 165708 239732 165714
rect 239680 165650 239732 165656
rect 239496 154692 239548 154698
rect 239496 154634 239548 154640
rect 239404 126948 239456 126954
rect 239404 126890 239456 126896
rect 239402 124536 239458 124545
rect 239402 124471 239458 124480
rect 238208 115864 238260 115870
rect 238208 115806 238260 115812
rect 238114 76528 238170 76537
rect 238114 76463 238170 76472
rect 238022 50280 238078 50289
rect 238022 50215 238078 50224
rect 238022 46200 238078 46209
rect 238022 46135 238078 46144
rect 238036 6186 238064 46135
rect 239416 15910 239444 124471
rect 239508 114510 239536 154634
rect 239692 135998 239720 165650
rect 240244 161430 240272 185574
rect 240324 180260 240376 180266
rect 240324 180202 240376 180208
rect 240232 161424 240284 161430
rect 240232 161366 240284 161372
rect 240336 156670 240364 180202
rect 240876 171216 240928 171222
rect 240876 171158 240928 171164
rect 240784 160132 240836 160138
rect 240784 160074 240836 160080
rect 240324 156664 240376 156670
rect 240324 156606 240376 156612
rect 239680 135992 239732 135998
rect 239680 135934 239732 135940
rect 239588 135924 239640 135930
rect 239588 135866 239640 135872
rect 239496 114504 239548 114510
rect 239496 114446 239548 114452
rect 239600 102066 239628 135866
rect 240796 124914 240824 160074
rect 240888 152425 240916 171158
rect 240968 169788 241020 169794
rect 240968 169730 241020 169736
rect 240874 152416 240930 152425
rect 240874 152351 240930 152360
rect 240874 149424 240930 149433
rect 240874 149359 240930 149368
rect 240784 124908 240836 124914
rect 240784 124850 240836 124856
rect 240784 120148 240836 120154
rect 240784 120090 240836 120096
rect 239678 104000 239734 104009
rect 239678 103935 239734 103944
rect 239588 102060 239640 102066
rect 239588 102002 239640 102008
rect 239494 98696 239550 98705
rect 239494 98631 239550 98640
rect 239508 42090 239536 98631
rect 239692 90438 239720 103935
rect 239680 90432 239732 90438
rect 239680 90374 239732 90380
rect 240138 42120 240194 42129
rect 239496 42084 239548 42090
rect 240138 42055 240194 42064
rect 239496 42026 239548 42032
rect 239404 15904 239456 15910
rect 239404 15846 239456 15852
rect 238024 6180 238076 6186
rect 238024 6122 238076 6128
rect 236642 4856 236698 4865
rect 236642 4791 236698 4800
rect 232504 4208 232556 4214
rect 232504 4150 232556 4156
rect 235816 4208 235868 4214
rect 235816 4150 235868 4156
rect 222844 2100 222896 2106
rect 222844 2042 222896 2048
rect 195242 2000 195298 2009
rect 195242 1935 195298 1944
rect 235828 480 235856 4150
rect 239310 2136 239366 2145
rect 239310 2071 239366 2080
rect 239324 480 239352 2071
rect 240152 490 240180 42055
rect 240796 17270 240824 120090
rect 240888 107545 240916 149359
rect 240980 147014 241008 169730
rect 241060 155984 241112 155990
rect 241060 155926 241112 155932
rect 240968 147008 241020 147014
rect 240968 146950 241020 146956
rect 240968 143608 241020 143614
rect 240968 143550 241020 143556
rect 240874 107536 240930 107545
rect 240874 107471 240930 107480
rect 240980 103426 241008 143550
rect 241072 117978 241100 155926
rect 241532 146985 241560 209063
rect 241610 198248 241666 198257
rect 241610 198183 241666 198192
rect 241624 168609 241652 198183
rect 242176 186425 242204 238682
rect 242268 216209 242296 240110
rect 242728 235793 242756 240244
rect 242714 235784 242770 235793
rect 242714 235719 242770 235728
rect 243280 228313 243308 240244
rect 243648 238921 243676 240244
rect 243924 240106 243952 240479
rect 243912 240100 243964 240106
rect 243912 240042 243964 240048
rect 243634 238912 243690 238921
rect 243634 238847 243690 238856
rect 243648 235278 243676 238847
rect 244016 238754 244044 248367
rect 244370 245168 244426 245177
rect 244370 245103 244426 245112
rect 244094 241360 244150 241369
rect 244094 241295 244150 241304
rect 244108 240174 244136 241295
rect 244096 240168 244148 240174
rect 244096 240110 244148 240116
rect 243924 238726 244044 238754
rect 243636 235272 243688 235278
rect 243636 235214 243688 235220
rect 243266 228304 243322 228313
rect 243266 228239 243322 228248
rect 242900 219428 242952 219434
rect 242900 219370 242952 219376
rect 242912 218822 242940 219370
rect 243924 218822 243952 238726
rect 244280 224936 244332 224942
rect 244280 224878 244332 224884
rect 244292 224777 244320 224878
rect 244278 224768 244334 224777
rect 244278 224703 244334 224712
rect 242900 218816 242952 218822
rect 242900 218758 242952 218764
rect 243912 218816 243964 218822
rect 243912 218758 243964 218764
rect 242254 216200 242310 216209
rect 242254 216135 242310 216144
rect 242162 186416 242218 186425
rect 242162 186351 242218 186360
rect 241702 184376 241758 184385
rect 241702 184311 241758 184320
rect 241610 168600 241666 168609
rect 241610 168535 241666 168544
rect 241716 162178 241744 184311
rect 242256 182844 242308 182850
rect 242256 182786 242308 182792
rect 242164 167136 242216 167142
rect 242164 167078 242216 167084
rect 241704 162172 241756 162178
rect 241704 162114 241756 162120
rect 241518 146976 241574 146985
rect 241518 146911 241574 146920
rect 242176 128314 242204 167078
rect 242268 158030 242296 182786
rect 242256 158024 242308 158030
rect 242256 157966 242308 157972
rect 242254 156632 242310 156641
rect 242254 156567 242310 156576
rect 242164 128308 242216 128314
rect 242164 128250 242216 128256
rect 241060 117972 241112 117978
rect 241060 117914 241112 117920
rect 242164 117360 242216 117366
rect 242164 117302 242216 117308
rect 241058 106312 241114 106321
rect 241058 106247 241114 106256
rect 240968 103420 241020 103426
rect 240968 103362 241020 103368
rect 241072 75313 241100 106247
rect 241520 77988 241572 77994
rect 241520 77930 241572 77936
rect 241058 75304 241114 75313
rect 241058 75239 241114 75248
rect 240784 17264 240836 17270
rect 240784 17206 240836 17212
rect 241532 16574 241560 77930
rect 242176 36582 242204 117302
rect 242268 117298 242296 156567
rect 242440 150476 242492 150482
rect 242440 150418 242492 150424
rect 242346 145344 242402 145353
rect 242346 145279 242402 145288
rect 242360 118017 242388 145279
rect 242346 118008 242402 118017
rect 242346 117943 242402 117952
rect 242256 117292 242308 117298
rect 242256 117234 242308 117240
rect 242348 114572 242400 114578
rect 242348 114514 242400 114520
rect 242254 109440 242310 109449
rect 242254 109375 242310 109384
rect 242268 54534 242296 109375
rect 242360 69601 242388 114514
rect 242452 110362 242480 150418
rect 242912 144226 242940 218758
rect 244384 213858 244412 245103
rect 244464 242956 244516 242962
rect 244464 242898 244516 242904
rect 244476 238066 244504 242898
rect 244464 238060 244516 238066
rect 244464 238002 244516 238008
rect 244372 213852 244424 213858
rect 244372 213794 244424 213800
rect 244384 209774 244412 213794
rect 244568 212430 244596 264415
rect 245844 264036 245896 264042
rect 245844 263978 245896 263984
rect 245856 263945 245884 263978
rect 245842 263936 245898 263945
rect 245842 263871 245898 263880
rect 245658 263120 245714 263129
rect 245658 263055 245714 263064
rect 245672 259978 245700 263055
rect 245752 260772 245804 260778
rect 245752 260714 245804 260720
rect 245764 260137 245792 260714
rect 245750 260128 245806 260137
rect 245750 260063 245806 260072
rect 245672 259950 245792 259978
rect 245660 258052 245712 258058
rect 245660 257994 245712 258000
rect 245672 257417 245700 257994
rect 245658 257408 245714 257417
rect 245658 257343 245714 257352
rect 245658 253056 245714 253065
rect 245658 252991 245714 253000
rect 245672 250578 245700 252991
rect 245660 250572 245712 250578
rect 245660 250514 245712 250520
rect 245106 250336 245162 250345
rect 245106 250271 245162 250280
rect 244646 243808 244702 243817
rect 244646 243743 244702 243752
rect 244660 242962 244688 243743
rect 244648 242956 244700 242962
rect 244648 242898 244700 242904
rect 245120 242214 245148 250271
rect 245108 242208 245160 242214
rect 245108 242150 245160 242156
rect 245764 221649 245792 259950
rect 245936 259412 245988 259418
rect 245936 259354 245988 259360
rect 245842 258768 245898 258777
rect 245842 258703 245898 258712
rect 245856 258126 245884 258703
rect 245948 258233 245976 259354
rect 245934 258224 245990 258233
rect 245934 258159 245990 258168
rect 245844 258120 245896 258126
rect 245844 258062 245896 258068
rect 245936 256624 245988 256630
rect 245934 256592 245936 256601
rect 245988 256592 245990 256601
rect 245934 256527 245990 256536
rect 245844 255264 245896 255270
rect 245844 255206 245896 255212
rect 245934 255232 245990 255241
rect 245856 254425 245884 255206
rect 245934 255167 245936 255176
rect 245988 255167 245990 255176
rect 245936 255138 245988 255144
rect 245842 254416 245898 254425
rect 245842 254351 245898 254360
rect 245936 253904 245988 253910
rect 245934 253872 245936 253881
rect 245988 253872 245990 253881
rect 245934 253807 245990 253816
rect 245844 252544 245896 252550
rect 245844 252486 245896 252492
rect 245856 251705 245884 252486
rect 245936 252340 245988 252346
rect 245936 252282 245988 252288
rect 245948 252249 245976 252282
rect 245934 252240 245990 252249
rect 245934 252175 245990 252184
rect 245842 251696 245898 251705
rect 245842 251631 245898 251640
rect 245936 249688 245988 249694
rect 245936 249630 245988 249636
rect 245948 249529 245976 249630
rect 245934 249520 245990 249529
rect 245934 249455 245990 249464
rect 245934 248160 245990 248169
rect 245934 248095 245990 248104
rect 245948 247722 245976 248095
rect 245936 247716 245988 247722
rect 245936 247658 245988 247664
rect 245842 246528 245898 246537
rect 245842 246463 245898 246472
rect 245856 245682 245884 246463
rect 245844 245676 245896 245682
rect 245844 245618 245896 245624
rect 245948 245562 245976 247658
rect 245856 245534 245976 245562
rect 245856 235929 245884 245534
rect 245934 244624 245990 244633
rect 245934 244559 245990 244568
rect 245948 244458 245976 244559
rect 245936 244452 245988 244458
rect 245936 244394 245988 244400
rect 245934 242448 245990 242457
rect 245934 242383 245990 242392
rect 245948 241534 245976 242383
rect 245936 241528 245988 241534
rect 245936 241470 245988 241476
rect 245842 235920 245898 235929
rect 245842 235855 245898 235864
rect 245844 225616 245896 225622
rect 245844 225558 245896 225564
rect 245750 221640 245806 221649
rect 245750 221575 245806 221584
rect 244556 212424 244608 212430
rect 244556 212366 244608 212372
rect 244292 209746 244412 209774
rect 242990 205184 243046 205193
rect 242990 205119 243046 205128
rect 243004 204950 243032 205119
rect 242992 204944 243044 204950
rect 242992 204886 243044 204892
rect 243004 157350 243032 204886
rect 243544 175364 243596 175370
rect 243544 175306 243596 175312
rect 242992 157344 243044 157350
rect 242992 157286 243044 157292
rect 242900 144220 242952 144226
rect 242900 144162 242952 144168
rect 242440 110356 242492 110362
rect 242440 110298 242492 110304
rect 243556 99278 243584 175306
rect 243634 160440 243690 160449
rect 243634 160375 243690 160384
rect 243648 119785 243676 160375
rect 244292 150346 244320 209746
rect 244568 200114 244596 212366
rect 245856 204241 245884 225558
rect 245842 204232 245898 204241
rect 245842 204167 245898 204176
rect 244384 200086 244596 200114
rect 244384 172417 244412 200086
rect 244464 189848 244516 189854
rect 244464 189790 244516 189796
rect 244370 172408 244426 172417
rect 244370 172343 244426 172352
rect 244476 151774 244504 189790
rect 245752 181620 245804 181626
rect 245752 181562 245804 181568
rect 244554 178120 244610 178129
rect 244554 178055 244610 178064
rect 244568 160002 244596 178055
rect 245200 162920 245252 162926
rect 245200 162862 245252 162868
rect 244556 159996 244608 160002
rect 244556 159938 244608 159944
rect 244924 159384 244976 159390
rect 244924 159326 244976 159332
rect 244464 151768 244516 151774
rect 244464 151710 244516 151716
rect 244280 150340 244332 150346
rect 244280 150282 244332 150288
rect 243820 144220 243872 144226
rect 243820 144162 243872 144168
rect 243634 119776 243690 119785
rect 243634 119711 243690 119720
rect 243726 107944 243782 107953
rect 243726 107879 243782 107888
rect 243634 102232 243690 102241
rect 243634 102167 243690 102176
rect 243544 99272 243596 99278
rect 243544 99214 243596 99220
rect 242346 69592 242402 69601
rect 242346 69527 242402 69536
rect 242256 54528 242308 54534
rect 242256 54470 242308 54476
rect 242164 36576 242216 36582
rect 242164 36518 242216 36524
rect 243648 31074 243676 102167
rect 243740 55894 243768 107879
rect 243832 104854 243860 144162
rect 244936 122738 244964 159326
rect 245108 149116 245160 149122
rect 245108 149058 245160 149064
rect 245014 142488 245070 142497
rect 245014 142423 245070 142432
rect 244924 122732 244976 122738
rect 244924 122674 244976 122680
rect 244924 110492 244976 110498
rect 244924 110434 244976 110440
rect 243820 104848 243872 104854
rect 243820 104790 243872 104796
rect 244278 96520 244334 96529
rect 244278 96455 244334 96464
rect 244292 95674 244320 96455
rect 244280 95668 244332 95674
rect 244280 95610 244332 95616
rect 243728 55888 243780 55894
rect 243728 55830 243780 55836
rect 244936 47666 244964 110434
rect 245028 100638 245056 142423
rect 245120 108934 245148 149058
rect 245212 142769 245240 162862
rect 245764 144809 245792 181562
rect 245844 178696 245896 178702
rect 245844 178638 245896 178644
rect 245856 154562 245884 178638
rect 245936 175976 245988 175982
rect 245936 175918 245988 175924
rect 245948 161537 245976 175918
rect 246040 164937 246068 277366
rect 246408 272241 246436 298726
rect 247052 283218 247080 336806
rect 247316 306400 247368 306406
rect 247316 306342 247368 306348
rect 247222 290184 247278 290193
rect 247222 290119 247278 290128
rect 247040 283212 247092 283218
rect 247040 283154 247092 283160
rect 246486 274544 246542 274553
rect 246486 274479 246542 274488
rect 246118 272232 246174 272241
rect 246118 272167 246174 272176
rect 246394 272232 246450 272241
rect 246394 272167 246450 272176
rect 246132 271017 246160 272167
rect 246118 271008 246174 271017
rect 246118 270943 246174 270952
rect 246302 270192 246358 270201
rect 246302 270127 246358 270136
rect 246316 269890 246344 270127
rect 246304 269884 246356 269890
rect 246304 269826 246356 269832
rect 246500 264246 246528 274479
rect 247040 269884 247092 269890
rect 247040 269826 247092 269832
rect 246488 264240 246540 264246
rect 246488 264182 246540 264188
rect 246396 261588 246448 261594
rect 246396 261530 246448 261536
rect 246408 260953 246436 261530
rect 246394 260944 246450 260953
rect 246394 260879 246450 260888
rect 246394 245984 246450 245993
rect 246394 245919 246450 245928
rect 246408 245750 246436 245919
rect 246396 245744 246448 245750
rect 246396 245686 246448 245692
rect 246304 221536 246356 221542
rect 246304 221478 246356 221484
rect 246316 179450 246344 221478
rect 246394 204232 246450 204241
rect 246394 204167 246450 204176
rect 246304 179444 246356 179450
rect 246304 179386 246356 179392
rect 246408 175982 246436 204167
rect 246396 175976 246448 175982
rect 246396 175918 246448 175924
rect 247052 173874 247080 269826
rect 247130 262304 247186 262313
rect 247130 262239 247186 262248
rect 247144 202162 247172 262239
rect 247236 256057 247264 290119
rect 247328 279002 247356 306342
rect 247408 289876 247460 289882
rect 247408 289818 247460 289824
rect 247316 278996 247368 279002
rect 247316 278938 247368 278944
rect 247420 261594 247448 289818
rect 248432 264042 248460 368455
rect 255412 356108 255464 356114
rect 255412 356050 255464 356056
rect 251272 351960 251324 351966
rect 251272 351902 251324 351908
rect 249892 350600 249944 350606
rect 249892 350542 249944 350548
rect 248604 329112 248656 329118
rect 248604 329054 248656 329060
rect 248512 319456 248564 319462
rect 248512 319398 248564 319404
rect 248420 264036 248472 264042
rect 248420 263978 248472 263984
rect 247408 261588 247460 261594
rect 247408 261530 247460 261536
rect 248420 261588 248472 261594
rect 248420 261530 248472 261536
rect 247222 256048 247278 256057
rect 247222 255983 247278 255992
rect 247224 245744 247276 245750
rect 247224 245686 247276 245692
rect 247236 231577 247264 245686
rect 247222 231568 247278 231577
rect 247222 231503 247278 231512
rect 247132 202156 247184 202162
rect 247132 202098 247184 202104
rect 247684 200184 247736 200190
rect 247684 200126 247736 200132
rect 247224 186992 247276 186998
rect 247224 186934 247276 186940
rect 247132 179444 247184 179450
rect 247132 179386 247184 179392
rect 247040 173868 247092 173874
rect 247040 173810 247092 173816
rect 246026 164928 246082 164937
rect 246026 164863 246082 164872
rect 245934 161528 245990 161537
rect 245934 161463 245990 161472
rect 246488 161492 246540 161498
rect 246488 161434 246540 161440
rect 246396 160200 246448 160206
rect 246396 160142 246448 160148
rect 245844 154556 245896 154562
rect 245844 154498 245896 154504
rect 245750 144800 245806 144809
rect 245750 144735 245806 144744
rect 245198 142760 245254 142769
rect 245198 142695 245254 142704
rect 246304 127016 246356 127022
rect 246304 126958 246356 126964
rect 245108 108928 245160 108934
rect 245108 108870 245160 108876
rect 245106 103728 245162 103737
rect 245106 103663 245162 103672
rect 245016 100632 245068 100638
rect 245016 100574 245068 100580
rect 245014 98832 245070 98841
rect 245014 98767 245070 98776
rect 244924 47660 244976 47666
rect 244924 47602 244976 47608
rect 245028 46238 245056 98767
rect 245120 89078 245148 103663
rect 245200 99408 245252 99414
rect 245200 99350 245252 99356
rect 245108 89072 245160 89078
rect 245108 89014 245160 89020
rect 245212 84862 245240 99350
rect 245200 84856 245252 84862
rect 245200 84798 245252 84804
rect 246316 59945 246344 126958
rect 246408 120057 246436 160142
rect 246500 121446 246528 161434
rect 247144 150414 247172 179386
rect 247236 162858 247264 186934
rect 247696 178809 247724 200126
rect 247682 178800 247738 178809
rect 247682 178735 247738 178744
rect 247776 173936 247828 173942
rect 247776 173878 247828 173884
rect 247684 172576 247736 172582
rect 247684 172518 247736 172524
rect 247224 162852 247276 162858
rect 247224 162794 247276 162800
rect 247132 150408 247184 150414
rect 247132 150350 247184 150356
rect 247696 135182 247724 172518
rect 247788 136610 247816 173878
rect 247868 151904 247920 151910
rect 247868 151846 247920 151852
rect 247776 136604 247828 136610
rect 247776 136546 247828 136552
rect 247684 135176 247736 135182
rect 247684 135118 247736 135124
rect 246578 134464 246634 134473
rect 246578 134399 246634 134408
rect 246488 121440 246540 121446
rect 246488 121382 246540 121388
rect 246394 120048 246450 120057
rect 246394 119983 246450 119992
rect 246396 100768 246448 100774
rect 246396 100710 246448 100716
rect 246302 59936 246358 59945
rect 246302 59871 246358 59880
rect 245016 46232 245068 46238
rect 245016 46174 245068 46180
rect 246408 43450 246436 100710
rect 246592 99346 246620 134399
rect 247684 132592 247736 132598
rect 247684 132534 247736 132540
rect 246580 99340 246632 99346
rect 246580 99282 246632 99288
rect 246486 95296 246542 95305
rect 246486 95231 246542 95240
rect 246500 79529 246528 95231
rect 246486 79520 246542 79529
rect 246486 79455 246542 79464
rect 247696 65657 247724 132534
rect 247880 111790 247908 151846
rect 248432 148374 248460 261530
rect 248524 238746 248552 319398
rect 248616 280838 248644 329054
rect 249800 327140 249852 327146
rect 249800 327082 249852 327088
rect 248694 294672 248750 294681
rect 248694 294607 248750 294616
rect 248604 280832 248656 280838
rect 248604 280774 248656 280780
rect 248708 252346 248736 294607
rect 249812 278118 249840 327082
rect 249800 278112 249852 278118
rect 249800 278054 249852 278060
rect 249800 255196 249852 255202
rect 249800 255138 249852 255144
rect 248696 252340 248748 252346
rect 248696 252282 248748 252288
rect 249812 248414 249840 255138
rect 249904 249694 249932 350542
rect 249982 291272 250038 291281
rect 249982 291207 250038 291216
rect 249996 278050 250024 291207
rect 251284 283529 251312 351902
rect 252652 342304 252704 342310
rect 252652 342246 252704 342252
rect 251362 338328 251418 338337
rect 251362 338263 251418 338272
rect 251270 283520 251326 283529
rect 251270 283455 251326 283464
rect 250076 283212 250128 283218
rect 250076 283154 250128 283160
rect 249984 278044 250036 278050
rect 249984 277986 250036 277992
rect 249892 249688 249944 249694
rect 249892 249630 249944 249636
rect 249812 248386 249932 248414
rect 248604 245676 248656 245682
rect 248604 245618 248656 245624
rect 248512 238740 248564 238746
rect 248512 238682 248564 238688
rect 248616 195945 248644 245618
rect 248696 244452 248748 244458
rect 248696 244394 248748 244400
rect 248708 207670 248736 244394
rect 249904 234598 249932 248386
rect 249892 234592 249944 234598
rect 249892 234534 249944 234540
rect 248696 207664 248748 207670
rect 248696 207606 248748 207612
rect 248602 195936 248658 195945
rect 248602 195871 248658 195880
rect 248510 189136 248566 189145
rect 248510 189071 248566 189080
rect 248524 156233 248552 189071
rect 248604 181484 248656 181490
rect 248604 181426 248656 181432
rect 248510 156224 248566 156233
rect 248510 156159 248566 156168
rect 248616 151065 248644 181426
rect 249248 169856 249300 169862
rect 249248 169798 249300 169804
rect 248602 151056 248658 151065
rect 248602 150991 248658 151000
rect 249154 150784 249210 150793
rect 249154 150719 249210 150728
rect 248420 148368 248472 148374
rect 248420 148310 248472 148316
rect 249062 132560 249118 132569
rect 249062 132495 249118 132504
rect 247958 123584 248014 123593
rect 247958 123519 248014 123528
rect 247868 111784 247920 111790
rect 247868 111726 247920 111732
rect 247774 110800 247830 110809
rect 247774 110735 247830 110744
rect 247682 65648 247738 65657
rect 247682 65583 247738 65592
rect 247788 51921 247816 110735
rect 247972 87650 248000 123519
rect 247960 87644 248012 87650
rect 247960 87586 248012 87592
rect 248418 71088 248474 71097
rect 248418 71023 248474 71032
rect 247774 51912 247830 51921
rect 247774 51847 247830 51856
rect 246396 43444 246448 43450
rect 246396 43386 246448 43392
rect 243636 31068 243688 31074
rect 243636 31010 243688 31016
rect 241532 16546 241744 16574
rect 240336 598 240548 626
rect 240336 490 240364 598
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240152 462 240364 490
rect 240520 480 240548 598
rect 241716 480 241744 16546
rect 245200 11824 245252 11830
rect 245200 11766 245252 11772
rect 244096 10328 244148 10334
rect 244096 10270 244148 10276
rect 242900 9036 242952 9042
rect 242900 8978 242952 8984
rect 242912 480 242940 8978
rect 244108 480 244136 10270
rect 245212 480 245240 11766
rect 246394 3632 246450 3641
rect 246394 3567 246450 3576
rect 246408 480 246436 3567
rect 247590 3496 247646 3505
rect 247590 3431 247646 3440
rect 247604 480 247632 3431
rect 248432 490 248460 71023
rect 249076 68377 249104 132495
rect 249168 109041 249196 150719
rect 249260 131102 249288 169798
rect 249904 164218 249932 234534
rect 249892 164212 249944 164218
rect 249892 164154 249944 164160
rect 249432 146668 249484 146674
rect 249432 146610 249484 146616
rect 249248 131096 249300 131102
rect 249248 131038 249300 131044
rect 249340 126336 249392 126342
rect 249340 126278 249392 126284
rect 249248 113280 249300 113286
rect 249248 113222 249300 113228
rect 249154 109032 249210 109041
rect 249154 108967 249210 108976
rect 249260 73817 249288 113222
rect 249352 90409 249380 126278
rect 249444 126274 249472 146610
rect 250088 143546 250116 283154
rect 251272 279472 251324 279478
rect 251272 279414 251324 279420
rect 251284 278905 251312 279414
rect 251270 278896 251326 278905
rect 251270 278831 251326 278840
rect 251284 278798 251312 278831
rect 251272 278792 251324 278798
rect 251272 278734 251324 278740
rect 251272 271924 251324 271930
rect 251272 271866 251324 271872
rect 251180 177336 251232 177342
rect 251180 177278 251232 177284
rect 250536 172644 250588 172650
rect 250536 172586 250588 172592
rect 250444 156052 250496 156058
rect 250444 155994 250496 156000
rect 250076 143540 250128 143546
rect 250076 143482 250128 143488
rect 249432 126268 249484 126274
rect 249432 126210 249484 126216
rect 250456 115841 250484 155994
rect 250548 133657 250576 172586
rect 250628 162988 250680 162994
rect 250628 162930 250680 162936
rect 250534 133648 250590 133657
rect 250534 133583 250590 133592
rect 250640 124098 250668 162930
rect 251192 142866 251220 177278
rect 251284 160070 251312 271866
rect 251376 265674 251404 338263
rect 251454 293992 251510 294001
rect 251454 293927 251510 293936
rect 251364 265668 251416 265674
rect 251364 265610 251416 265616
rect 251376 262886 251404 265610
rect 251364 262880 251416 262886
rect 251364 262822 251416 262828
rect 251468 260778 251496 293927
rect 252558 292768 252614 292777
rect 252558 292703 252614 292712
rect 251546 292632 251602 292641
rect 251546 292567 251602 292576
rect 251456 260772 251508 260778
rect 251456 260714 251508 260720
rect 251560 170377 251588 292567
rect 251824 193928 251876 193934
rect 251824 193870 251876 193876
rect 251836 181490 251864 193870
rect 251824 181484 251876 181490
rect 251824 181426 251876 181432
rect 251546 170368 251602 170377
rect 251546 170303 251602 170312
rect 251822 165744 251878 165753
rect 251822 165679 251878 165688
rect 251272 160064 251324 160070
rect 251272 160006 251324 160012
rect 251180 142860 251232 142866
rect 251180 142802 251232 142808
rect 250720 138712 250772 138718
rect 250720 138654 250772 138660
rect 250628 124092 250680 124098
rect 250628 124034 250680 124040
rect 250442 115832 250498 115841
rect 250442 115767 250498 115776
rect 250442 108080 250498 108089
rect 250442 108015 250498 108024
rect 249800 95668 249852 95674
rect 249800 95610 249852 95616
rect 249812 93838 249840 95610
rect 249800 93832 249852 93838
rect 249800 93774 249852 93780
rect 249338 90400 249394 90409
rect 249338 90335 249394 90344
rect 249246 73808 249302 73817
rect 249246 73743 249302 73752
rect 249062 68368 249118 68377
rect 249062 68303 249118 68312
rect 250456 58682 250484 108015
rect 250536 107704 250588 107710
rect 250536 107646 250588 107652
rect 250548 67017 250576 107646
rect 250732 107574 250760 138654
rect 251836 129033 251864 165679
rect 252572 158001 252600 292703
rect 252664 269890 252692 342246
rect 254032 316056 254084 316062
rect 254032 315998 254084 316004
rect 253204 299600 253256 299606
rect 253204 299542 253256 299548
rect 252836 270564 252888 270570
rect 252836 270506 252888 270512
rect 252652 269884 252704 269890
rect 252652 269826 252704 269832
rect 252744 242208 252796 242214
rect 252744 242150 252796 242156
rect 252756 229090 252784 242150
rect 252848 240106 252876 270506
rect 253216 259554 253244 299542
rect 253940 291304 253992 291310
rect 253940 291246 253992 291252
rect 253204 259548 253256 259554
rect 253204 259490 253256 259496
rect 253216 259418 253244 259490
rect 253204 259412 253256 259418
rect 253204 259354 253256 259360
rect 252836 240100 252888 240106
rect 252836 240042 252888 240048
rect 252928 235952 252980 235958
rect 252926 235920 252928 235929
rect 252980 235920 252982 235929
rect 252926 235855 252982 235864
rect 252940 234666 252968 235855
rect 252928 234660 252980 234666
rect 252928 234602 252980 234608
rect 252744 229084 252796 229090
rect 252744 229026 252796 229032
rect 252756 228410 252784 229026
rect 252744 228404 252796 228410
rect 252744 228346 252796 228352
rect 252652 202224 252704 202230
rect 252652 202166 252704 202172
rect 252558 157992 252614 158001
rect 252558 157927 252614 157936
rect 251916 157412 251968 157418
rect 251916 157354 251968 157360
rect 251822 129024 251878 129033
rect 251822 128959 251878 128968
rect 250812 127628 250864 127634
rect 250812 127570 250864 127576
rect 250720 107568 250772 107574
rect 250720 107510 250772 107516
rect 250824 102921 250852 127570
rect 251928 118658 251956 157354
rect 252008 149728 252060 149734
rect 252008 149670 252060 149676
rect 251916 118652 251968 118658
rect 251916 118594 251968 118600
rect 251822 117600 251878 117609
rect 251822 117535 251878 117544
rect 250810 102912 250866 102921
rect 250810 102847 250866 102856
rect 250628 102196 250680 102202
rect 250628 102138 250680 102144
rect 250640 93129 250668 102138
rect 250626 93120 250682 93129
rect 250626 93055 250682 93064
rect 250534 67008 250590 67017
rect 250534 66943 250590 66952
rect 250444 58676 250496 58682
rect 250444 58618 250496 58624
rect 249800 44872 249852 44878
rect 249800 44814 249852 44820
rect 249812 16574 249840 44814
rect 251836 35222 251864 117535
rect 252020 110430 252048 149670
rect 252664 137970 252692 202166
rect 253952 182850 253980 291246
rect 254044 276010 254072 315998
rect 254124 297492 254176 297498
rect 254124 297434 254176 297440
rect 254136 282878 254164 297434
rect 255320 287088 255372 287094
rect 255320 287030 255372 287036
rect 254124 282872 254176 282878
rect 254124 282814 254176 282820
rect 254032 276004 254084 276010
rect 254032 275946 254084 275952
rect 254032 273284 254084 273290
rect 254032 273226 254084 273232
rect 253940 182844 253992 182850
rect 253940 182786 253992 182792
rect 254044 176633 254072 273226
rect 254030 176624 254086 176633
rect 254030 176559 254086 176568
rect 253940 175976 253992 175982
rect 253940 175918 253992 175924
rect 253952 175302 253980 175918
rect 253940 175296 253992 175302
rect 253940 175238 253992 175244
rect 253202 168464 253258 168473
rect 253202 168399 253258 168408
rect 252652 137964 252704 137970
rect 252652 137906 252704 137912
rect 253216 128353 253244 168399
rect 253296 158024 253348 158030
rect 253296 157966 253348 157972
rect 253202 128344 253258 128353
rect 253202 128279 253258 128288
rect 252100 121508 252152 121514
rect 252100 121450 252152 121456
rect 252008 110424 252060 110430
rect 252008 110366 252060 110372
rect 251916 106344 251968 106350
rect 251916 106286 251968 106292
rect 251928 60042 251956 106286
rect 252112 86193 252140 121450
rect 253308 120086 253336 157966
rect 253480 147688 253532 147694
rect 253480 147630 253532 147636
rect 253296 120080 253348 120086
rect 253296 120022 253348 120028
rect 253204 117428 253256 117434
rect 253204 117370 253256 117376
rect 252098 86184 252154 86193
rect 252098 86119 252154 86128
rect 251916 60036 251968 60042
rect 251916 59978 251968 59984
rect 251824 35216 251876 35222
rect 251824 35158 251876 35164
rect 249812 16546 250024 16574
rect 248616 598 248828 626
rect 248616 490 248644 598
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248432 462 248644 490
rect 248800 480 248828 598
rect 249996 480 250024 16546
rect 253216 13122 253244 117370
rect 253296 116000 253348 116006
rect 253296 115942 253348 115948
rect 253308 37942 253336 115942
rect 253492 107642 253520 147630
rect 253480 107636 253532 107642
rect 253480 107578 253532 107584
rect 253388 106412 253440 106418
rect 253388 106354 253440 106360
rect 253400 61402 253428 106354
rect 253952 105602 253980 175238
rect 254674 172816 254730 172825
rect 254674 172751 254730 172760
rect 254582 170232 254638 170241
rect 254582 170167 254638 170176
rect 254596 141506 254624 170167
rect 254688 146946 254716 172751
rect 255332 149054 255360 287030
rect 255424 269074 255452 356050
rect 255504 325032 255556 325038
rect 255504 324974 255556 324980
rect 255412 269068 255464 269074
rect 255412 269010 255464 269016
rect 255424 268394 255452 269010
rect 255412 268388 255464 268394
rect 255412 268330 255464 268336
rect 255516 255270 255544 324974
rect 256700 303680 256752 303686
rect 256700 303622 256752 303628
rect 255596 302252 255648 302258
rect 255596 302194 255648 302200
rect 255608 258058 255636 302194
rect 255596 258052 255648 258058
rect 255596 257994 255648 258000
rect 255608 257378 255636 257994
rect 255596 257372 255648 257378
rect 255596 257314 255648 257320
rect 255504 255264 255556 255270
rect 255504 255206 255556 255212
rect 255504 241528 255556 241534
rect 255504 241470 255556 241476
rect 255412 221468 255464 221474
rect 255412 221410 255464 221416
rect 255320 149048 255372 149054
rect 255320 148990 255372 148996
rect 254676 146940 254728 146946
rect 254676 146882 254728 146888
rect 254676 142180 254728 142186
rect 254676 142122 254728 142128
rect 254584 141500 254636 141506
rect 254584 141442 254636 141448
rect 254584 136672 254636 136678
rect 254584 136614 254636 136620
rect 254596 123457 254624 136614
rect 254582 123448 254638 123457
rect 254582 123383 254638 123392
rect 254582 114880 254638 114889
rect 254582 114815 254638 114824
rect 253940 105596 253992 105602
rect 253940 105538 253992 105544
rect 253480 98388 253532 98394
rect 253480 98330 253532 98336
rect 253492 91866 253520 98330
rect 253480 91860 253532 91866
rect 253480 91802 253532 91808
rect 253388 61396 253440 61402
rect 253388 61338 253440 61344
rect 254596 47598 254624 114815
rect 254688 102134 254716 142122
rect 255424 139398 255452 221410
rect 255516 216578 255544 241470
rect 255504 216572 255556 216578
rect 255504 216514 255556 216520
rect 255516 215354 255544 216514
rect 255504 215348 255556 215354
rect 255504 215290 255556 215296
rect 255964 215348 256016 215354
rect 255964 215290 256016 215296
rect 255976 193934 256004 215290
rect 255964 193928 256016 193934
rect 255964 193870 256016 193876
rect 256712 174321 256740 303622
rect 256790 297392 256846 297401
rect 256790 297327 256846 297336
rect 256804 270502 256832 297327
rect 256884 289944 256936 289950
rect 256884 289886 256936 289892
rect 256792 270496 256844 270502
rect 256792 270438 256844 270444
rect 256804 269822 256832 270438
rect 256792 269816 256844 269822
rect 256792 269758 256844 269764
rect 256790 261216 256846 261225
rect 256790 261151 256846 261160
rect 256804 211070 256832 261151
rect 256896 253910 256924 289886
rect 256884 253904 256936 253910
rect 256884 253846 256936 253852
rect 256896 253230 256924 253846
rect 256884 253224 256936 253230
rect 256884 253166 256936 253172
rect 258092 240145 258120 371214
rect 262218 358048 262274 358057
rect 262218 357983 262274 357992
rect 258172 340944 258224 340950
rect 258172 340886 258224 340892
rect 258078 240136 258134 240145
rect 258078 240071 258134 240080
rect 258184 238649 258212 340886
rect 259460 339516 259512 339522
rect 259460 339458 259512 339464
rect 259472 271930 259500 339458
rect 261576 305040 261628 305046
rect 261576 304982 261628 304988
rect 261484 302320 261536 302326
rect 261484 302262 261536 302268
rect 259552 295996 259604 296002
rect 259552 295938 259604 295944
rect 259460 271924 259512 271930
rect 259460 271866 259512 271872
rect 259460 262880 259512 262886
rect 259460 262822 259512 262828
rect 258170 238640 258226 238649
rect 258170 238575 258226 238584
rect 256792 211064 256844 211070
rect 256792 211006 256844 211012
rect 256698 174312 256754 174321
rect 256698 174247 256754 174256
rect 255964 174004 256016 174010
rect 255964 173946 256016 173952
rect 255976 141438 256004 173946
rect 256804 162489 256832 211006
rect 257434 171592 257490 171601
rect 257434 171527 257490 171536
rect 256790 162480 256846 162489
rect 256790 162415 256846 162424
rect 257344 161560 257396 161566
rect 257344 161502 257396 161508
rect 256240 146940 256292 146946
rect 256240 146882 256292 146888
rect 255964 141432 256016 141438
rect 255964 141374 256016 141380
rect 256056 140820 256108 140826
rect 256056 140762 256108 140768
rect 255412 139392 255464 139398
rect 255412 139334 255464 139340
rect 254766 112024 254822 112033
rect 254766 111959 254822 111968
rect 254676 102128 254728 102134
rect 254676 102070 254728 102076
rect 254780 75206 254808 111959
rect 255964 110560 256016 110566
rect 255964 110502 256016 110508
rect 254860 104848 254912 104854
rect 254860 104790 254912 104796
rect 254872 86358 254900 104790
rect 254860 86352 254912 86358
rect 254860 86294 254912 86300
rect 254768 75200 254820 75206
rect 254768 75142 254820 75148
rect 255976 50386 256004 110502
rect 256068 97918 256096 140762
rect 256148 139460 256200 139466
rect 256148 139402 256200 139408
rect 256160 98394 256188 139402
rect 256252 109002 256280 146882
rect 257356 146674 257384 161502
rect 257344 146668 257396 146674
rect 257344 146610 257396 146616
rect 257344 133952 257396 133958
rect 257344 133894 257396 133900
rect 256240 108996 256292 109002
rect 256240 108938 256292 108944
rect 256148 98388 256200 98394
rect 256148 98330 256200 98336
rect 256240 98048 256292 98054
rect 256240 97990 256292 97996
rect 256056 97912 256108 97918
rect 256056 97854 256108 97860
rect 256148 96688 256200 96694
rect 256148 96630 256200 96636
rect 256160 80753 256188 96630
rect 256146 80744 256202 80753
rect 256146 80679 256202 80688
rect 256252 68241 256280 97990
rect 256238 68232 256294 68241
rect 256238 68167 256294 68176
rect 257356 64161 257384 133894
rect 257448 132462 257476 171527
rect 259472 153105 259500 262822
rect 259564 256630 259592 295938
rect 260102 287464 260158 287473
rect 260102 287399 260158 287408
rect 260116 272542 260144 287399
rect 260104 272536 260156 272542
rect 260104 272478 260156 272484
rect 259552 256624 259604 256630
rect 259552 256566 259604 256572
rect 260748 256624 260800 256630
rect 260748 256566 260800 256572
rect 260760 256018 260788 256566
rect 260748 256012 260800 256018
rect 260748 255954 260800 255960
rect 260102 174448 260158 174457
rect 260102 174383 260158 174392
rect 259458 153096 259514 153105
rect 259458 153031 259514 153040
rect 258814 152008 258870 152017
rect 258814 151943 258870 151952
rect 257526 146568 257582 146577
rect 257526 146503 257582 146512
rect 257436 132456 257488 132462
rect 257436 132398 257488 132404
rect 257540 124817 257568 146503
rect 257620 138032 257672 138038
rect 257620 137974 257672 137980
rect 257526 124808 257582 124817
rect 257526 124743 257582 124752
rect 257528 122868 257580 122874
rect 257528 122810 257580 122816
rect 257436 109064 257488 109070
rect 257436 109006 257488 109012
rect 257342 64152 257398 64161
rect 257342 64087 257398 64096
rect 257448 53106 257476 109006
rect 257540 76673 257568 122810
rect 257632 104854 257660 137974
rect 258724 135312 258776 135318
rect 258724 135254 258776 135260
rect 258736 127634 258764 135254
rect 258724 127628 258776 127634
rect 258724 127570 258776 127576
rect 258724 125656 258776 125662
rect 258724 125598 258776 125604
rect 257620 104848 257672 104854
rect 257620 104790 257672 104796
rect 257526 76664 257582 76673
rect 257526 76599 257582 76608
rect 257436 53100 257488 53106
rect 257436 53042 257488 53048
rect 255964 50380 256016 50386
rect 255964 50322 256016 50328
rect 254584 47592 254636 47598
rect 254584 47534 254636 47540
rect 253296 37936 253348 37942
rect 253296 37878 253348 37884
rect 258078 35184 258134 35193
rect 258078 35119 258134 35128
rect 255318 19952 255374 19961
rect 255318 19887 255374 19896
rect 255332 16574 255360 19887
rect 258092 16574 258120 35119
rect 258736 32502 258764 125598
rect 258828 110401 258856 151943
rect 259090 148336 259146 148345
rect 259090 148271 259146 148280
rect 259104 147937 259132 148271
rect 259090 147928 259146 147937
rect 259090 147863 259146 147872
rect 259000 146872 259052 146878
rect 259000 146814 259052 146820
rect 258906 113384 258962 113393
rect 258906 113319 258962 113328
rect 258814 110392 258870 110401
rect 258814 110327 258870 110336
rect 258816 104984 258868 104990
rect 258816 104926 258868 104932
rect 258828 44946 258856 104926
rect 258920 77897 258948 113319
rect 259012 113082 259040 146814
rect 260116 135250 260144 174383
rect 260196 158772 260248 158778
rect 260196 158714 260248 158720
rect 260208 140078 260236 158714
rect 260288 142248 260340 142254
rect 260288 142190 260340 142196
rect 260196 140072 260248 140078
rect 260196 140014 260248 140020
rect 260104 135244 260156 135250
rect 260104 135186 260156 135192
rect 260102 121680 260158 121689
rect 260102 121615 260158 121624
rect 259000 113076 259052 113082
rect 259000 113018 259052 113024
rect 259000 107772 259052 107778
rect 259000 107714 259052 107720
rect 259012 93158 259040 107714
rect 259000 93152 259052 93158
rect 259000 93094 259052 93100
rect 258906 77888 258962 77897
rect 258906 77823 258962 77832
rect 258816 44940 258868 44946
rect 258816 44882 258868 44888
rect 259460 43512 259512 43518
rect 259460 43454 259512 43460
rect 258724 32496 258776 32502
rect 258724 32438 258776 32444
rect 255332 16546 255912 16574
rect 258092 16546 258304 16574
rect 253204 13116 253256 13122
rect 253204 13058 253256 13064
rect 251178 11656 251234 11665
rect 251178 11591 251234 11600
rect 251192 480 251220 11591
rect 253480 7608 253532 7614
rect 253480 7550 253532 7556
rect 252374 3496 252430 3505
rect 252374 3431 252430 3440
rect 252388 480 252416 3431
rect 253492 480 253520 7550
rect 254676 2168 254728 2174
rect 254676 2110 254728 2116
rect 254688 480 254716 2110
rect 255884 480 255912 16546
rect 257068 3528 257120 3534
rect 257068 3470 257120 3476
rect 257080 480 257108 3470
rect 258276 480 258304 16546
rect 259472 11762 259500 43454
rect 260116 40798 260144 121615
rect 260196 104916 260248 104922
rect 260196 104858 260248 104864
rect 260208 49026 260236 104858
rect 260300 101425 260328 142190
rect 260380 139528 260432 139534
rect 260380 139470 260432 139476
rect 260392 106282 260420 139470
rect 260472 111852 260524 111858
rect 260472 111794 260524 111800
rect 260380 106276 260432 106282
rect 260380 106218 260432 106224
rect 260286 101416 260342 101425
rect 260286 101351 260342 101360
rect 260380 100836 260432 100842
rect 260380 100778 260432 100784
rect 260392 83473 260420 100778
rect 260484 89010 260512 111794
rect 261496 93770 261524 302262
rect 261588 242214 261616 304982
rect 262232 252550 262260 357983
rect 320180 353320 320232 353326
rect 320180 353262 320232 353268
rect 263690 349208 263746 349217
rect 263690 349143 263746 349152
rect 262862 285832 262918 285841
rect 262862 285767 262918 285776
rect 262220 252544 262272 252550
rect 262220 252486 262272 252492
rect 262680 252544 262732 252550
rect 262680 252486 262732 252492
rect 262692 251870 262720 252486
rect 262680 251864 262732 251870
rect 262680 251806 262732 251812
rect 261576 242208 261628 242214
rect 261576 242150 261628 242156
rect 262876 203658 262904 285767
rect 263704 266529 263732 349143
rect 304998 335472 305054 335481
rect 304998 335407 305054 335416
rect 300952 317484 301004 317490
rect 300952 317426 301004 317432
rect 282184 311908 282236 311914
rect 282184 311850 282236 311856
rect 267002 310584 267058 310593
rect 267002 310519 267058 310528
rect 265624 298172 265676 298178
rect 265624 298114 265676 298120
rect 264242 284472 264298 284481
rect 264242 284407 264298 284416
rect 263690 266520 263746 266529
rect 263690 266455 263746 266464
rect 263600 266416 263652 266422
rect 263600 266358 263652 266364
rect 263612 224913 263640 266358
rect 263704 265674 263732 266455
rect 263692 265668 263744 265674
rect 263692 265610 263744 265616
rect 264256 259418 264284 284407
rect 264244 259412 264296 259418
rect 264244 259354 264296 259360
rect 265636 250510 265664 298114
rect 265716 261520 265768 261526
rect 265716 261462 265768 261468
rect 265624 250504 265676 250510
rect 265624 250446 265676 250452
rect 265624 242956 265676 242962
rect 265624 242898 265676 242904
rect 263598 224904 263654 224913
rect 263598 224839 263654 224848
rect 263612 224505 263640 224839
rect 263598 224496 263654 224505
rect 263598 224431 263654 224440
rect 264242 224496 264298 224505
rect 264242 224431 264298 224440
rect 262864 203652 262916 203658
rect 262864 203594 262916 203600
rect 264256 202162 264284 224431
rect 264244 202156 264296 202162
rect 264244 202098 264296 202104
rect 265636 182850 265664 242898
rect 265728 237386 265756 261462
rect 265716 237380 265768 237386
rect 265716 237322 265768 237328
rect 267016 194041 267044 310519
rect 273904 307828 273956 307834
rect 273904 307770 273956 307776
rect 271144 306468 271196 306474
rect 271144 306410 271196 306416
rect 269948 300892 270000 300898
rect 269948 300834 270000 300840
rect 268382 295488 268438 295497
rect 268382 295423 268438 295432
rect 267002 194032 267058 194041
rect 267002 193967 267058 193976
rect 268396 192574 268424 295423
rect 269764 285728 269816 285734
rect 269764 285670 269816 285676
rect 268476 193928 268528 193934
rect 268476 193870 268528 193876
rect 268384 192568 268436 192574
rect 268384 192510 268436 192516
rect 265624 182844 265676 182850
rect 265624 182786 265676 182792
rect 268488 177342 268516 193870
rect 269776 181529 269804 285670
rect 269856 250572 269908 250578
rect 269856 250514 269908 250520
rect 269762 181520 269818 181529
rect 269762 181455 269818 181464
rect 269868 180198 269896 250514
rect 269960 242282 269988 300834
rect 269948 242276 270000 242282
rect 269948 242218 270000 242224
rect 271156 185745 271184 306410
rect 272522 305008 272578 305017
rect 272522 304943 272578 304952
rect 271236 257372 271288 257378
rect 271236 257314 271288 257320
rect 271142 185736 271198 185745
rect 271142 185671 271198 185680
rect 269856 180192 269908 180198
rect 269856 180134 269908 180140
rect 271248 178702 271276 257314
rect 271236 178696 271288 178702
rect 271236 178638 271288 178644
rect 272536 177449 272564 304943
rect 273916 181558 273944 307770
rect 278044 294024 278096 294030
rect 278044 293966 278096 293972
rect 273996 280220 274048 280226
rect 273996 280162 274048 280168
rect 273904 181552 273956 181558
rect 273904 181494 273956 181500
rect 272522 177440 272578 177449
rect 274008 177410 274036 280162
rect 276664 259548 276716 259554
rect 276664 259490 276716 259496
rect 276676 184278 276704 259490
rect 276754 216064 276810 216073
rect 276754 215999 276810 216008
rect 276664 184272 276716 184278
rect 276664 184214 276716 184220
rect 276768 178945 276796 215999
rect 278056 179489 278084 293966
rect 280160 288516 280212 288522
rect 280160 288458 280212 288464
rect 278136 276684 278188 276690
rect 278136 276626 278188 276632
rect 278042 179480 278098 179489
rect 278042 179415 278098 179424
rect 276754 178936 276810 178945
rect 276754 178871 276810 178880
rect 272522 177375 272578 177384
rect 273996 177404 274048 177410
rect 273996 177346 274048 177352
rect 268476 177336 268528 177342
rect 268476 177278 268528 177284
rect 278148 176254 278176 276626
rect 279424 258120 279476 258126
rect 279424 258062 279476 258068
rect 278228 242208 278280 242214
rect 278228 242150 278280 242156
rect 278240 178974 278268 242150
rect 279056 195288 279108 195294
rect 279056 195230 279108 195236
rect 278780 180124 278832 180130
rect 278780 180066 278832 180072
rect 278792 179110 278820 180066
rect 278780 179104 278832 179110
rect 278780 179046 278832 179052
rect 278228 178968 278280 178974
rect 278228 178910 278280 178916
rect 278780 178968 278832 178974
rect 278780 178910 278832 178916
rect 278792 177041 278820 178910
rect 278778 177032 278834 177041
rect 278778 176967 278834 176976
rect 278136 176248 278188 176254
rect 278136 176190 278188 176196
rect 264978 175672 265034 175681
rect 264978 175607 265034 175616
rect 264992 175370 265020 175607
rect 264980 175364 265032 175370
rect 264980 175306 265032 175312
rect 265070 175264 265126 175273
rect 265070 175199 265126 175208
rect 264978 174856 265034 174865
rect 264978 174791 265034 174800
rect 264992 174010 265020 174791
rect 264980 174004 265032 174010
rect 264980 173946 265032 173952
rect 265084 173942 265112 175199
rect 265072 173936 265124 173942
rect 265072 173878 265124 173884
rect 265070 173632 265126 173641
rect 265070 173567 265126 173576
rect 264978 172680 265034 172689
rect 264978 172615 264980 172624
rect 265032 172615 265034 172624
rect 264980 172586 265032 172592
rect 265084 172582 265112 173567
rect 265072 172576 265124 172582
rect 265072 172518 265124 172524
rect 265070 172272 265126 172281
rect 265070 172207 265126 172216
rect 264978 171456 265034 171465
rect 264978 171391 265034 171400
rect 264992 171222 265020 171391
rect 264980 171216 265032 171222
rect 264980 171158 265032 171164
rect 265084 171154 265112 172207
rect 265072 171148 265124 171154
rect 265072 171090 265124 171096
rect 265070 171048 265126 171057
rect 265070 170983 265126 170992
rect 264978 170096 265034 170105
rect 264978 170031 265034 170040
rect 264992 169862 265020 170031
rect 264980 169856 265032 169862
rect 264980 169798 265032 169804
rect 265084 169794 265112 170983
rect 265072 169788 265124 169794
rect 265072 169730 265124 169736
rect 264978 169688 265034 169697
rect 264978 169623 265034 169632
rect 264242 169280 264298 169289
rect 264242 169215 264298 169224
rect 261758 164520 261814 164529
rect 261758 164455 261814 164464
rect 261668 140888 261720 140894
rect 261668 140830 261720 140836
rect 261576 131232 261628 131238
rect 261576 131174 261628 131180
rect 261484 93764 261536 93770
rect 261484 93706 261536 93712
rect 260472 89004 260524 89010
rect 260472 88946 260524 88952
rect 260378 83464 260434 83473
rect 260378 83399 260434 83408
rect 261588 54505 261616 131174
rect 261680 100706 261708 140830
rect 261772 124166 261800 164455
rect 263046 162888 263102 162897
rect 263046 162823 263102 162832
rect 262862 138272 262918 138281
rect 262862 138207 262918 138216
rect 261760 124160 261812 124166
rect 261760 124102 261812 124108
rect 262128 123072 262180 123078
rect 262128 123014 262180 123020
rect 262140 120737 262168 123014
rect 262126 120728 262182 120737
rect 262126 120663 262182 120672
rect 262310 119504 262366 119513
rect 262310 119439 262366 119448
rect 262324 119105 262352 119439
rect 262310 119096 262366 119105
rect 262310 119031 262366 119040
rect 262218 116920 262274 116929
rect 262218 116855 262274 116864
rect 262232 116113 262260 116855
rect 262218 116104 262274 116113
rect 262218 116039 262274 116048
rect 262770 108352 262826 108361
rect 262770 108287 262826 108296
rect 262784 107953 262812 108287
rect 262770 107944 262826 107953
rect 262770 107879 262826 107888
rect 261758 100872 261814 100881
rect 261758 100807 261814 100816
rect 261668 100700 261720 100706
rect 261668 100642 261720 100648
rect 261772 73953 261800 100807
rect 262678 96384 262734 96393
rect 262678 96319 262734 96328
rect 262692 95266 262720 96319
rect 262680 95260 262732 95266
rect 262680 95202 262732 95208
rect 261758 73944 261814 73953
rect 261758 73879 261814 73888
rect 262218 69728 262274 69737
rect 262218 69663 262274 69672
rect 261574 54496 261630 54505
rect 261574 54431 261630 54440
rect 260196 49020 260248 49026
rect 260196 48962 260248 48968
rect 260104 40792 260156 40798
rect 260104 40734 260156 40740
rect 262232 16574 262260 69663
rect 262876 24138 262904 138207
rect 262954 135688 263010 135697
rect 262954 135623 263010 135632
rect 262968 58585 262996 135623
rect 263060 122806 263088 162823
rect 263140 147756 263192 147762
rect 263140 147698 263192 147704
rect 263048 122800 263100 122806
rect 263048 122742 263100 122748
rect 263152 115938 263180 147698
rect 264256 129742 264284 169215
rect 264992 168434 265020 169623
rect 265162 168872 265218 168881
rect 265162 168807 265218 168816
rect 264980 168428 265032 168434
rect 264980 168370 265032 168376
rect 264978 167920 265034 167929
rect 264978 167855 265034 167864
rect 264992 167142 265020 167855
rect 265070 167512 265126 167521
rect 265070 167447 265126 167456
rect 264980 167136 265032 167142
rect 264980 167078 265032 167084
rect 265084 167074 265112 167447
rect 265072 167068 265124 167074
rect 265072 167010 265124 167016
rect 265070 166696 265126 166705
rect 265070 166631 265126 166640
rect 264978 166288 265034 166297
rect 264978 166223 265034 166232
rect 264992 165714 265020 166223
rect 264980 165708 265032 165714
rect 264980 165650 265032 165656
rect 265084 165646 265112 166631
rect 265072 165640 265124 165646
rect 265072 165582 265124 165588
rect 264978 165336 265034 165345
rect 264978 165271 265034 165280
rect 264992 164286 265020 165271
rect 265176 164898 265204 168807
rect 265164 164892 265216 164898
rect 265164 164834 265216 164840
rect 267830 164656 267886 164665
rect 267830 164591 267886 164600
rect 267844 164393 267872 164591
rect 265622 164384 265678 164393
rect 265622 164319 265678 164328
rect 267830 164384 267886 164393
rect 267830 164319 267886 164328
rect 264980 164280 265032 164286
rect 264980 164222 265032 164228
rect 265070 164112 265126 164121
rect 265070 164047 265126 164056
rect 264978 163704 265034 163713
rect 264978 163639 265034 163648
rect 264992 162994 265020 163639
rect 264980 162988 265032 162994
rect 264980 162930 265032 162936
rect 265084 162926 265112 164047
rect 265072 162920 265124 162926
rect 265072 162862 265124 162868
rect 265162 162344 265218 162353
rect 265162 162279 265218 162288
rect 265070 161936 265126 161945
rect 265070 161871 265126 161880
rect 264980 161560 265032 161566
rect 264978 161528 264980 161537
rect 265032 161528 265034 161537
rect 265084 161498 265112 161871
rect 264978 161463 265034 161472
rect 265072 161492 265124 161498
rect 265072 161434 265124 161440
rect 265070 161120 265126 161129
rect 265070 161055 265126 161064
rect 264978 160304 265034 160313
rect 264978 160239 265034 160248
rect 264992 160206 265020 160239
rect 264980 160200 265032 160206
rect 264980 160142 265032 160148
rect 265084 160138 265112 161055
rect 265072 160132 265124 160138
rect 265072 160074 265124 160080
rect 265070 159760 265126 159769
rect 265070 159695 265126 159704
rect 264978 158944 265034 158953
rect 264978 158879 265034 158888
rect 264992 158778 265020 158879
rect 264980 158772 265032 158778
rect 264980 158714 265032 158720
rect 264978 158536 265034 158545
rect 264978 158471 265034 158480
rect 264992 157418 265020 158471
rect 265084 158030 265112 159695
rect 265176 159390 265204 162279
rect 265164 159384 265216 159390
rect 265164 159326 265216 159332
rect 265162 158128 265218 158137
rect 265162 158063 265218 158072
rect 265072 158024 265124 158030
rect 265072 157966 265124 157972
rect 264980 157412 265032 157418
rect 264980 157354 265032 157360
rect 265070 157176 265126 157185
rect 265070 157111 265126 157120
rect 264978 156768 265034 156777
rect 264978 156703 265034 156712
rect 264992 156058 265020 156703
rect 264980 156052 265032 156058
rect 264980 155994 265032 156000
rect 265084 155990 265112 157111
rect 265176 156641 265204 158063
rect 265162 156632 265218 156641
rect 265162 156567 265218 156576
rect 265072 155984 265124 155990
rect 265072 155926 265124 155932
rect 265162 155952 265218 155961
rect 265162 155887 265218 155896
rect 264980 154692 265032 154698
rect 264980 154634 265032 154640
rect 264992 154601 265020 154634
rect 265176 154630 265204 155887
rect 265164 154624 265216 154630
rect 264978 154592 265034 154601
rect 265164 154566 265216 154572
rect 264978 154527 265034 154536
rect 265636 153882 265664 164319
rect 265714 156360 265770 156369
rect 265714 156295 265770 156304
rect 265624 153876 265676 153882
rect 265624 153818 265676 153824
rect 265254 153776 265310 153785
rect 265254 153711 265310 153720
rect 264520 153468 264572 153474
rect 264520 153410 264572 153416
rect 264532 151814 264560 153410
rect 265070 152960 265126 152969
rect 265070 152895 265126 152904
rect 264978 152552 265034 152561
rect 264978 152487 265034 152496
rect 264992 151910 265020 152487
rect 264980 151904 265032 151910
rect 264980 151846 265032 151852
rect 265084 151842 265112 152895
rect 264440 151786 264560 151814
rect 265072 151836 265124 151842
rect 264244 129736 264296 129742
rect 264244 129678 264296 129684
rect 264242 118960 264298 118969
rect 264242 118895 264298 118904
rect 263232 116068 263284 116074
rect 263232 116010 263284 116016
rect 263140 115932 263192 115938
rect 263140 115874 263192 115880
rect 263046 102640 263102 102649
rect 263046 102575 263102 102584
rect 263060 82113 263088 102575
rect 263244 97889 263272 116010
rect 263230 97880 263286 97889
rect 263230 97815 263286 97824
rect 263140 96756 263192 96762
rect 263140 96698 263192 96704
rect 263152 89049 263180 96698
rect 263138 89040 263194 89049
rect 263138 88975 263194 88984
rect 263046 82104 263102 82113
rect 263046 82039 263102 82048
rect 262954 58576 263010 58585
rect 262954 58511 263010 58520
rect 263598 30968 263654 30977
rect 263598 30903 263654 30912
rect 262864 24132 262916 24138
rect 262864 24074 262916 24080
rect 263612 16574 263640 30903
rect 262232 16546 262536 16574
rect 263612 16546 264192 16574
rect 261758 13016 261814 13025
rect 261758 12951 261814 12960
rect 259460 11756 259512 11762
rect 259460 11698 259512 11704
rect 260656 11756 260708 11762
rect 260656 11698 260708 11704
rect 259458 10296 259514 10305
rect 259458 10231 259514 10240
rect 259472 480 259500 10231
rect 260668 480 260696 11698
rect 261772 480 261800 12951
rect 262508 490 262536 16546
rect 262784 598 262996 626
rect 262784 490 262812 598
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 462 262812 490
rect 262968 480 262996 598
rect 264164 480 264192 16546
rect 264256 8974 264284 118895
rect 264336 118040 264388 118046
rect 264336 117982 264388 117988
rect 264348 80889 264376 117982
rect 264440 114481 264468 151786
rect 265072 151778 265124 151784
rect 264978 151600 265034 151609
rect 264978 151535 265034 151544
rect 264520 150544 264572 150550
rect 264520 150486 264572 150492
rect 264426 114472 264482 114481
rect 264426 114407 264482 114416
rect 264532 113150 264560 150486
rect 264992 150482 265020 151535
rect 265070 151192 265126 151201
rect 265070 151127 265126 151136
rect 264980 150476 265032 150482
rect 264980 150418 265032 150424
rect 264978 150376 265034 150385
rect 264978 150311 265034 150320
rect 264992 149122 265020 150311
rect 265084 149734 265112 151127
rect 265162 149968 265218 149977
rect 265162 149903 265218 149912
rect 265072 149728 265124 149734
rect 265072 149670 265124 149676
rect 264980 149116 265032 149122
rect 264980 149058 265032 149064
rect 264978 149016 265034 149025
rect 264978 148951 265034 148960
rect 264992 147694 265020 148951
rect 264980 147688 265032 147694
rect 264980 147630 265032 147636
rect 265176 146946 265204 149903
rect 265164 146940 265216 146946
rect 265164 146882 265216 146888
rect 265268 146878 265296 153711
rect 265622 148608 265678 148617
rect 265622 148543 265678 148552
rect 265256 146872 265308 146878
rect 265256 146814 265308 146820
rect 265162 146432 265218 146441
rect 265162 146367 265218 146376
rect 265070 146024 265126 146033
rect 265070 145959 265126 145968
rect 264978 145208 265034 145217
rect 264978 145143 265034 145152
rect 264992 144974 265020 145143
rect 265084 145042 265112 145959
rect 265072 145036 265124 145042
rect 265072 144978 265124 144984
rect 264980 144968 265032 144974
rect 264980 144910 265032 144916
rect 264978 144800 265034 144809
rect 264978 144735 265034 144744
rect 264992 143614 265020 144735
rect 265176 144226 265204 146367
rect 265164 144220 265216 144226
rect 265164 144162 265216 144168
rect 265254 143848 265310 143857
rect 265254 143783 265310 143792
rect 264980 143608 265032 143614
rect 264980 143550 265032 143556
rect 264978 143440 265034 143449
rect 264978 143375 265034 143384
rect 264992 142186 265020 143375
rect 265162 143032 265218 143041
rect 265162 142967 265218 142976
rect 265072 142248 265124 142254
rect 265070 142216 265072 142225
rect 265124 142216 265126 142225
rect 264980 142180 265032 142186
rect 265070 142151 265126 142160
rect 264980 142122 265032 142128
rect 265176 140894 265204 142967
rect 265164 140888 265216 140894
rect 264978 140856 265034 140865
rect 265164 140830 265216 140836
rect 264978 140791 264980 140800
rect 265032 140791 265034 140800
rect 264980 140762 265032 140768
rect 264978 139632 265034 139641
rect 264978 139567 265034 139576
rect 264992 139466 265020 139567
rect 264980 139460 265032 139466
rect 264980 139402 265032 139408
rect 264978 138680 265034 138689
rect 264978 138615 265034 138624
rect 264992 138038 265020 138615
rect 264980 138032 265032 138038
rect 264980 137974 265032 137980
rect 264978 137456 265034 137465
rect 264978 137391 265034 137400
rect 264992 136678 265020 137391
rect 264980 136672 265032 136678
rect 264980 136614 265032 136620
rect 265070 136640 265126 136649
rect 265070 136575 265126 136584
rect 265084 135318 265112 136575
rect 265268 135930 265296 143783
rect 265346 141808 265402 141817
rect 265346 141743 265402 141752
rect 265256 135924 265308 135930
rect 265256 135866 265308 135872
rect 265072 135312 265124 135318
rect 265072 135254 265124 135260
rect 265360 134473 265388 141743
rect 265636 138718 265664 148543
rect 265728 147762 265756 156295
rect 265806 155544 265862 155553
rect 265806 155479 265862 155488
rect 265820 153474 265848 155479
rect 266266 154184 266322 154193
rect 266266 154119 266322 154128
rect 265808 153468 265860 153474
rect 265808 153410 265860 153416
rect 266280 150550 266308 154119
rect 279068 151814 279096 195230
rect 279146 188592 279202 188601
rect 279146 188527 279202 188536
rect 279160 161474 279188 188527
rect 279436 180266 279464 258062
rect 279424 180260 279476 180266
rect 279424 180202 279476 180208
rect 279422 179072 279478 179081
rect 279422 179007 279478 179016
rect 279238 176760 279294 176769
rect 279238 176695 279294 176704
rect 279252 166994 279280 176695
rect 279332 175432 279384 175438
rect 279332 175374 279384 175380
rect 279344 175273 279372 175374
rect 279330 175264 279386 175273
rect 279330 175199 279386 175208
rect 279436 174457 279464 179007
rect 279422 174448 279478 174457
rect 279422 174383 279478 174392
rect 279252 166966 279372 166994
rect 279344 165889 279372 166966
rect 279330 165880 279386 165889
rect 279330 165815 279386 165824
rect 279160 161446 279464 161474
rect 279068 151786 279372 151814
rect 279344 150657 279372 151786
rect 279330 150648 279386 150657
rect 279330 150583 279386 150592
rect 266268 150544 266320 150550
rect 266268 150486 266320 150492
rect 265716 147756 265768 147762
rect 265716 147698 265768 147704
rect 265898 147384 265954 147393
rect 265898 147319 265954 147328
rect 265806 140040 265862 140049
rect 265806 139975 265862 139984
rect 265624 138712 265676 138718
rect 265624 138654 265676 138660
rect 265346 134464 265402 134473
rect 265346 134399 265402 134408
rect 265622 134464 265678 134473
rect 265622 134399 265678 134408
rect 264978 134056 265034 134065
rect 264978 133991 265034 134000
rect 264992 133958 265020 133991
rect 264980 133952 265032 133958
rect 264980 133894 265032 133900
rect 265070 133648 265126 133657
rect 265070 133583 265126 133592
rect 264978 133104 265034 133113
rect 264978 133039 265034 133048
rect 264992 132598 265020 133039
rect 264980 132592 265032 132598
rect 264980 132534 265032 132540
rect 265084 132530 265112 133583
rect 265072 132524 265124 132530
rect 265072 132466 265124 132472
rect 264978 131880 265034 131889
rect 264978 131815 265034 131824
rect 264992 131170 265020 131815
rect 265070 131472 265126 131481
rect 265070 131407 265126 131416
rect 265084 131238 265112 131407
rect 265072 131232 265124 131238
rect 265072 131174 265124 131180
rect 264980 131164 265032 131170
rect 264980 131106 265032 131112
rect 264978 130520 265034 130529
rect 264978 130455 265034 130464
rect 264992 129810 265020 130455
rect 264980 129804 265032 129810
rect 264980 129746 265032 129752
rect 264978 129704 265034 129713
rect 264978 129639 265034 129648
rect 264992 128382 265020 129639
rect 264980 128376 265032 128382
rect 264980 128318 265032 128324
rect 264978 127528 265034 127537
rect 264978 127463 265034 127472
rect 264992 127022 265020 127463
rect 264980 127016 265032 127022
rect 264980 126958 265032 126964
rect 264978 126304 265034 126313
rect 264978 126239 265034 126248
rect 264992 125662 265020 126239
rect 264980 125656 265032 125662
rect 264980 125598 265032 125604
rect 264610 125352 264666 125361
rect 264610 125287 264666 125296
rect 264624 118046 264652 125287
rect 264978 124944 265034 124953
rect 264978 124879 265034 124888
rect 264992 124234 265020 124879
rect 264980 124228 265032 124234
rect 264980 124170 265032 124176
rect 264978 124128 265034 124137
rect 264978 124063 265034 124072
rect 264992 122874 265020 124063
rect 265070 123312 265126 123321
rect 265070 123247 265126 123256
rect 265084 123078 265112 123247
rect 265072 123072 265124 123078
rect 265072 123014 265124 123020
rect 264980 122868 265032 122874
rect 264980 122810 265032 122816
rect 264978 122360 265034 122369
rect 264978 122295 265034 122304
rect 264992 121514 265020 122295
rect 264980 121508 265032 121514
rect 264980 121450 265032 121456
rect 264978 121136 265034 121145
rect 264978 121071 265034 121080
rect 264992 120154 265020 121071
rect 264980 120148 265032 120154
rect 264980 120090 265032 120096
rect 265070 118552 265126 118561
rect 265070 118487 265126 118496
rect 264978 118144 265034 118153
rect 264978 118079 265034 118088
rect 264612 118040 264664 118046
rect 264612 117982 264664 117988
rect 264992 117366 265020 118079
rect 265084 117434 265112 118487
rect 265072 117428 265124 117434
rect 265072 117370 265124 117376
rect 264980 117360 265032 117366
rect 264980 117302 265032 117308
rect 264978 117192 265034 117201
rect 264978 117127 265034 117136
rect 264992 116006 265020 117127
rect 265070 116376 265126 116385
rect 265070 116311 265126 116320
rect 265084 116074 265112 116311
rect 265072 116068 265124 116074
rect 265072 116010 265124 116016
rect 264980 116000 265032 116006
rect 264980 115942 265032 115948
rect 264978 115560 265034 115569
rect 264978 115495 265034 115504
rect 264992 114578 265020 115495
rect 264980 114572 265032 114578
rect 264980 114514 265032 114520
rect 265070 114200 265126 114209
rect 265070 114135 265126 114144
rect 264978 113792 265034 113801
rect 264978 113727 265034 113736
rect 264992 113218 265020 113727
rect 265084 113286 265112 114135
rect 265072 113280 265124 113286
rect 265072 113222 265124 113228
rect 264980 113212 265032 113218
rect 264980 113154 265032 113160
rect 264520 113144 264572 113150
rect 264520 113086 264572 113092
rect 264978 112568 265034 112577
rect 264978 112503 265034 112512
rect 264992 111858 265020 112503
rect 264980 111852 265032 111858
rect 264980 111794 265032 111800
rect 265070 111616 265126 111625
rect 265070 111551 265126 111560
rect 264978 111208 265034 111217
rect 264978 111143 265034 111152
rect 264992 110566 265020 111143
rect 264980 110560 265032 110566
rect 264980 110502 265032 110508
rect 265084 110498 265112 111551
rect 265072 110492 265124 110498
rect 265072 110434 265124 110440
rect 264426 110392 264482 110401
rect 264426 110327 264482 110336
rect 264334 80880 264390 80889
rect 264334 80815 264390 80824
rect 264440 71233 264468 110327
rect 264978 109984 265034 109993
rect 264978 109919 265034 109928
rect 264992 109070 265020 109919
rect 264980 109064 265032 109070
rect 264980 109006 265032 109012
rect 265070 109032 265126 109041
rect 265070 108967 265126 108976
rect 264978 107808 265034 107817
rect 264978 107743 264980 107752
rect 265032 107743 265034 107752
rect 264980 107714 265032 107720
rect 265084 107710 265112 108967
rect 265072 107704 265124 107710
rect 265072 107646 265124 107652
rect 265070 107400 265126 107409
rect 265070 107335 265126 107344
rect 264978 106992 265034 107001
rect 264978 106927 265034 106936
rect 264992 106418 265020 106927
rect 264980 106412 265032 106418
rect 264980 106354 265032 106360
rect 265084 106350 265112 107335
rect 265072 106344 265124 106350
rect 265072 106286 265124 106292
rect 264978 106040 265034 106049
rect 264978 105975 265034 105984
rect 264992 104922 265020 105975
rect 265070 105632 265126 105641
rect 265070 105567 265126 105576
rect 265084 104990 265112 105567
rect 265072 104984 265124 104990
rect 265072 104926 265124 104932
rect 264980 104916 265032 104922
rect 264980 104858 265032 104864
rect 264978 104816 265034 104825
rect 264978 104751 265034 104760
rect 264992 103562 265020 104751
rect 264980 103556 265032 103562
rect 264980 103498 265032 103504
rect 264978 103456 265034 103465
rect 264978 103391 265034 103400
rect 264794 103048 264850 103057
rect 264794 102983 264850 102992
rect 264808 98705 264836 102983
rect 264992 102202 265020 103391
rect 264980 102196 265032 102202
rect 264980 102138 265032 102144
rect 264978 101824 265034 101833
rect 264978 101759 265034 101768
rect 264992 100774 265020 101759
rect 265070 101280 265126 101289
rect 265070 101215 265126 101224
rect 265084 100842 265112 101215
rect 265072 100836 265124 100842
rect 265072 100778 265124 100784
rect 264980 100768 265032 100774
rect 264980 100710 265032 100716
rect 264978 99648 265034 99657
rect 264978 99583 265034 99592
rect 264992 99414 265020 99583
rect 264980 99408 265032 99414
rect 264980 99350 265032 99356
rect 264794 98696 264850 98705
rect 264794 98631 264850 98640
rect 264978 98696 265034 98705
rect 264978 98631 265034 98640
rect 264992 98054 265020 98631
rect 264980 98048 265032 98054
rect 264980 97990 265032 97996
rect 264978 97472 265034 97481
rect 264978 97407 265034 97416
rect 264992 96694 265020 97407
rect 265072 96756 265124 96762
rect 265072 96698 265124 96704
rect 264980 96688 265032 96694
rect 265084 96665 265112 96698
rect 264980 96630 265032 96636
rect 265070 96656 265126 96665
rect 265070 96591 265126 96600
rect 264426 71224 264482 71233
rect 264426 71159 264482 71168
rect 265636 61441 265664 134399
rect 265714 125896 265770 125905
rect 265714 125831 265770 125840
rect 265728 76566 265756 125831
rect 265820 91798 265848 139975
rect 265912 139534 265940 147319
rect 279436 147121 279464 161446
rect 279422 147112 279478 147121
rect 279422 147047 279478 147056
rect 280172 145897 280200 288458
rect 281908 284436 281960 284442
rect 281908 284378 281960 284384
rect 280252 206304 280304 206310
rect 280252 206246 280304 206252
rect 280158 145888 280214 145897
rect 280158 145823 280214 145832
rect 265900 139528 265952 139534
rect 265900 139470 265952 139476
rect 267094 136232 267150 136241
rect 267094 136167 267150 136176
rect 265898 135280 265954 135289
rect 265898 135215 265954 135224
rect 265912 126342 265940 135215
rect 265900 126336 265952 126342
rect 265900 126278 265952 126284
rect 267002 122904 267058 122913
rect 267002 122839 267058 122848
rect 265898 97064 265954 97073
rect 265898 96999 265954 97008
rect 265808 91792 265860 91798
rect 265808 91734 265860 91740
rect 265912 79393 265940 96999
rect 265898 79384 265954 79393
rect 265898 79319 265954 79328
rect 265716 76560 265768 76566
rect 265716 76502 265768 76508
rect 265622 61432 265678 61441
rect 265622 61367 265678 61376
rect 264978 28248 265034 28257
rect 264978 28183 265034 28192
rect 264244 8968 264296 8974
rect 264244 8910 264296 8916
rect 264992 490 265020 28183
rect 267016 4894 267044 122839
rect 267108 62830 267136 136167
rect 267278 120728 267334 120737
rect 267278 120663 267334 120672
rect 267186 105224 267242 105233
rect 267186 105159 267242 105168
rect 267096 62824 267148 62830
rect 267096 62766 267148 62772
rect 267200 33862 267228 105159
rect 267292 90370 267320 120663
rect 280264 117609 280292 206246
rect 281816 191140 281868 191146
rect 281816 191082 281868 191088
rect 281632 182844 281684 182850
rect 281632 182786 281684 182792
rect 280434 179480 280490 179489
rect 280434 179415 280490 179424
rect 280344 179104 280396 179110
rect 280344 179046 280396 179052
rect 280356 174729 280384 179046
rect 280342 174720 280398 174729
rect 280342 174655 280398 174664
rect 280448 170241 280476 179415
rect 281540 172508 281592 172514
rect 281540 172450 281592 172456
rect 281552 171737 281580 172450
rect 281538 171728 281594 171737
rect 281538 171663 281594 171672
rect 280434 170232 280490 170241
rect 280434 170167 280490 170176
rect 281540 169652 281592 169658
rect 281540 169594 281592 169600
rect 281552 169425 281580 169594
rect 281538 169416 281594 169425
rect 281538 169351 281594 169360
rect 281644 151881 281672 182786
rect 281722 181384 281778 181393
rect 281722 181319 281778 181328
rect 281736 152697 281764 181319
rect 281828 168745 281856 191082
rect 281814 168736 281870 168745
rect 281814 168671 281870 168680
rect 281920 157321 281948 284378
rect 282196 227050 282224 311850
rect 287336 305108 287388 305114
rect 287336 305050 287388 305056
rect 282920 283892 282972 283898
rect 282920 283834 282972 283840
rect 282184 227044 282236 227050
rect 282184 226986 282236 226992
rect 282274 226944 282330 226953
rect 282274 226879 282330 226888
rect 282182 202328 282238 202337
rect 282182 202263 282238 202272
rect 282196 182850 282224 202263
rect 282288 182918 282316 226879
rect 282276 182912 282328 182918
rect 282276 182854 282328 182860
rect 282184 182844 282236 182850
rect 282184 182786 282236 182792
rect 282826 172544 282882 172553
rect 282932 172530 282960 283834
rect 285680 242276 285732 242282
rect 285680 242218 285732 242224
rect 284300 235272 284352 235278
rect 284300 235214 284352 235220
rect 283010 218104 283066 218113
rect 283010 218039 283066 218048
rect 282882 172502 282960 172530
rect 282826 172479 282882 172488
rect 282828 166456 282880 166462
rect 282826 166424 282828 166433
rect 282880 166424 282882 166433
rect 282826 166359 282882 166368
rect 282828 165572 282880 165578
rect 282828 165514 282880 165520
rect 282840 164937 282868 165514
rect 282826 164928 282882 164937
rect 282826 164863 282882 164872
rect 282828 164212 282880 164218
rect 282828 164154 282880 164160
rect 282840 164121 282868 164154
rect 282826 164112 282882 164121
rect 282826 164047 282882 164056
rect 282826 163296 282882 163305
rect 282826 163231 282882 163240
rect 282840 163198 282868 163231
rect 282828 163192 282880 163198
rect 282828 163134 282880 163140
rect 282736 162852 282788 162858
rect 282736 162794 282788 162800
rect 282748 161809 282776 162794
rect 282828 162784 282880 162790
rect 282828 162726 282880 162732
rect 282840 162625 282868 162726
rect 282826 162616 282882 162625
rect 282826 162551 282882 162560
rect 282734 161800 282790 161809
rect 282734 161735 282790 161744
rect 282736 161424 282788 161430
rect 282736 161366 282788 161372
rect 282748 160313 282776 161366
rect 282828 161356 282880 161362
rect 282828 161298 282880 161304
rect 282840 161129 282868 161298
rect 282826 161120 282882 161129
rect 282826 161055 282882 161064
rect 282734 160304 282790 160313
rect 282734 160239 282790 160248
rect 282460 160064 282512 160070
rect 282460 160006 282512 160012
rect 282472 158817 282500 160006
rect 282552 159792 282604 159798
rect 282552 159734 282604 159740
rect 282564 159497 282592 159734
rect 282550 159488 282606 159497
rect 282550 159423 282606 159432
rect 282458 158808 282514 158817
rect 282458 158743 282514 158752
rect 282092 158704 282144 158710
rect 282092 158646 282144 158652
rect 282104 158001 282132 158646
rect 282276 158024 282328 158030
rect 282090 157992 282146 158001
rect 282276 157966 282328 157972
rect 282090 157927 282146 157936
rect 281906 157312 281962 157321
rect 281906 157247 281962 157256
rect 282184 155916 282236 155922
rect 282184 155858 282236 155864
rect 282196 155009 282224 155858
rect 282182 155000 282238 155009
rect 282182 154935 282238 154944
rect 282092 154488 282144 154494
rect 282092 154430 282144 154436
rect 282104 154193 282132 154430
rect 282090 154184 282146 154193
rect 282090 154119 282146 154128
rect 281722 152688 281778 152697
rect 281722 152623 281778 152632
rect 281630 151872 281686 151881
rect 281630 151807 281686 151816
rect 281540 148912 281592 148918
rect 281538 148880 281540 148889
rect 281592 148880 281594 148889
rect 281538 148815 281594 148824
rect 282288 145081 282316 157966
rect 282828 155848 282880 155854
rect 282828 155790 282880 155796
rect 282840 155689 282868 155790
rect 282826 155680 282882 155689
rect 282826 155615 282882 155624
rect 282368 154556 282420 154562
rect 282368 154498 282420 154504
rect 282380 153513 282408 154498
rect 282366 153504 282422 153513
rect 282366 153439 282422 153448
rect 282828 151768 282880 151774
rect 282828 151710 282880 151716
rect 282840 151201 282868 151710
rect 282826 151192 282882 151201
rect 282826 151127 282882 151136
rect 282828 148980 282880 148986
rect 282828 148922 282880 148928
rect 282840 148073 282868 148922
rect 282826 148064 282882 148073
rect 282826 147999 282882 148008
rect 282828 147620 282880 147626
rect 282828 147562 282880 147568
rect 282840 147393 282868 147562
rect 282826 147384 282882 147393
rect 282826 147319 282882 147328
rect 282274 145072 282330 145081
rect 282274 145007 282330 145016
rect 282460 144900 282512 144906
rect 282460 144842 282512 144848
rect 281908 144832 281960 144838
rect 281908 144774 281960 144780
rect 281920 144265 281948 144774
rect 281906 144256 281962 144265
rect 281906 144191 281962 144200
rect 282472 143585 282500 144842
rect 282458 143576 282514 143585
rect 282092 143540 282144 143546
rect 282458 143511 282514 143520
rect 282092 143482 282144 143488
rect 282104 142769 282132 143482
rect 282090 142760 282146 142769
rect 282090 142695 282146 142704
rect 283024 142154 283052 218039
rect 283102 180160 283158 180169
rect 283102 180095 283158 180104
rect 282932 142126 283052 142154
rect 281908 142112 281960 142118
rect 281906 142080 281908 142089
rect 281960 142080 281962 142089
rect 281906 142015 281962 142024
rect 282276 141364 282328 141370
rect 282276 141306 282328 141312
rect 282288 141273 282316 141306
rect 282274 141264 282330 141273
rect 282274 141199 282330 141208
rect 282276 140752 282328 140758
rect 282276 140694 282328 140700
rect 281724 140684 281776 140690
rect 281724 140626 281776 140632
rect 281736 140457 281764 140626
rect 281722 140448 281778 140457
rect 281722 140383 281778 140392
rect 282288 139777 282316 140694
rect 282274 139768 282330 139777
rect 282274 139703 282330 139712
rect 282276 139392 282328 139398
rect 282276 139334 282328 139340
rect 282288 138961 282316 139334
rect 282828 139324 282880 139330
rect 282828 139266 282880 139272
rect 282274 138952 282330 138961
rect 282274 138887 282330 138896
rect 282840 138281 282868 139266
rect 282826 138272 282882 138281
rect 282826 138207 282882 138216
rect 281724 137964 281776 137970
rect 281724 137906 281776 137912
rect 281736 137465 281764 137906
rect 281722 137456 281778 137465
rect 281722 137391 281778 137400
rect 282826 136640 282882 136649
rect 282932 136626 282960 142126
rect 282882 136598 282960 136626
rect 282826 136575 282882 136584
rect 281908 136536 281960 136542
rect 281908 136478 281960 136484
rect 281920 135969 281948 136478
rect 281906 135960 281962 135969
rect 281906 135895 281962 135904
rect 282092 135244 282144 135250
rect 282092 135186 282144 135192
rect 282104 134473 282132 135186
rect 282090 134464 282146 134473
rect 282090 134399 282146 134408
rect 282276 133884 282328 133890
rect 282276 133826 282328 133832
rect 282288 132841 282316 133826
rect 282828 133816 282880 133822
rect 282828 133758 282880 133764
rect 282840 133657 282868 133758
rect 282826 133648 282882 133657
rect 282826 133583 282882 133592
rect 282274 132832 282330 132841
rect 282274 132767 282330 132776
rect 282736 132456 282788 132462
rect 282736 132398 282788 132404
rect 282748 131345 282776 132398
rect 282828 132388 282880 132394
rect 282828 132330 282880 132336
rect 282840 132161 282868 132330
rect 282826 132152 282882 132161
rect 282826 132087 282882 132096
rect 282734 131336 282790 131345
rect 282734 131271 282790 131280
rect 282276 131096 282328 131102
rect 282276 131038 282328 131044
rect 282288 130665 282316 131038
rect 282274 130656 282330 130665
rect 281540 130620 281592 130626
rect 282274 130591 282330 130600
rect 281540 130562 281592 130568
rect 281552 129849 281580 130562
rect 281538 129840 281594 129849
rect 281538 129775 281594 129784
rect 282092 129736 282144 129742
rect 282092 129678 282144 129684
rect 282104 129033 282132 129678
rect 282090 129024 282146 129033
rect 282090 128959 282146 128968
rect 282826 128344 282882 128353
rect 282826 128279 282828 128288
rect 282880 128279 282882 128288
rect 282828 128250 282880 128256
rect 282736 128240 282788 128246
rect 282736 128182 282788 128188
rect 282748 127537 282776 128182
rect 282734 127528 282790 127537
rect 282734 127463 282790 127472
rect 282276 126948 282328 126954
rect 282276 126890 282328 126896
rect 282288 126041 282316 126890
rect 282274 126032 282330 126041
rect 282274 125967 282330 125976
rect 282828 125588 282880 125594
rect 282828 125530 282880 125536
rect 282092 125520 282144 125526
rect 282092 125462 282144 125468
rect 282104 125225 282132 125462
rect 282090 125216 282146 125225
rect 282090 125151 282146 125160
rect 282840 124545 282868 125530
rect 282826 124536 282882 124545
rect 282826 124471 282882 124480
rect 282276 124160 282328 124166
rect 282276 124102 282328 124108
rect 282288 123729 282316 124102
rect 282828 124092 282880 124098
rect 282828 124034 282880 124040
rect 282274 123720 282330 123729
rect 282274 123655 282330 123664
rect 282840 123049 282868 124034
rect 282826 123040 282882 123049
rect 282826 122975 282882 122984
rect 283116 122834 283144 180095
rect 283196 177336 283248 177342
rect 283196 177278 283248 177284
rect 283208 148918 283236 177278
rect 283196 148912 283248 148918
rect 283196 148854 283248 148860
rect 282932 122806 283144 122834
rect 282460 122800 282512 122806
rect 282460 122742 282512 122748
rect 282472 122233 282500 122742
rect 282458 122224 282514 122233
rect 282458 122159 282514 122168
rect 282644 122120 282696 122126
rect 282644 122062 282696 122068
rect 282092 120080 282144 120086
rect 282092 120022 282144 120028
rect 282104 119241 282132 120022
rect 282656 119921 282684 122062
rect 282828 121440 282880 121446
rect 282826 121408 282828 121417
rect 282880 121408 282882 121417
rect 282826 121343 282882 121352
rect 282642 119912 282698 119921
rect 282642 119847 282698 119856
rect 282184 119400 282236 119406
rect 282184 119342 282236 119348
rect 282090 119232 282146 119241
rect 282090 119167 282146 119176
rect 281816 118448 281868 118454
rect 281814 118416 281816 118425
rect 281868 118416 281870 118425
rect 281814 118351 281870 118360
rect 280250 117600 280306 117609
rect 280250 117535 280306 117544
rect 282000 113076 282052 113082
rect 282000 113018 282052 113024
rect 282012 112305 282040 113018
rect 281998 112296 282054 112305
rect 281998 112231 282054 112240
rect 281724 108928 281776 108934
rect 281724 108870 281776 108876
rect 281736 108497 281764 108870
rect 281722 108488 281778 108497
rect 281722 108423 281778 108432
rect 282196 107817 282224 119342
rect 282828 117292 282880 117298
rect 282828 117234 282880 117240
rect 282368 117156 282420 117162
rect 282368 117098 282420 117104
rect 282380 116113 282408 117098
rect 282840 116929 282868 117234
rect 282826 116920 282882 116929
rect 282826 116855 282882 116864
rect 282366 116104 282422 116113
rect 282366 116039 282422 116048
rect 282828 115932 282880 115938
rect 282828 115874 282880 115880
rect 282840 115433 282868 115874
rect 282826 115424 282882 115433
rect 282276 115388 282328 115394
rect 282826 115359 282882 115368
rect 282276 115330 282328 115336
rect 282288 114617 282316 115330
rect 282274 114608 282330 114617
rect 282274 114543 282330 114552
rect 282826 113792 282882 113801
rect 282932 113778 282960 122806
rect 282882 113750 282960 113778
rect 282826 113727 282882 113736
rect 282828 113144 282880 113150
rect 282826 113112 282828 113121
rect 282880 113112 282882 113121
rect 282826 113047 282882 113056
rect 282828 111784 282880 111790
rect 282828 111726 282880 111732
rect 282840 110809 282868 111726
rect 282826 110800 282882 110809
rect 282826 110735 282882 110744
rect 282276 110424 282328 110430
rect 282276 110366 282328 110372
rect 282288 109993 282316 110366
rect 282274 109984 282330 109993
rect 282274 109919 282330 109928
rect 282828 109812 282880 109818
rect 282828 109754 282880 109760
rect 282840 109313 282868 109754
rect 282826 109304 282882 109313
rect 282826 109239 282882 109248
rect 284312 108934 284340 235214
rect 284392 227792 284444 227798
rect 284392 227734 284444 227740
rect 284404 118454 284432 227734
rect 284484 184204 284536 184210
rect 284484 184146 284536 184152
rect 284496 130626 284524 184146
rect 284576 177404 284628 177410
rect 284576 177346 284628 177352
rect 284588 142118 284616 177346
rect 284576 142112 284628 142118
rect 284576 142054 284628 142060
rect 284484 130620 284536 130626
rect 284484 130562 284536 130568
rect 284392 118448 284444 118454
rect 284392 118390 284444 118396
rect 285692 115394 285720 242218
rect 287242 233880 287298 233889
rect 287242 233815 287298 233824
rect 287152 229764 287204 229770
rect 287152 229706 287204 229712
rect 285772 213240 285824 213246
rect 285772 213182 285824 213188
rect 285784 120086 285812 213182
rect 286324 198008 286376 198014
rect 286324 197950 286376 197956
rect 285864 178696 285916 178702
rect 285864 178638 285916 178644
rect 285876 141370 285904 178638
rect 286336 178022 286364 197950
rect 286324 178016 286376 178022
rect 286324 177958 286376 177964
rect 287060 178016 287112 178022
rect 287060 177958 287112 177964
rect 285956 176248 286008 176254
rect 285956 176190 286008 176196
rect 285968 159798 285996 176190
rect 287072 169658 287100 177958
rect 287060 169652 287112 169658
rect 287060 169594 287112 169600
rect 285956 159792 286008 159798
rect 285956 159734 286008 159740
rect 285864 141364 285916 141370
rect 285864 141306 285916 141312
rect 285772 120080 285824 120086
rect 285772 120022 285824 120028
rect 287164 117162 287192 229706
rect 287256 128246 287284 233815
rect 287244 128240 287296 128246
rect 287244 128182 287296 128188
rect 287152 117156 287204 117162
rect 287152 117098 287204 117104
rect 285680 115388 285732 115394
rect 285680 115330 285732 115336
rect 287348 109818 287376 305050
rect 299572 304292 299624 304298
rect 299572 304234 299624 304240
rect 298742 302288 298798 302297
rect 298742 302223 298798 302232
rect 295340 297424 295392 297430
rect 295340 297366 295392 297372
rect 288438 287328 288494 287337
rect 288438 287263 288494 287272
rect 287336 109812 287388 109818
rect 287336 109754 287388 109760
rect 284300 108928 284352 108934
rect 284300 108870 284352 108876
rect 282276 108316 282328 108322
rect 282276 108258 282328 108264
rect 282182 107808 282238 107817
rect 282182 107743 282238 107752
rect 282000 104780 282052 104786
rect 282000 104722 282052 104728
rect 282012 104009 282040 104722
rect 281998 104000 282054 104009
rect 281998 103935 282054 103944
rect 281538 100872 281594 100881
rect 281538 100807 281594 100816
rect 279422 98832 279478 98841
rect 279422 98767 279478 98776
rect 267738 98288 267794 98297
rect 267738 98223 267794 98232
rect 267280 90364 267332 90370
rect 267280 90306 267332 90312
rect 267752 64190 267780 98223
rect 279330 98152 279386 98161
rect 279330 98087 279386 98096
rect 269118 94888 269174 94897
rect 269118 94823 269174 94832
rect 267740 64184 267792 64190
rect 267740 64126 267792 64132
rect 269132 36650 269160 94823
rect 274008 93838 274036 96084
rect 279344 95169 279372 98087
rect 279330 95160 279386 95169
rect 279330 95095 279386 95104
rect 279436 95033 279464 98767
rect 280066 95840 280122 95849
rect 280066 95775 280122 95784
rect 279422 95024 279478 95033
rect 279422 94959 279478 94968
rect 273996 93832 274048 93838
rect 273996 93774 274048 93780
rect 280080 93673 280108 95775
rect 281552 95198 281580 100807
rect 281724 100700 281776 100706
rect 281724 100642 281776 100648
rect 281736 100201 281764 100642
rect 281722 100192 281778 100201
rect 281722 100127 281778 100136
rect 282288 97889 282316 108258
rect 282828 106276 282880 106282
rect 282828 106218 282880 106224
rect 282840 105505 282868 106218
rect 282826 105496 282882 105505
rect 282826 105431 282882 105440
rect 282828 104848 282880 104854
rect 282828 104790 282880 104796
rect 282840 104689 282868 104790
rect 282826 104680 282882 104689
rect 282826 104615 282882 104624
rect 282828 103488 282880 103494
rect 282828 103430 282880 103436
rect 282840 103193 282868 103430
rect 282826 103184 282882 103193
rect 282736 103148 282788 103154
rect 288452 103154 288480 287263
rect 288532 267028 288584 267034
rect 288532 266970 288584 266976
rect 288544 126954 288572 266970
rect 291200 259480 291252 259486
rect 291200 259422 291252 259428
rect 289820 250504 289872 250510
rect 289820 250446 289872 250452
rect 288624 188352 288676 188358
rect 288624 188294 288676 188300
rect 288636 163198 288664 188294
rect 288714 178936 288770 178945
rect 288714 178871 288770 178880
rect 288728 166462 288756 178871
rect 288716 166456 288768 166462
rect 288716 166398 288768 166404
rect 288624 163192 288676 163198
rect 288624 163134 288676 163140
rect 289832 135250 289860 250446
rect 289910 210488 289966 210497
rect 289910 210423 289966 210432
rect 289820 135244 289872 135250
rect 289820 135186 289872 135192
rect 288532 126948 288584 126954
rect 288532 126890 288584 126896
rect 289924 103494 289952 210423
rect 290002 198112 290058 198121
rect 290002 198047 290058 198056
rect 290016 111790 290044 198047
rect 290096 180260 290148 180266
rect 290096 180202 290148 180208
rect 290108 148986 290136 180202
rect 290096 148980 290148 148986
rect 290096 148922 290148 148928
rect 291212 113082 291240 259422
rect 294052 253224 294104 253230
rect 294052 253166 294104 253172
rect 292580 231872 292632 231878
rect 292580 231814 292632 231820
rect 291384 217320 291436 217326
rect 291384 217262 291436 217268
rect 291292 203584 291344 203590
rect 291292 203526 291344 203532
rect 291200 113076 291252 113082
rect 291200 113018 291252 113024
rect 290004 111784 290056 111790
rect 290004 111726 290056 111732
rect 291304 106282 291332 203526
rect 291396 172514 291424 217262
rect 291476 180192 291528 180198
rect 291476 180134 291528 180140
rect 291384 172508 291436 172514
rect 291384 172450 291436 172456
rect 291488 137970 291516 180134
rect 291476 137964 291528 137970
rect 291476 137906 291528 137912
rect 291292 106276 291344 106282
rect 291292 106218 291344 106224
rect 292592 104786 292620 231814
rect 292672 227044 292724 227050
rect 292672 226986 292724 226992
rect 292684 133822 292712 226986
rect 293958 187096 294014 187105
rect 293958 187031 294014 187040
rect 292856 184272 292908 184278
rect 292856 184214 292908 184220
rect 292762 178800 292818 178809
rect 292762 178735 292818 178744
rect 292672 133816 292724 133822
rect 292672 133758 292724 133764
rect 292776 117298 292804 178735
rect 292868 158710 292896 184214
rect 292856 158704 292908 158710
rect 292856 158646 292908 158652
rect 292764 117292 292816 117298
rect 292764 117234 292816 117240
rect 292580 104780 292632 104786
rect 292580 104722 292632 104728
rect 289912 103488 289964 103494
rect 289912 103430 289964 103436
rect 282826 103119 282882 103128
rect 288440 103148 288492 103154
rect 282736 103090 282788 103096
rect 288440 103090 288492 103096
rect 282748 102377 282776 103090
rect 282734 102368 282790 102377
rect 282734 102303 282790 102312
rect 282828 102128 282880 102134
rect 282828 102070 282880 102076
rect 282840 101697 282868 102070
rect 282826 101688 282882 101697
rect 282826 101623 282882 101632
rect 282274 97880 282330 97889
rect 282274 97815 282330 97824
rect 281722 97064 281778 97073
rect 281722 96999 281778 97008
rect 281540 95192 281592 95198
rect 281540 95134 281592 95140
rect 281736 93770 281764 96999
rect 281724 93764 281776 93770
rect 281724 93706 281776 93712
rect 280066 93664 280122 93673
rect 280066 93599 280122 93608
rect 277398 91760 277454 91769
rect 277398 91695 277454 91704
rect 270498 84824 270554 84833
rect 270498 84759 270554 84768
rect 269120 36644 269172 36650
rect 269120 36586 269172 36592
rect 267188 33856 267240 33862
rect 267188 33798 267240 33804
rect 269120 21480 269172 21486
rect 269120 21422 269172 21428
rect 269132 16574 269160 21422
rect 270512 16574 270540 84759
rect 273258 82240 273314 82249
rect 273258 82175 273314 82184
rect 269132 16546 269712 16574
rect 270512 16546 270816 16574
rect 268382 14512 268438 14521
rect 268382 14447 268438 14456
rect 267740 6180 267792 6186
rect 267740 6122 267792 6128
rect 267004 4888 267056 4894
rect 267004 4830 267056 4836
rect 266542 3632 266598 3641
rect 266542 3567 266598 3576
rect 265176 598 265388 626
rect 265176 490 265204 598
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 264992 462 265204 490
rect 265360 480 265388 598
rect 266556 480 266584 3567
rect 267752 480 267780 6122
rect 268396 490 268424 14447
rect 269684 2938 269712 16546
rect 269764 15972 269816 15978
rect 269764 15914 269816 15920
rect 269776 3126 269804 15914
rect 269764 3120 269816 3126
rect 269764 3062 269816 3068
rect 269684 2910 270080 2938
rect 268672 598 268884 626
rect 268672 490 268700 598
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268396 462 268700 490
rect 268856 480 268884 598
rect 270052 480 270080 2910
rect 270788 490 270816 16546
rect 272432 3120 272484 3126
rect 272432 3062 272484 3068
rect 271064 598 271276 626
rect 271064 490 271092 598
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 270788 462 271092 490
rect 271248 480 271276 598
rect 272444 480 272472 3062
rect 273272 490 273300 82175
rect 276018 65512 276074 65521
rect 276018 65447 276074 65456
rect 276032 16574 276060 65447
rect 277412 16574 277440 91695
rect 280158 87544 280214 87553
rect 280158 87479 280214 87488
rect 278780 33788 278832 33794
rect 278780 33730 278832 33736
rect 278792 16574 278820 33730
rect 280172 16574 280200 87479
rect 281540 83496 281592 83502
rect 281540 83438 281592 83444
rect 280802 22808 280858 22817
rect 280802 22743 280858 22752
rect 276032 16546 276704 16574
rect 277412 16546 278360 16574
rect 278792 16546 279096 16574
rect 280172 16546 280752 16574
rect 274822 3496 274878 3505
rect 274822 3431 274878 3440
rect 273456 598 273668 626
rect 273456 490 273484 598
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273272 462 273484 490
rect 273640 480 273668 598
rect 274836 480 274864 3431
rect 276018 3360 276074 3369
rect 276018 3295 276074 3304
rect 276032 480 276060 3295
rect 276676 490 276704 16546
rect 276952 598 277164 626
rect 276952 490 276980 598
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276676 462 276980 490
rect 277136 480 277164 598
rect 278332 480 278360 16546
rect 279068 490 279096 16546
rect 279344 598 279556 626
rect 279344 490 279372 598
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279068 462 279372 490
rect 279528 480 279556 598
rect 280724 480 280752 16546
rect 280816 3194 280844 22743
rect 280804 3188 280856 3194
rect 280804 3130 280856 3136
rect 281552 490 281580 83438
rect 284298 72448 284354 72457
rect 284298 72383 284354 72392
rect 283104 3188 283156 3194
rect 283104 3130 283156 3136
rect 281736 598 281948 626
rect 281736 490 281764 598
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281552 462 281764 490
rect 281920 480 281948 598
rect 283116 480 283144 3130
rect 284312 480 284340 72383
rect 292578 37904 292634 37913
rect 292578 37839 292634 37848
rect 289820 19984 289872 19990
rect 289820 19926 289872 19932
rect 286598 3496 286654 3505
rect 285404 3460 285456 3466
rect 286598 3431 286654 3440
rect 287794 3496 287850 3505
rect 287794 3431 287850 3440
rect 288990 3496 289046 3505
rect 288990 3431 289046 3440
rect 285404 3402 285456 3408
rect 285416 480 285444 3402
rect 286612 480 286640 3431
rect 287808 480 287836 3431
rect 289004 480 289032 3431
rect 289832 490 289860 19926
rect 291382 3496 291438 3505
rect 291382 3431 291438 3440
rect 290016 598 290228 626
rect 290016 490 290044 598
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289832 462 290044 490
rect 290200 480 290228 598
rect 291396 480 291424 3431
rect 292592 480 292620 37839
rect 293972 6914 294000 187031
rect 294064 124098 294092 253166
rect 294144 207732 294196 207738
rect 294144 207674 294196 207680
rect 294156 133890 294184 207674
rect 294236 182912 294288 182918
rect 294236 182854 294288 182860
rect 294248 154494 294276 182854
rect 294236 154488 294288 154494
rect 294236 154430 294288 154436
rect 295352 143546 295380 297366
rect 296720 256012 296772 256018
rect 296720 255954 296772 255960
rect 295432 231192 295484 231198
rect 295432 231134 295484 231140
rect 295340 143540 295392 143546
rect 295340 143482 295392 143488
rect 294144 133884 294196 133890
rect 294144 133826 294196 133832
rect 294052 124092 294104 124098
rect 294052 124034 294104 124040
rect 295444 100706 295472 231134
rect 295616 196648 295668 196654
rect 295616 196590 295668 196596
rect 295524 181552 295576 181558
rect 295524 181494 295576 181500
rect 295536 122126 295564 181494
rect 295628 154562 295656 196590
rect 295616 154556 295668 154562
rect 295616 154498 295668 154504
rect 295524 122120 295576 122126
rect 295524 122062 295576 122068
rect 296732 108322 296760 255954
rect 298192 245676 298244 245682
rect 298192 245618 298244 245624
rect 298098 220144 298154 220153
rect 298098 220079 298154 220088
rect 296904 198756 296956 198762
rect 296904 198698 296956 198704
rect 296812 192568 296864 192574
rect 296812 192510 296864 192516
rect 296824 110430 296852 192510
rect 296916 139330 296944 198698
rect 296996 185632 297048 185638
rect 296996 185574 297048 185580
rect 297008 161362 297036 185574
rect 296996 161356 297048 161362
rect 296996 161298 297048 161304
rect 296904 139324 296956 139330
rect 296904 139266 296956 139272
rect 296812 110424 296864 110430
rect 296812 110366 296864 110372
rect 296720 108316 296772 108322
rect 296720 108258 296772 108264
rect 295432 100700 295484 100706
rect 295432 100642 295484 100648
rect 296720 32428 296772 32434
rect 296720 32370 296772 32376
rect 296732 16574 296760 32370
rect 296732 16546 297312 16574
rect 293696 6886 294000 6914
rect 293696 480 293724 6886
rect 296076 4140 296128 4146
rect 296076 4082 296128 4088
rect 294878 3904 294934 3913
rect 294878 3839 294934 3848
rect 294892 480 294920 3839
rect 296088 480 296116 4082
rect 297284 480 297312 16546
rect 298112 4146 298140 220079
rect 298204 125526 298232 245618
rect 298756 215966 298784 302223
rect 298744 215960 298796 215966
rect 298744 215902 298796 215908
rect 298744 209092 298796 209098
rect 298744 209034 298796 209040
rect 298284 181484 298336 181490
rect 298284 181426 298336 181432
rect 298296 144838 298324 181426
rect 298756 178090 298784 209034
rect 299478 202192 299534 202201
rect 299478 202127 299534 202136
rect 298744 178084 298796 178090
rect 298744 178026 298796 178032
rect 298374 177304 298430 177313
rect 298374 177239 298430 177248
rect 298388 158030 298416 177239
rect 298376 158024 298428 158030
rect 298376 157966 298428 157972
rect 298284 144832 298336 144838
rect 298284 144774 298336 144780
rect 298192 125520 298244 125526
rect 298192 125462 298244 125468
rect 299492 16574 299520 202127
rect 299584 161430 299612 304234
rect 299664 264240 299716 264246
rect 299664 264182 299716 264188
rect 299572 161424 299624 161430
rect 299572 161366 299624 161372
rect 299676 132394 299704 264182
rect 300858 189952 300914 189961
rect 300858 189887 300914 189896
rect 299756 178084 299808 178090
rect 299756 178026 299808 178032
rect 299768 164218 299796 178026
rect 299756 164212 299808 164218
rect 299756 164154 299808 164160
rect 299664 132388 299716 132394
rect 299664 132330 299716 132336
rect 300872 16574 300900 189887
rect 300964 140690 300992 317426
rect 303620 299532 303672 299538
rect 303620 299474 303672 299480
rect 302240 272536 302292 272542
rect 302240 272478 302292 272484
rect 301044 220108 301096 220114
rect 301044 220050 301096 220056
rect 300952 140684 301004 140690
rect 300952 140626 301004 140632
rect 301056 136542 301084 220050
rect 301134 205048 301190 205057
rect 301134 204983 301190 204992
rect 301148 162790 301176 204983
rect 301136 162784 301188 162790
rect 301136 162726 301188 162732
rect 302252 139398 302280 272478
rect 302422 223000 302478 223009
rect 302422 222935 302478 222944
rect 302332 193860 302384 193866
rect 302332 193802 302384 193808
rect 302240 139392 302292 139398
rect 302240 139334 302292 139340
rect 301044 136536 301096 136542
rect 301044 136478 301096 136484
rect 302344 115938 302372 193802
rect 302436 165578 302464 222935
rect 302516 209160 302568 209166
rect 302516 209102 302568 209108
rect 302424 165572 302476 165578
rect 302424 165514 302476 165520
rect 302528 160070 302556 209102
rect 302516 160064 302568 160070
rect 302516 160006 302568 160012
rect 303632 122806 303660 299474
rect 304262 284336 304318 284345
rect 304262 284271 304318 284280
rect 303710 229800 303766 229809
rect 303710 229735 303766 229744
rect 303620 122800 303672 122806
rect 303620 122742 303672 122748
rect 302332 115932 302384 115938
rect 302332 115874 302384 115880
rect 303724 113150 303752 229735
rect 304276 219434 304304 284271
rect 304264 219428 304316 219434
rect 304264 219370 304316 219376
rect 304262 211984 304318 211993
rect 304262 211919 304318 211928
rect 303804 196716 303856 196722
rect 303804 196658 303856 196664
rect 303816 155854 303844 196658
rect 303804 155848 303856 155854
rect 303804 155790 303856 155796
rect 303712 113144 303764 113150
rect 303712 113086 303764 113092
rect 302240 17332 302292 17338
rect 302240 17274 302292 17280
rect 302252 16574 302280 17274
rect 299492 16546 299704 16574
rect 300872 16546 301544 16574
rect 302252 16546 303200 16574
rect 298100 4140 298152 4146
rect 298100 4082 298152 4088
rect 298466 4040 298522 4049
rect 298466 3975 298522 3984
rect 298480 480 298508 3975
rect 299676 480 299704 16546
rect 300766 3496 300822 3505
rect 300766 3431 300822 3440
rect 300780 480 300808 3431
rect 301516 490 301544 16546
rect 301792 598 302004 626
rect 301792 490 301820 598
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301516 462 301820 490
rect 301976 480 302004 598
rect 303172 480 303200 16546
rect 304276 4010 304304 211919
rect 305012 6914 305040 335407
rect 306380 329180 306432 329186
rect 306380 329122 306432 329128
rect 305184 231124 305236 231130
rect 305184 231066 305236 231072
rect 305090 188320 305146 188329
rect 305090 188255 305146 188264
rect 304920 6886 305040 6914
rect 304356 5568 304408 5574
rect 304356 5510 304408 5516
rect 304264 4004 304316 4010
rect 304264 3946 304316 3952
rect 304368 480 304396 5510
rect 304920 3505 304948 6886
rect 305104 5574 305132 188255
rect 305196 151774 305224 231066
rect 305276 192500 305328 192506
rect 305276 192442 305328 192448
rect 305184 151768 305236 151774
rect 305184 151710 305236 151716
rect 305288 121446 305316 192442
rect 305276 121440 305328 121446
rect 305276 121382 305328 121388
rect 305092 5568 305144 5574
rect 305092 5510 305144 5516
rect 304906 3496 304962 3505
rect 304906 3431 304962 3440
rect 305550 3496 305606 3505
rect 305550 3431 305606 3440
rect 305564 480 305592 3431
rect 306392 490 306420 329122
rect 313924 324964 313976 324970
rect 313924 324906 313976 324912
rect 309140 311160 309192 311166
rect 309140 311102 309192 311108
rect 306564 291236 306616 291242
rect 306564 291178 306616 291184
rect 306470 218648 306526 218657
rect 306470 218583 306526 218592
rect 306484 3466 306512 218583
rect 306576 162858 306604 291178
rect 307758 273320 307814 273329
rect 307758 273255 307814 273264
rect 306656 203652 306708 203658
rect 306656 203594 306708 203600
rect 306564 162852 306616 162858
rect 306564 162794 306616 162800
rect 306668 132462 306696 203594
rect 306656 132456 306708 132462
rect 306656 132398 306708 132404
rect 307772 124166 307800 273255
rect 307850 237416 307906 237425
rect 307850 237351 307906 237360
rect 307760 124160 307812 124166
rect 307760 124102 307812 124108
rect 307864 119406 307892 237351
rect 307944 214600 307996 214606
rect 307944 214542 307996 214548
rect 307956 147626 307984 214542
rect 307944 147620 307996 147626
rect 307944 147562 307996 147568
rect 307852 119400 307904 119406
rect 307852 119342 307904 119348
rect 307850 22672 307906 22681
rect 307850 22607 307906 22616
rect 307864 11762 307892 22607
rect 309152 16574 309180 311102
rect 310518 285696 310574 285705
rect 310518 285631 310574 285640
rect 309230 270600 309286 270609
rect 309230 270535 309286 270544
rect 309244 155922 309272 270535
rect 309324 215960 309376 215966
rect 309324 215902 309376 215908
rect 309232 155916 309284 155922
rect 309232 155858 309284 155864
rect 309336 102134 309364 215902
rect 309416 182844 309468 182850
rect 309416 182786 309468 182792
rect 309428 129742 309456 182786
rect 309416 129736 309468 129742
rect 309416 129678 309468 129684
rect 310532 104854 310560 285631
rect 311992 280832 312044 280838
rect 311992 280774 312044 280780
rect 310612 202156 310664 202162
rect 310612 202098 310664 202104
rect 310624 144906 310652 202098
rect 311898 199336 311954 199345
rect 311898 199271 311954 199280
rect 310612 144900 310664 144906
rect 310612 144842 310664 144848
rect 310520 104848 310572 104854
rect 310520 104790 310572 104796
rect 309324 102128 309376 102134
rect 309324 102070 309376 102076
rect 310520 18624 310572 18630
rect 310520 18566 310572 18572
rect 310532 16574 310560 18566
rect 311912 16574 311940 199271
rect 312004 140758 312032 280774
rect 313372 228404 313424 228410
rect 313372 228346 313424 228352
rect 313280 226364 313332 226370
rect 313280 226306 313332 226312
rect 311992 140752 312044 140758
rect 311992 140694 312044 140700
rect 313292 128314 313320 226306
rect 313384 131102 313412 228346
rect 313372 131096 313424 131102
rect 313372 131038 313424 131044
rect 313280 128308 313332 128314
rect 313280 128250 313332 128256
rect 309152 16546 309824 16574
rect 310532 16546 311480 16574
rect 311912 16546 312216 16574
rect 307852 11756 307904 11762
rect 307852 11698 307904 11704
rect 309048 11756 309100 11762
rect 309048 11698 309100 11704
rect 307944 4004 307996 4010
rect 307944 3946 307996 3952
rect 306472 3460 306524 3466
rect 306472 3402 306524 3408
rect 306576 598 306788 626
rect 306576 490 306604 598
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306392 462 306604 490
rect 306760 480 306788 598
rect 307956 480 307984 3946
rect 309060 480 309088 11698
rect 309796 490 309824 16546
rect 310072 598 310284 626
rect 310072 490 310100 598
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 309796 462 310100 490
rect 310256 480 310284 598
rect 311452 480 311480 16546
rect 312188 490 312216 16546
rect 313830 4856 313886 4865
rect 313830 4791 313886 4800
rect 312464 598 312676 626
rect 312464 490 312492 598
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312188 462 312492 490
rect 312648 480 312676 598
rect 313844 480 313872 4791
rect 313936 3534 313964 324906
rect 318062 306504 318118 306513
rect 318062 306439 318118 306448
rect 316682 300928 316738 300937
rect 316682 300863 316738 300872
rect 314658 282976 314714 282985
rect 314658 282911 314714 282920
rect 314672 125594 314700 282911
rect 316038 206408 316094 206417
rect 316038 206343 316094 206352
rect 314660 125588 314712 125594
rect 314660 125530 314712 125536
rect 316052 3534 316080 206343
rect 316696 195294 316724 300863
rect 316684 195288 316736 195294
rect 316130 195256 316186 195265
rect 316684 195230 316736 195236
rect 316130 195191 316186 195200
rect 316144 16574 316172 195191
rect 317418 17232 317474 17241
rect 317418 17167 317474 17176
rect 317432 16574 317460 17167
rect 316144 16546 316264 16574
rect 317432 16546 318012 16574
rect 313924 3528 313976 3534
rect 313924 3470 313976 3476
rect 315028 3528 315080 3534
rect 315028 3470 315080 3476
rect 316040 3528 316092 3534
rect 316040 3470 316092 3476
rect 315040 480 315068 3470
rect 316236 480 316264 16546
rect 317328 3528 317380 3534
rect 317328 3470 317380 3476
rect 317340 480 317368 3470
rect 317984 490 318012 16546
rect 318076 4826 318104 306439
rect 318798 191040 318854 191049
rect 318798 190975 318854 190984
rect 318812 16574 318840 190975
rect 320192 16574 320220 353262
rect 321572 16574 321600 371311
rect 327080 367124 327132 367130
rect 327080 367066 327132 367072
rect 324318 342272 324374 342281
rect 324318 342207 324374 342216
rect 323582 322144 323638 322153
rect 323582 322079 323638 322088
rect 322938 210352 322994 210361
rect 322938 210287 322994 210296
rect 318812 16546 319760 16574
rect 320192 16546 320496 16574
rect 321572 16546 322152 16574
rect 318064 4820 318116 4826
rect 318064 4762 318116 4768
rect 318352 598 318564 626
rect 318352 490 318380 598
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 317984 462 318380 490
rect 318536 480 318564 598
rect 319732 480 319760 16546
rect 320468 490 320496 16546
rect 320744 598 320956 626
rect 320744 490 320772 598
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320468 462 320772 490
rect 320928 480 320956 598
rect 322124 480 322152 16546
rect 322952 490 322980 210287
rect 323596 3466 323624 322079
rect 324332 3534 324360 342207
rect 325700 195288 325752 195294
rect 325700 195230 325752 195236
rect 324412 29640 324464 29646
rect 324412 29582 324464 29588
rect 324320 3528 324372 3534
rect 324320 3470 324372 3476
rect 323584 3460 323636 3466
rect 323584 3402 323636 3408
rect 323136 598 323348 626
rect 323136 490 323164 598
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 322952 462 323164 490
rect 323320 480 323348 598
rect 324424 480 324452 29582
rect 325712 16574 325740 195230
rect 327092 16574 327120 367066
rect 582378 365120 582434 365129
rect 582378 365055 582434 365064
rect 331218 353424 331274 353433
rect 331218 353359 331274 353368
rect 329838 185600 329894 185609
rect 329838 185535 329894 185544
rect 329852 16574 329880 185535
rect 325712 16546 326384 16574
rect 327092 16546 328040 16574
rect 329852 16546 330432 16574
rect 325608 3528 325660 3534
rect 325608 3470 325660 3476
rect 325620 480 325648 3470
rect 326356 490 326384 16546
rect 326632 598 326844 626
rect 326632 490 326660 598
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326356 462 326660 490
rect 326816 480 326844 598
rect 328012 480 328040 16546
rect 329196 4820 329248 4826
rect 329196 4762 329248 4768
rect 329208 480 329236 4762
rect 330404 480 330432 16546
rect 331232 490 331260 353359
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580184 349081 580212 351863
rect 580170 349072 580226 349081
rect 580170 349007 580226 349016
rect 582392 347750 582420 365055
rect 582380 347744 582432 347750
rect 582380 347686 582432 347692
rect 357438 345128 357494 345137
rect 357438 345063 357494 345072
rect 336002 340912 336058 340921
rect 336002 340847 336058 340856
rect 333978 313984 334034 313993
rect 333978 313919 334034 313928
rect 332690 196616 332746 196625
rect 332690 196551 332746 196560
rect 332704 11762 332732 196551
rect 333992 16574 334020 313919
rect 335358 189680 335414 189689
rect 335358 189615 335414 189624
rect 335372 16574 335400 189615
rect 333992 16546 334664 16574
rect 335372 16546 335952 16574
rect 332692 11756 332744 11762
rect 332692 11698 332744 11704
rect 333888 11756 333940 11762
rect 333888 11698 333940 11704
rect 332692 3460 332744 3466
rect 332692 3402 332744 3408
rect 331416 598 331628 626
rect 331416 490 331444 598
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 462 331444 490
rect 331600 480 331628 598
rect 332704 480 332732 3402
rect 333900 480 333928 11698
rect 334636 490 334664 16546
rect 335924 3346 335952 16546
rect 336016 3534 336044 340847
rect 339498 338192 339554 338201
rect 339498 338127 339554 338136
rect 338118 308408 338174 308417
rect 338118 308343 338174 308352
rect 338132 16574 338160 308343
rect 338132 16546 338712 16574
rect 336004 3528 336056 3534
rect 336004 3470 336056 3476
rect 337476 3528 337528 3534
rect 337476 3470 337528 3476
rect 335924 3318 336320 3346
rect 334912 598 335124 626
rect 334912 490 334940 598
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 334636 462 334940 490
rect 335096 480 335124 598
rect 336292 480 336320 3318
rect 337488 480 337516 3470
rect 338684 480 338712 16546
rect 339512 490 339540 338127
rect 349160 323604 349212 323610
rect 349160 323546 349212 323552
rect 342258 217288 342314 217297
rect 342258 217223 342314 217232
rect 340878 213208 340934 213217
rect 340878 213143 340934 213152
rect 340892 3534 340920 213143
rect 342272 16574 342300 217223
rect 345018 207632 345074 207641
rect 345018 207567 345074 207576
rect 345032 16574 345060 207567
rect 347042 57216 347098 57225
rect 347042 57151 347098 57160
rect 342272 16546 342944 16574
rect 345032 16546 345336 16574
rect 340972 6180 341024 6186
rect 340972 6122 341024 6128
rect 340880 3528 340932 3534
rect 340880 3470 340932 3476
rect 339696 598 339908 626
rect 339696 490 339724 598
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 462 339724 490
rect 339880 480 339908 598
rect 340984 480 341012 6122
rect 342168 3528 342220 3534
rect 342168 3470 342220 3476
rect 342180 480 342208 3470
rect 342916 490 342944 16546
rect 344558 3360 344614 3369
rect 344558 3295 344614 3304
rect 343192 598 343404 626
rect 343192 490 343220 598
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 342916 462 343220 490
rect 343376 480 343404 598
rect 344572 480 344600 3295
rect 345308 490 345336 16546
rect 346952 3324 347004 3330
rect 346952 3266 347004 3272
rect 345584 598 345796 626
rect 345584 490 345612 598
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345308 462 345612 490
rect 345768 480 345796 598
rect 346964 480 346992 3266
rect 347056 3126 347084 57151
rect 349172 6186 349200 323546
rect 356058 215928 356114 215937
rect 356058 215863 356114 215872
rect 351918 211848 351974 211857
rect 351918 211783 351974 211792
rect 349160 6180 349212 6186
rect 349160 6122 349212 6128
rect 351642 3632 351698 3641
rect 351642 3567 351698 3576
rect 350448 3528 350500 3534
rect 348054 3496 348110 3505
rect 350448 3470 350500 3476
rect 348054 3431 348110 3440
rect 347044 3120 347096 3126
rect 347044 3062 347096 3068
rect 348068 480 348096 3431
rect 349252 3120 349304 3126
rect 349252 3062 349304 3068
rect 349264 480 349292 3062
rect 350460 480 350488 3470
rect 351656 480 351684 3567
rect 351932 3330 351960 211783
rect 353298 208992 353354 209001
rect 353298 208927 353354 208936
rect 353312 3534 353340 208927
rect 353300 3528 353352 3534
rect 353300 3470 353352 3476
rect 356072 3369 356100 215863
rect 357452 3505 357480 345063
rect 582378 343768 582434 343777
rect 582378 343703 582434 343712
rect 580264 309188 580316 309194
rect 580264 309130 580316 309136
rect 574742 296848 574798 296857
rect 574742 296783 574798 296792
rect 358818 197976 358874 197985
rect 358818 197911 358874 197920
rect 358832 3641 358860 197911
rect 574756 179382 574784 296783
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 580170 245576 580226 245585
rect 580170 245511 580226 245520
rect 580184 240145 580212 245511
rect 580170 240136 580226 240145
rect 580170 240071 580226 240080
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 580276 192545 580304 309130
rect 580354 272232 580410 272241
rect 580354 272167 580410 272176
rect 580368 261526 580396 272167
rect 580356 261520 580408 261526
rect 580356 261462 580408 261468
rect 580908 220992 580960 220998
rect 580908 220934 580960 220940
rect 580262 192536 580318 192545
rect 580262 192471 580318 192480
rect 580262 186960 580318 186969
rect 580262 186895 580318 186904
rect 574744 179376 574796 179382
rect 574744 179318 574796 179324
rect 580172 179376 580224 179382
rect 580172 179318 580224 179324
rect 580184 179217 580212 179318
rect 580170 179208 580226 179217
rect 580170 179143 580226 179152
rect 580276 59673 580304 186895
rect 580920 126041 580948 220934
rect 580906 126032 580962 126041
rect 580906 125967 580962 125976
rect 580262 59664 580318 59673
rect 580262 59599 580318 59608
rect 582392 16574 582420 343703
rect 582484 291825 582512 418231
rect 582562 404968 582618 404977
rect 582562 404903 582618 404912
rect 582470 291816 582526 291825
rect 582470 291751 582526 291760
rect 582576 291145 582604 404903
rect 582562 291136 582618 291145
rect 582562 291071 582618 291080
rect 582668 276010 582696 471407
rect 582746 378448 582802 378457
rect 582746 378383 582802 378392
rect 582760 282878 582788 378383
rect 582838 325272 582894 325281
rect 582838 325207 582894 325216
rect 582748 282872 582800 282878
rect 582748 282814 582800 282820
rect 582656 276004 582708 276010
rect 582656 275946 582708 275952
rect 582656 268388 582708 268394
rect 582656 268330 582708 268336
rect 582668 232393 582696 268330
rect 582852 247722 582880 325207
rect 583022 312080 583078 312089
rect 583022 312015 583078 312024
rect 582930 298208 582986 298217
rect 582930 298143 582986 298152
rect 582840 247716 582892 247722
rect 582840 247658 582892 247664
rect 582840 234660 582892 234666
rect 582840 234602 582892 234608
rect 582654 232384 582710 232393
rect 582654 232319 582710 232328
rect 582654 225040 582710 225049
rect 582654 224975 582710 224984
rect 582472 223644 582524 223650
rect 582472 223586 582524 223592
rect 582484 86193 582512 223586
rect 582470 86184 582526 86193
rect 582470 86119 582526 86128
rect 582392 16546 582604 16574
rect 358818 3632 358874 3641
rect 358818 3567 358874 3576
rect 582196 3528 582248 3534
rect 357438 3496 357494 3505
rect 582196 3470 582248 3476
rect 357438 3431 357494 3440
rect 356058 3360 356114 3369
rect 351920 3324 351972 3330
rect 356058 3295 356114 3304
rect 351920 3266 351972 3272
rect 581000 3052 581052 3058
rect 581000 2994 581052 3000
rect 581012 480 581040 2994
rect 582208 480 582236 3470
rect 582576 2938 582604 16546
rect 582668 6633 582696 224975
rect 582748 222896 582800 222902
rect 582748 222838 582800 222844
rect 582760 33153 582788 222838
rect 582852 46345 582880 234602
rect 582944 112849 582972 298143
rect 583036 270502 583064 312015
rect 583114 299568 583170 299577
rect 583114 299503 583170 299512
rect 583024 270496 583076 270502
rect 583024 270438 583076 270444
rect 583024 265668 583076 265674
rect 583024 265610 583076 265616
rect 582930 112840 582986 112849
rect 582930 112775 582986 112784
rect 583036 99521 583064 265610
rect 583128 139369 583156 299503
rect 583390 298752 583446 298761
rect 583390 298687 583446 298696
rect 583404 296714 583432 298687
rect 583404 296686 583524 296714
rect 583392 292596 583444 292602
rect 583392 292538 583444 292544
rect 583208 278792 583260 278798
rect 583208 278734 583260 278740
rect 583220 220998 583248 278734
rect 583300 278044 583352 278050
rect 583300 277986 583352 277992
rect 583208 220992 583260 220998
rect 583208 220934 583260 220940
rect 583312 152697 583340 277986
rect 583404 205737 583432 292538
rect 583496 237289 583524 296686
rect 583666 295352 583722 295361
rect 583666 295287 583722 295296
rect 583576 251864 583628 251870
rect 583576 251806 583628 251812
rect 583482 237280 583538 237289
rect 583482 237215 583538 237224
rect 583390 205728 583446 205737
rect 583390 205663 583446 205672
rect 583390 204912 583446 204921
rect 583390 204847 583446 204856
rect 583298 152688 583354 152697
rect 583298 152623 583354 152632
rect 583114 139360 583170 139369
rect 583114 139295 583170 139304
rect 583022 99512 583078 99521
rect 583022 99447 583078 99456
rect 582838 46336 582894 46345
rect 582838 46271 582894 46280
rect 582746 33144 582802 33153
rect 582746 33079 582802 33088
rect 582654 6624 582710 6633
rect 582654 6559 582710 6568
rect 583404 3058 583432 204847
rect 583482 200696 583538 200705
rect 583482 200631 583538 200640
rect 583496 3534 583524 200631
rect 583588 166433 583616 251806
rect 583574 166424 583630 166433
rect 583574 166359 583630 166368
rect 583680 20369 583708 295287
rect 583758 294536 583814 294545
rect 583758 294471 583814 294480
rect 583772 73273 583800 294471
rect 583758 73264 583814 73273
rect 583758 73199 583814 73208
rect 583666 20360 583722 20369
rect 583666 20295 583722 20304
rect 583484 3528 583536 3534
rect 583484 3470 583536 3476
rect 583392 3052 583444 3058
rect 583392 2994 583444 3000
rect 582576 2910 583432 2938
rect 583404 480 583432 2910
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658164 3478 658200
rect 3422 658144 3424 658164
rect 3424 658144 3476 658164
rect 3476 658144 3478 658164
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 2778 619132 2834 619168
rect 2778 619112 2780 619132
rect 2780 619112 2832 619132
rect 2832 619112 2834 619132
rect 3238 606056 3294 606112
rect 3422 579944 3478 580000
rect 3422 566888 3478 566944
rect 3330 553832 3386 553888
rect 52274 590688 52330 590744
rect 3422 527856 3478 527912
rect 3330 501744 3386 501800
rect 2778 462596 2834 462632
rect 2778 462576 2780 462596
rect 2780 462576 2832 462596
rect 2832 462576 2834 462596
rect 3514 514820 3570 514856
rect 3514 514800 3516 514820
rect 3516 514800 3568 514820
rect 3568 514800 3570 514820
rect 4066 475632 4122 475688
rect 3146 449520 3202 449576
rect 3146 423544 3202 423600
rect 3422 410488 3478 410544
rect 2778 397432 2834 397488
rect 3422 388728 3478 388784
rect 3422 371320 3478 371376
rect 2778 345344 2834 345400
rect 3514 358400 3570 358456
rect 7562 328480 7618 328536
rect 4066 319232 4122 319288
rect 3422 306176 3478 306232
rect 2778 293120 2834 293176
rect 3422 267144 3478 267200
rect 3422 254088 3478 254144
rect 3422 241068 3424 241088
rect 3424 241068 3476 241088
rect 3476 241068 3478 241088
rect 3422 241032 3478 241068
rect 3330 214920 3386 214976
rect 3514 207576 3570 207632
rect 3422 201864 3478 201920
rect 3238 162832 3294 162888
rect 2778 149776 2834 149832
rect 3514 188808 3570 188864
rect 3514 136720 3570 136776
rect 3422 110608 3478 110664
rect 3422 97552 3478 97608
rect 41326 449112 41382 449168
rect 32402 328616 32458 328672
rect 33782 327392 33838 327448
rect 3146 84632 3202 84688
rect 30286 83408 30342 83464
rect 12346 80688 12402 80744
rect 5446 79464 5502 79520
rect 3422 71576 3478 71632
rect 3054 58520 3110 58576
rect 3422 45500 3424 45520
rect 3424 45500 3476 45520
rect 3476 45500 3478 45520
rect 3422 45464 3478 45500
rect 3146 32408 3202 32464
rect 110 24112 166 24168
rect 18 6704 74 6760
rect 3974 25472 4030 25528
rect 3422 19352 3478 19408
rect 10966 51720 11022 51776
rect 15842 79328 15898 79384
rect 13726 77832 13782 77888
rect 15106 66816 15162 66872
rect 19246 75112 19302 75168
rect 17866 55800 17922 55856
rect 23386 73752 23442 73808
rect 20534 59880 20590 59936
rect 26146 68176 26202 68232
rect 24766 39208 24822 39264
rect 15934 3304 15990 3360
rect 28906 26832 28962 26888
rect 28814 21256 28870 21312
rect 33046 62736 33102 62792
rect 32402 58656 32458 58712
rect 40682 327256 40738 327312
rect 36542 222944 36598 223000
rect 35806 69536 35862 69592
rect 43994 240080 44050 240136
rect 41234 82048 41290 82104
rect 41142 72392 41198 72448
rect 38566 50224 38622 50280
rect 37186 48864 37242 48920
rect 43994 76472 44050 76528
rect 41878 7656 41934 7712
rect 48134 235728 48190 235784
rect 45282 15816 45338 15872
rect 49606 231784 49662 231840
rect 52366 385600 52422 385656
rect 50894 239944 50950 240000
rect 50894 72528 50950 72584
rect 51722 224168 51778 224224
rect 52274 226208 52330 226264
rect 53470 213832 53526 213888
rect 53562 206896 53618 206952
rect 52366 202816 52422 202872
rect 53654 54440 53710 54496
rect 57702 366288 57758 366344
rect 59174 445848 59230 445904
rect 59082 388864 59138 388920
rect 59266 411304 59322 411360
rect 59174 351872 59230 351928
rect 57886 241440 57942 241496
rect 60554 353912 60610 353968
rect 58990 237904 59046 237960
rect 59082 220768 59138 220824
rect 56506 69672 56562 69728
rect 57886 53080 57942 53136
rect 55034 17176 55090 17232
rect 60554 237088 60610 237144
rect 60462 223488 60518 223544
rect 61106 313112 61162 313168
rect 61382 313112 61438 313168
rect 61842 233144 61898 233200
rect 66074 579672 66130 579728
rect 66810 588240 66866 588296
rect 66258 586508 66260 586528
rect 66260 586508 66312 586528
rect 66312 586508 66314 586528
rect 66258 586472 66314 586508
rect 66810 582412 66866 582448
rect 66810 582392 66812 582412
rect 66812 582392 66864 582412
rect 66864 582392 66866 582412
rect 66994 581052 67050 581088
rect 66994 581032 66996 581052
rect 66996 581032 67048 581052
rect 67048 581032 67050 581052
rect 66902 575592 66958 575648
rect 67454 575320 67510 575376
rect 66442 573144 66498 573200
rect 66442 571784 66498 571840
rect 67270 570152 67326 570208
rect 66810 568792 66866 568848
rect 66902 567432 66958 567488
rect 66626 564576 66682 564632
rect 66442 564032 66498 564088
rect 66442 561992 66498 562048
rect 66626 560360 66682 560416
rect 66626 559000 66682 559056
rect 66350 555192 66406 555248
rect 66258 554684 66260 554704
rect 66260 554684 66312 554704
rect 66312 554684 66314 554704
rect 66258 554648 66314 554684
rect 66534 549616 66590 549672
rect 66534 548256 66590 548312
rect 66810 547576 66866 547632
rect 66166 546352 66222 546408
rect 66810 544856 66866 544912
rect 66810 542680 66866 542736
rect 67086 541728 67142 541784
rect 65982 447752 66038 447808
rect 64602 387640 64658 387696
rect 65890 390904 65946 390960
rect 67546 566752 67602 566808
rect 67730 589872 67786 589928
rect 72974 699488 73030 699544
rect 72422 590824 72478 590880
rect 73618 590688 73674 590744
rect 73158 590008 73214 590064
rect 77942 592048 77998 592104
rect 75642 588784 75698 588840
rect 82542 590960 82598 591016
rect 83738 591912 83794 591968
rect 86866 590824 86922 590880
rect 84106 590688 84162 590744
rect 84382 588648 84438 588704
rect 87878 588648 87934 588704
rect 88890 588376 88946 588432
rect 67730 585792 67786 585848
rect 67730 583752 67786 583808
rect 67638 558864 67694 558920
rect 67362 556280 67418 556336
rect 66994 439864 67050 439920
rect 66810 437688 66866 437744
rect 66810 435240 66866 435296
rect 66902 433064 66958 433120
rect 66902 430888 66958 430944
rect 66810 428440 66866 428496
rect 66258 426264 66314 426320
rect 66258 424088 66314 424144
rect 66258 421912 66314 421968
rect 66902 417288 66958 417344
rect 66442 415148 66444 415168
rect 66444 415148 66496 415168
rect 66496 415148 66498 415168
rect 66442 415112 66498 415148
rect 66534 408312 66590 408368
rect 66626 406136 66682 406192
rect 66350 403688 66406 403744
rect 66810 401548 66812 401568
rect 66812 401548 66864 401568
rect 66864 401548 66866 401568
rect 66810 401512 66866 401548
rect 66350 399336 66406 399392
rect 66994 396888 67050 396944
rect 66258 392536 66314 392592
rect 66166 389136 66222 389192
rect 64602 332832 64658 332888
rect 61934 199280 61990 199336
rect 60646 71032 60702 71088
rect 59266 22616 59322 22672
rect 64602 224848 64658 224904
rect 65982 346296 66038 346352
rect 67454 552200 67510 552256
rect 67362 419464 67418 419520
rect 67454 412664 67510 412720
rect 67362 396888 67418 396944
rect 67362 347656 67418 347712
rect 67178 341128 67234 341184
rect 66074 336912 66130 336968
rect 65982 320184 66038 320240
rect 65522 304680 65578 304736
rect 66074 302504 66130 302560
rect 67178 328344 67234 328400
rect 66810 324808 66866 324864
rect 66810 323720 66866 323776
rect 67270 322632 67326 322688
rect 66258 319368 66314 319424
rect 66350 318280 66406 318336
rect 66258 317500 66260 317520
rect 66260 317500 66312 317520
rect 66312 317500 66314 317520
rect 66258 317464 66314 317500
rect 66442 315288 66498 315344
rect 66258 314220 66314 314256
rect 66258 314200 66260 314220
rect 66260 314200 66312 314220
rect 66312 314200 66314 314220
rect 66258 312024 66314 312080
rect 66810 310936 66866 310992
rect 66626 309848 66682 309904
rect 66810 301416 66866 301472
rect 66442 300600 66498 300656
rect 66810 299512 66866 299568
rect 66626 297336 66682 297392
rect 67822 576952 67878 577008
rect 68650 540776 68706 540832
rect 68466 535472 68522 535528
rect 69662 535472 69718 535528
rect 70674 535472 70730 535528
rect 67730 442040 67786 442096
rect 67546 394712 67602 394768
rect 67638 380160 67694 380216
rect 67546 330112 67602 330168
rect 67086 309032 67142 309088
rect 67178 307944 67234 308000
rect 66442 296248 66498 296304
rect 66810 294092 66866 294128
rect 66810 294072 66812 294092
rect 66812 294072 66864 294092
rect 66864 294072 66866 294092
rect 66994 292984 67050 293040
rect 66902 292168 66958 292224
rect 66810 291080 66866 291136
rect 66810 289992 66866 290048
rect 66718 288904 66774 288960
rect 66626 287816 66682 287872
rect 66810 286728 66866 286784
rect 66810 281580 66866 281616
rect 66810 281560 66812 281580
rect 66812 281560 66864 281580
rect 66864 281560 66866 281580
rect 66810 280472 66866 280528
rect 66442 278296 66498 278352
rect 66810 277208 66866 277264
rect 66166 276120 66222 276176
rect 66810 275304 66866 275360
rect 66810 274216 66866 274272
rect 66810 273128 66866 273184
rect 65890 272040 65946 272096
rect 66810 270952 66866 271008
rect 66810 269864 66866 269920
rect 66626 267688 66682 267744
rect 65982 257352 66038 257408
rect 65890 243344 65946 243400
rect 66810 265784 66866 265840
rect 66718 264696 66774 264752
rect 66810 263608 66866 263664
rect 66810 262520 66866 262576
rect 66810 261432 66866 261488
rect 66258 258068 66260 258088
rect 66260 258068 66312 258088
rect 66312 258068 66314 258088
rect 66258 258032 66314 258068
rect 66810 256264 66866 256320
rect 66810 254088 66866 254144
rect 66994 285640 67050 285696
rect 67362 305768 67418 305824
rect 67546 298424 67602 298480
rect 67546 295160 67602 295216
rect 67086 284552 67142 284608
rect 67546 282648 67602 282704
rect 67178 279384 67234 279440
rect 66810 253000 66866 253056
rect 66442 250008 66498 250064
rect 66810 247832 66866 247888
rect 67270 246744 67326 246800
rect 66626 244568 66682 244624
rect 66810 243480 66866 243536
rect 67086 242800 67142 242856
rect 66166 235864 66222 235920
rect 66074 230424 66130 230480
rect 64694 217232 64750 217288
rect 67454 255176 67510 255232
rect 67454 241712 67510 241768
rect 70306 449112 70362 449168
rect 68742 444760 68798 444816
rect 76746 538056 76802 538112
rect 75918 535472 75974 535528
rect 76746 535472 76802 535528
rect 76562 467744 76618 467800
rect 82726 536696 82782 536752
rect 81438 462848 81494 462904
rect 82726 453192 82782 453248
rect 78770 447752 78826 447808
rect 84750 536016 84806 536072
rect 84106 454688 84162 454744
rect 83462 451288 83518 451344
rect 86958 461488 87014 461544
rect 86866 457408 86922 457464
rect 86222 447752 86278 447808
rect 85578 445848 85634 445904
rect 88338 456048 88394 456104
rect 89166 593408 89222 593464
rect 88798 445712 88854 445768
rect 89902 585656 89958 585712
rect 89810 560088 89866 560144
rect 91098 581576 91154 581632
rect 91098 578856 91154 578912
rect 91098 577496 91154 577552
rect 91926 584568 91982 584624
rect 91926 583652 91928 583672
rect 91928 583652 91980 583672
rect 91980 583652 91982 583672
rect 91926 583616 91982 583652
rect 91190 576680 91246 576736
rect 91098 573416 91154 573472
rect 91190 572056 91246 572112
rect 91098 571412 91100 571432
rect 91100 571412 91152 571432
rect 91152 571412 91154 571432
rect 91098 571376 91154 571412
rect 91098 570016 91154 570072
rect 91926 574796 91982 574832
rect 91926 574776 91928 574796
rect 91928 574776 91980 574796
rect 91980 574776 91982 574796
rect 91742 568656 91798 568712
rect 91282 567860 91338 567896
rect 91282 567840 91284 567860
rect 91284 567840 91336 567860
rect 91336 567840 91338 567860
rect 91098 565836 91100 565856
rect 91100 565836 91152 565856
rect 91152 565836 91154 565856
rect 91098 565800 91154 565836
rect 91098 564460 91154 564496
rect 91098 564440 91100 564460
rect 91100 564440 91152 564460
rect 91152 564440 91154 564460
rect 91098 563100 91154 563136
rect 91098 563080 91100 563100
rect 91100 563080 91152 563100
rect 91152 563080 91154 563100
rect 91098 560904 91154 560960
rect 91190 558184 91246 558240
rect 91190 556824 91246 556880
rect 91190 555464 91246 555520
rect 91282 552744 91338 552800
rect 91190 552100 91192 552120
rect 91192 552100 91244 552120
rect 91244 552100 91246 552120
rect 91190 552064 91246 552100
rect 91190 549344 91246 549400
rect 91190 547848 91246 547904
rect 91282 546508 91338 546544
rect 91282 546488 91284 546508
rect 91284 546488 91336 546508
rect 91336 546488 91338 546508
rect 91282 545400 91338 545456
rect 91282 544040 91338 544096
rect 91282 542428 91338 542464
rect 91282 542408 91284 542428
rect 91284 542408 91336 542428
rect 91336 542408 91338 542428
rect 91282 541320 91338 541376
rect 91282 539708 91338 539744
rect 91282 539688 91284 539708
rect 91284 539688 91336 539708
rect 91336 539688 91338 539708
rect 91834 560088 91890 560144
rect 90132 444488 90188 444544
rect 95882 590824 95938 590880
rect 93766 581576 93822 581632
rect 93122 512624 93178 512680
rect 96434 467064 96490 467120
rect 96526 464344 96582 464400
rect 94410 445712 94466 445768
rect 98642 592048 98698 592104
rect 97906 580896 97962 580952
rect 97906 580216 97962 580272
rect 97262 458088 97318 458144
rect 96618 445712 96674 445768
rect 97354 445712 97410 445768
rect 98734 588648 98790 588704
rect 100666 447752 100722 447808
rect 98642 445712 98698 445768
rect 104254 463528 104310 463584
rect 104162 458224 104218 458280
rect 102138 445712 102194 445768
rect 105542 445848 105598 445904
rect 107106 590960 107162 591016
rect 107014 461488 107070 461544
rect 108302 449928 108358 449984
rect 108946 447888 109002 447944
rect 112442 585384 112498 585440
rect 110418 445712 110474 445768
rect 111430 445712 111486 445768
rect 109498 444624 109554 444680
rect 114466 444760 114522 444816
rect 118698 460128 118754 460184
rect 117318 445712 117374 445768
rect 119020 444624 119076 444680
rect 120814 439864 120870 439920
rect 120814 435240 120870 435296
rect 120722 418920 120778 418976
rect 120630 404232 120686 404288
rect 68650 391176 68706 391232
rect 86314 390904 86370 390960
rect 92846 390904 92902 390960
rect 69938 390360 69994 390416
rect 71870 390360 71926 390416
rect 68466 389000 68522 389056
rect 72054 389000 72110 389056
rect 73066 389000 73122 389056
rect 71042 355272 71098 355328
rect 70030 334192 70086 334248
rect 69294 331200 69350 331256
rect 69294 326984 69350 327040
rect 69938 327004 69994 327040
rect 69938 326984 69940 327004
rect 69940 326984 69992 327004
rect 69992 326984 69994 327004
rect 73066 339632 73122 339688
rect 76562 362208 76618 362264
rect 80058 390360 80114 390416
rect 80610 390360 80666 390416
rect 80058 389136 80114 389192
rect 79322 387640 79378 387696
rect 76562 359216 76618 359272
rect 77206 359216 77262 359272
rect 74630 335552 74686 335608
rect 77206 358808 77262 358864
rect 77298 349696 77354 349752
rect 80058 364928 80114 364984
rect 78586 342216 78642 342272
rect 80794 340992 80850 341048
rect 84106 360848 84162 360904
rect 86222 351056 86278 351112
rect 89810 390360 89866 390416
rect 89718 389000 89774 389056
rect 88890 388864 88946 388920
rect 91282 390360 91338 390416
rect 90362 388728 90418 388784
rect 86866 351056 86922 351112
rect 84106 330248 84162 330304
rect 83646 327528 83702 327584
rect 85670 338272 85726 338328
rect 102138 390904 102194 390960
rect 97354 390360 97410 390416
rect 95882 389000 95938 389056
rect 86498 327528 86554 327584
rect 96434 369552 96490 369608
rect 96434 368464 96490 368520
rect 93766 364248 93822 364304
rect 93122 363024 93178 363080
rect 93766 363024 93822 363080
rect 92386 356632 92442 356688
rect 89442 338408 89498 338464
rect 88614 334056 88670 334112
rect 89810 335416 89866 335472
rect 91742 336776 91798 336832
rect 92662 353232 92718 353288
rect 91236 327664 91292 327720
rect 92386 332424 92442 332480
rect 92386 327664 92442 327720
rect 96526 357992 96582 358048
rect 93858 353504 93914 353560
rect 95054 333240 95110 333296
rect 98826 390360 98882 390416
rect 100666 390360 100722 390416
rect 118698 390904 118754 390960
rect 115754 390632 115810 390688
rect 101126 389000 101182 389056
rect 101954 389000 102010 389056
rect 99286 364384 99342 364440
rect 99194 350648 99250 350704
rect 97906 339496 97962 339552
rect 100022 363704 100078 363760
rect 101402 360848 101458 360904
rect 105082 390360 105138 390416
rect 102046 371320 102102 371376
rect 101402 358944 101458 359000
rect 101954 358944 102010 359000
rect 100022 330384 100078 330440
rect 102690 331336 102746 331392
rect 106554 390360 106610 390416
rect 108026 390360 108082 390416
rect 109498 390360 109554 390416
rect 107474 351056 107530 351112
rect 105542 345616 105598 345672
rect 108854 370640 108910 370696
rect 109682 358672 109738 358728
rect 109682 357448 109738 357504
rect 108946 349288 109002 349344
rect 105542 342352 105598 342408
rect 108854 343712 108910 343768
rect 107842 339768 107898 339824
rect 106002 332560 106058 332616
rect 111338 356088 111394 356144
rect 110418 355816 110474 355872
rect 111798 389000 111854 389056
rect 112626 389000 112682 389056
rect 113178 388592 113234 388648
rect 114098 388592 114154 388648
rect 111706 355816 111762 355872
rect 111706 354728 111762 354784
rect 115938 390360 115994 390416
rect 114558 352008 114614 352064
rect 115846 352008 115902 352064
rect 113086 347928 113142 347984
rect 109958 330248 110014 330304
rect 111706 340856 111762 340912
rect 120722 390632 120778 390688
rect 120170 390360 120226 390416
rect 119342 368328 119398 368384
rect 117318 349152 117374 349208
rect 115938 345752 115994 345808
rect 112166 334328 112222 334384
rect 114742 335688 114798 335744
rect 118606 345072 118662 345128
rect 117134 332696 117190 332752
rect 121550 428440 121606 428496
rect 121550 417288 121606 417344
rect 121458 396888 121514 396944
rect 121642 410488 121698 410544
rect 122930 433064 122986 433120
rect 122838 428440 122894 428496
rect 122654 393216 122710 393272
rect 122746 392536 122802 392592
rect 122654 385600 122710 385656
rect 120814 375400 120870 375456
rect 119342 343848 119398 343904
rect 119342 330384 119398 330440
rect 121458 361664 121514 361720
rect 121458 356632 121514 356688
rect 123022 424088 123078 424144
rect 123022 421912 123078 421968
rect 123114 412664 123170 412720
rect 122930 392536 122986 392592
rect 124126 444216 124182 444272
rect 124126 442040 124182 442096
rect 124126 439864 124182 439920
rect 124126 437688 124182 437744
rect 124126 433064 124182 433120
rect 124126 415148 124128 415168
rect 124128 415148 124180 415168
rect 124180 415148 124182 415168
rect 124126 415112 124182 415148
rect 124126 408312 124182 408368
rect 123206 406156 123262 406192
rect 123206 406136 123208 406156
rect 123208 406136 123260 406156
rect 123260 406136 123262 406156
rect 124126 401532 124182 401568
rect 124126 401512 124128 401532
rect 124128 401512 124180 401532
rect 124180 401512 124182 401532
rect 123482 399336 123538 399392
rect 123666 394712 123722 394768
rect 123022 380160 123078 380216
rect 122838 370504 122894 370560
rect 122930 367648 122986 367704
rect 83922 327120 83978 327176
rect 114466 327392 114522 327448
rect 124954 406272 125010 406328
rect 123298 360168 123354 360224
rect 123298 355272 123354 355328
rect 122930 328616 122986 328672
rect 125506 338136 125562 338192
rect 124954 328480 125010 328536
rect 129002 536016 129058 536072
rect 127622 367104 127678 367160
rect 125690 357992 125746 358048
rect 129002 364248 129058 364304
rect 129002 363568 129058 363624
rect 126978 350512 127034 350568
rect 127714 350512 127770 350568
rect 132498 582936 132554 582992
rect 130382 536696 130438 536752
rect 154118 702480 154174 702536
rect 582378 697176 582434 697232
rect 580262 670656 580318 670712
rect 580170 590960 580226 591016
rect 580170 589872 580226 589928
rect 580262 577632 580318 577688
rect 133142 377304 133198 377360
rect 130382 358128 130438 358184
rect 129094 356632 129150 356688
rect 129646 354864 129702 354920
rect 132038 330384 132094 330440
rect 133878 328480 133934 328536
rect 579802 537784 579858 537840
rect 582470 683848 582526 683904
rect 582562 644000 582618 644056
rect 582378 536016 582434 536072
rect 582654 630808 582710 630864
rect 582746 617480 582802 617536
rect 582746 593408 582802 593464
rect 582746 564304 582802 564360
rect 582470 524456 582526 524512
rect 580170 511284 580226 511320
rect 580170 511264 580172 511284
rect 580172 511264 580224 511284
rect 580224 511264 580226 511284
rect 582378 484608 582434 484664
rect 142802 448568 142858 448624
rect 137282 444488 137338 444544
rect 135902 366968 135958 367024
rect 136546 366968 136602 367024
rect 136546 365744 136602 365800
rect 136546 349832 136602 349888
rect 135166 346976 135222 347032
rect 137282 345208 137338 345264
rect 135166 342488 135222 342544
rect 135258 337048 135314 337104
rect 135074 328616 135130 328672
rect 138018 349832 138074 349888
rect 142066 353368 142122 353424
rect 141974 328752 142030 328808
rect 143354 331472 143410 331528
rect 143354 330384 143410 330440
rect 142802 330112 142858 330168
rect 142894 329976 142950 330032
rect 142802 329024 142858 329080
rect 145562 375944 145618 376000
rect 151726 363704 151782 363760
rect 151082 360848 151138 360904
rect 151174 357312 151230 357368
rect 151726 357312 151782 357368
rect 144918 349696 144974 349752
rect 145562 349696 145618 349752
rect 144182 330112 144238 330168
rect 123574 327392 123630 327448
rect 122838 327256 122894 327312
rect 123666 327256 123722 327312
rect 146206 327664 146262 327720
rect 149886 327392 149942 327448
rect 150714 327120 150770 327176
rect 157338 364928 157394 364984
rect 153842 345616 153898 345672
rect 153382 328752 153438 328808
rect 152830 327120 152886 327176
rect 155222 327664 155278 327720
rect 153382 326984 153438 327040
rect 67822 321544 67878 321600
rect 154854 326848 154910 326904
rect 154670 318280 154726 318336
rect 67730 306856 67786 306912
rect 67638 268776 67694 268832
rect 155406 332832 155462 332888
rect 156694 353912 156750 353968
rect 156050 326440 156106 326496
rect 156142 325352 156198 325408
rect 156050 324264 156106 324320
rect 156050 322088 156106 322144
rect 155958 318008 156014 318064
rect 156602 318008 156658 318064
rect 155406 305632 155462 305688
rect 156050 304136 156106 304192
rect 156418 297880 156474 297936
rect 156326 294616 156382 294672
rect 156510 293528 156566 293584
rect 156050 291624 156106 291680
rect 156418 285096 156474 285152
rect 155314 279248 155370 279304
rect 155314 276664 155370 276720
rect 155222 264152 155278 264208
rect 67822 260344 67878 260400
rect 67730 250824 67786 250880
rect 67638 245656 67694 245712
rect 67362 236544 67418 236600
rect 67270 215872 67326 215928
rect 154946 243208 155002 243264
rect 70306 241848 70362 241904
rect 69662 241712 69718 241768
rect 67086 200640 67142 200696
rect 69754 215192 69810 215248
rect 72974 230288 73030 230344
rect 73158 238176 73214 238232
rect 73802 220632 73858 220688
rect 75366 240896 75422 240952
rect 74722 239944 74778 240000
rect 75458 239944 75514 240000
rect 75090 237904 75146 237960
rect 75090 234504 75146 234560
rect 74722 232872 74778 232928
rect 77298 240080 77354 240136
rect 77942 240080 77998 240136
rect 77206 222808 77262 222864
rect 76562 209616 76618 209672
rect 73066 197920 73122 197976
rect 79322 228656 79378 228712
rect 79874 206216 79930 206272
rect 77942 197240 77998 197296
rect 81254 211928 81310 211984
rect 82956 241440 83012 241496
rect 84106 241440 84162 241496
rect 84014 239808 84070 239864
rect 84106 224712 84162 224768
rect 82726 218728 82782 218784
rect 88246 210296 88302 210352
rect 85486 192480 85542 192536
rect 90914 220088 90970 220144
rect 89626 189760 89682 189816
rect 92386 213152 92442 213208
rect 93858 217776 93914 217832
rect 93766 214512 93822 214568
rect 95146 211792 95202 211848
rect 96618 238448 96674 238504
rect 97906 191120 97962 191176
rect 101954 221448 102010 221504
rect 102138 235592 102194 235648
rect 102138 234640 102194 234696
rect 102782 234640 102838 234696
rect 102782 228792 102838 228848
rect 102046 210432 102102 210488
rect 104254 212472 104310 212528
rect 104162 198464 104218 198520
rect 107474 195744 107530 195800
rect 108302 216552 108358 216608
rect 107566 193840 107622 193896
rect 111614 218592 111670 218648
rect 112534 239944 112590 240000
rect 111706 214648 111762 214704
rect 114374 231104 114430 231160
rect 114466 204176 114522 204232
rect 111062 193160 111118 193216
rect 115846 208936 115902 208992
rect 115294 205536 115350 205592
rect 120262 238312 120318 238368
rect 119342 235728 119398 235784
rect 119434 224984 119490 225040
rect 122654 217912 122710 217968
rect 122746 213288 122802 213344
rect 122930 240760 122986 240816
rect 124310 240216 124366 240272
rect 125414 222128 125470 222184
rect 122838 208256 122894 208312
rect 126702 240896 126758 240952
rect 126242 240760 126298 240816
rect 128174 231648 128230 231704
rect 129554 230152 129610 230208
rect 129002 227296 129058 227352
rect 128266 219272 128322 219328
rect 119342 201320 119398 201376
rect 130382 233008 130438 233064
rect 129646 200776 129702 200832
rect 118606 199416 118662 199472
rect 133602 236544 133658 236600
rect 132406 204992 132462 205048
rect 130382 195880 130438 195936
rect 135166 224984 135222 225040
rect 135994 241984 136050 242040
rect 133786 206352 133842 206408
rect 137098 237224 137154 237280
rect 137098 236816 137154 236872
rect 136638 235592 136694 235648
rect 136638 234640 136694 234696
rect 137374 234640 137430 234696
rect 137466 225528 137522 225584
rect 137282 221992 137338 222048
rect 138202 241984 138258 242040
rect 146758 241984 146814 242040
rect 135166 198600 135222 198656
rect 142342 235728 142398 235784
rect 143446 231104 143502 231160
rect 143354 210976 143410 211032
rect 140686 196560 140742 196616
rect 145930 240352 145986 240408
rect 149058 241460 149114 241496
rect 149058 241440 149060 241460
rect 149060 241440 149112 241460
rect 149112 241440 149114 241460
rect 149150 240760 149206 240816
rect 146758 226072 146814 226128
rect 133142 190984 133198 191040
rect 149058 237224 149114 237280
rect 150438 234368 150494 234424
rect 151082 208936 151138 208992
rect 148966 189896 149022 189952
rect 99286 188264 99342 188320
rect 91006 185680 91062 185736
rect 100666 183640 100722 183696
rect 98918 182144 98974 182200
rect 98918 177520 98974 177576
rect 100758 180920 100814 180976
rect 100758 177520 100814 177576
rect 119526 182280 119582 182336
rect 115846 180784 115902 180840
rect 110234 179424 110290 179480
rect 106186 177520 106242 177576
rect 108946 177520 109002 177576
rect 115846 177520 115902 177576
rect 110234 176976 110290 177032
rect 112258 176976 112314 177032
rect 119526 177520 119582 177576
rect 122746 177520 122802 177576
rect 124126 177520 124182 177576
rect 152554 241984 152610 242040
rect 151818 233008 151874 233064
rect 152462 219272 152518 219328
rect 154026 241596 154082 241632
rect 154026 241576 154028 241596
rect 154028 241576 154080 241596
rect 154080 241576 154082 241596
rect 153842 234232 153898 234288
rect 153014 204040 153070 204096
rect 151726 195200 151782 195256
rect 151082 187040 151138 187096
rect 154394 209072 154450 209128
rect 156510 273672 156566 273728
rect 156418 268232 156474 268288
rect 156326 267416 156382 267472
rect 156418 263064 156474 263120
rect 156510 255720 156566 255776
rect 156510 249464 156566 249520
rect 155406 242936 155462 242992
rect 156050 244024 156106 244080
rect 156234 242120 156290 242176
rect 155498 225528 155554 225584
rect 156970 326848 157026 326904
rect 157246 319948 157248 319968
rect 157248 319948 157300 319968
rect 157300 319948 157302 319968
rect 157246 319912 157302 319948
rect 157246 318844 157302 318880
rect 157246 318824 157248 318844
rect 157248 318824 157300 318844
rect 157300 318824 157302 318844
rect 157246 316920 157302 316976
rect 157154 315832 157210 315888
rect 157246 314744 157302 314800
rect 157246 312568 157302 312624
rect 157246 311480 157302 311536
rect 157246 310392 157302 310448
rect 157154 309576 157210 309632
rect 157246 309168 157302 309224
rect 157246 308488 157302 308544
rect 157246 306332 157302 306368
rect 157246 306312 157248 306332
rect 157248 306312 157300 306332
rect 157300 306312 157302 306332
rect 157246 305244 157302 305280
rect 157246 305224 157248 305244
rect 157248 305224 157300 305244
rect 157300 305224 157302 305244
rect 157246 303048 157302 303104
rect 157246 298968 157302 299024
rect 156694 296792 156750 296848
rect 157246 292712 157302 292768
rect 156786 291080 156842 291136
rect 157246 290536 157302 290592
rect 156786 290128 156842 290184
rect 156694 259800 156750 259856
rect 156602 224576 156658 224632
rect 156602 222944 156658 223000
rect 156602 213832 156658 213888
rect 154486 202136 154542 202192
rect 157246 289448 157302 289504
rect 157246 288360 157302 288416
rect 157062 286184 157118 286240
rect 157154 285504 157210 285560
rect 157154 284280 157210 284336
rect 157246 283212 157302 283248
rect 157246 283192 157248 283212
rect 157248 283192 157300 283212
rect 157300 283192 157302 283212
rect 157246 281016 157302 281072
rect 157246 279928 157302 279984
rect 157246 278840 157302 278896
rect 157246 277752 157302 277808
rect 156878 275848 156934 275904
rect 157246 274760 157302 274816
rect 156970 272584 157026 272640
rect 157246 270408 157302 270464
rect 157246 266364 157248 266384
rect 157248 266364 157300 266384
rect 157300 266364 157302 266384
rect 157246 266328 157302 266364
rect 157246 265240 157302 265296
rect 156970 261976 157026 262032
rect 157246 260908 157302 260944
rect 157246 260888 157248 260908
rect 157248 260888 157300 260908
rect 157300 260888 157302 260908
rect 156878 257932 156880 257952
rect 156880 257932 156932 257952
rect 156932 257932 156934 257952
rect 156878 257896 156934 257932
rect 157246 256808 157302 256864
rect 157246 254652 157302 254688
rect 157246 254632 157248 254652
rect 157248 254632 157300 254652
rect 157300 254632 157302 254652
rect 157246 253580 157248 253600
rect 157248 253580 157300 253600
rect 157300 253580 157302 253600
rect 157246 253544 157302 253580
rect 157154 252456 157210 252512
rect 157246 251368 157302 251424
rect 157246 250552 157302 250608
rect 156970 248376 157026 248432
rect 156786 247288 156842 247344
rect 157246 246200 157302 246256
rect 156786 246064 156842 246120
rect 158074 358128 158130 358184
rect 157338 232872 157394 232928
rect 156786 213832 156842 213888
rect 156694 208936 156750 208992
rect 157338 207032 157394 207088
rect 161478 370640 161534 370696
rect 160098 366288 160154 366344
rect 159638 336912 159694 336968
rect 159454 308352 159510 308408
rect 160742 357312 160798 357368
rect 160742 337320 160798 337376
rect 160926 337048 160982 337104
rect 160742 331336 160798 331392
rect 159362 302776 159418 302832
rect 159362 293120 159418 293176
rect 158718 247152 158774 247208
rect 158718 241576 158774 241632
rect 158074 223080 158130 223136
rect 158718 223080 158774 223136
rect 158258 217776 158314 217832
rect 157982 198464 158038 198520
rect 159454 267008 159510 267064
rect 160834 295296 160890 295352
rect 160834 255856 160890 255912
rect 160742 245112 160798 245168
rect 159454 227296 159510 227352
rect 159362 220632 159418 220688
rect 158718 195744 158774 195800
rect 156602 194112 156658 194168
rect 153106 186904 153162 186960
rect 161018 257216 161074 257272
rect 162122 311072 162178 311128
rect 160834 188400 160890 188456
rect 162674 254496 162730 254552
rect 162766 236952 162822 237008
rect 163594 331472 163650 331528
rect 163686 319368 163742 319424
rect 164146 299376 164202 299432
rect 164974 343848 165030 343904
rect 164882 291216 164938 291272
rect 164882 286320 164938 286376
rect 164882 275304 164938 275360
rect 163594 234368 163650 234424
rect 163502 230288 163558 230344
rect 166906 337320 166962 337376
rect 166354 329024 166410 329080
rect 165710 297356 165766 297392
rect 165710 297336 165712 297356
rect 165712 297336 165764 297356
rect 165764 297336 165766 297356
rect 164974 233824 165030 233880
rect 165526 226072 165582 226128
rect 163686 223488 163742 223544
rect 162306 218728 162362 218784
rect 163042 218728 163098 218784
rect 163042 210976 163098 211032
rect 169206 339768 169262 339824
rect 166446 304136 166502 304192
rect 167642 285504 167698 285560
rect 167642 253136 167698 253192
rect 169114 327256 169170 327312
rect 169206 315288 169262 315344
rect 169206 284416 169262 284472
rect 168378 241440 168434 241496
rect 169206 234504 169262 234560
rect 166262 207576 166318 207632
rect 160742 182824 160798 182880
rect 160006 179968 160062 180024
rect 125966 177520 126022 177576
rect 128266 177520 128322 177576
rect 129646 177520 129702 177576
rect 132406 177520 132462 177576
rect 133142 177520 133198 177576
rect 135166 177520 135222 177576
rect 148230 177520 148286 177576
rect 100666 176704 100722 176760
rect 103426 176704 103482 176760
rect 116950 176704 117006 176760
rect 120998 176704 121054 176760
rect 124494 176704 124550 176760
rect 128174 176740 128176 176760
rect 128176 176740 128228 176760
rect 128228 176740 128230 176760
rect 128174 176704 128230 176740
rect 136086 176724 136142 176760
rect 136086 176704 136088 176724
rect 136088 176704 136140 176724
rect 136140 176704 136142 176724
rect 158994 176724 159050 176760
rect 158994 176704 158996 176724
rect 158996 176704 159048 176724
rect 159048 176704 159050 176724
rect 130750 175616 130806 175672
rect 164882 175208 164938 175264
rect 168378 194384 168434 194440
rect 167642 186904 167698 186960
rect 166354 181328 166410 181384
rect 166538 180920 166594 180976
rect 166354 175480 166410 175536
rect 167734 171536 167790 171592
rect 169114 182280 169170 182336
rect 169206 176976 169262 177032
rect 169298 175208 169354 175264
rect 67454 129240 67510 129296
rect 65338 128016 65394 128072
rect 64786 127064 64842 127120
rect 65338 127064 65394 127120
rect 64694 120128 64750 120184
rect 66166 125160 66222 125216
rect 66074 122576 66130 122632
rect 65890 120808 65946 120864
rect 65890 120128 65946 120184
rect 65982 102312 66038 102368
rect 66074 93064 66130 93120
rect 67362 123528 67418 123584
rect 67270 100680 67326 100736
rect 67546 126248 67602 126304
rect 162122 94832 162178 94888
rect 110142 94696 110198 94752
rect 125414 94696 125470 94752
rect 108118 93472 108174 93528
rect 100022 92384 100078 92440
rect 105726 92384 105782 92440
rect 86498 91704 86554 91760
rect 75274 91160 75330 91216
rect 85486 91160 85542 91216
rect 75274 88168 75330 88224
rect 67270 86808 67326 86864
rect 65982 85448 66038 85504
rect 73066 75248 73122 75304
rect 71042 73888 71098 73944
rect 64786 68312 64842 68368
rect 63406 65456 63462 65512
rect 60830 8880 60886 8936
rect 68926 65592 68982 65648
rect 66718 7520 66774 7576
rect 70214 39344 70270 39400
rect 75826 64096 75882 64152
rect 73802 4800 73858 4856
rect 95146 91296 95202 91352
rect 97906 91296 97962 91352
rect 86774 91160 86830 91216
rect 88246 91160 88302 91216
rect 89626 91160 89682 91216
rect 91006 91160 91062 91216
rect 91926 91160 91982 91216
rect 93214 91160 93270 91216
rect 95054 91160 95110 91216
rect 86498 89528 86554 89584
rect 88246 82728 88302 82784
rect 89626 78512 89682 78568
rect 91926 86672 91982 86728
rect 94962 66952 95018 67008
rect 87602 61376 87658 61432
rect 85670 3440 85726 3496
rect 82082 1944 82138 2000
rect 89626 58520 89682 58576
rect 96526 91160 96582 91216
rect 97814 91160 97870 91216
rect 99194 91160 99250 91216
rect 97906 80008 97962 80064
rect 104530 91704 104586 91760
rect 101954 91296 102010 91352
rect 100574 91160 100630 91216
rect 102046 91160 102102 91216
rect 103334 91160 103390 91216
rect 101954 85312 102010 85368
rect 104714 91160 104770 91216
rect 105542 91160 105598 91216
rect 104530 89664 104586 89720
rect 104162 73072 104218 73128
rect 106186 76608 106242 76664
rect 104806 71168 104862 71224
rect 107566 91160 107622 91216
rect 108026 91160 108082 91216
rect 108026 88032 108082 88088
rect 110326 91296 110382 91352
rect 110234 91160 110290 91216
rect 108302 81368 108358 81424
rect 106922 74432 106978 74488
rect 121458 94424 121514 94480
rect 121734 93472 121790 93528
rect 122102 93064 122158 93120
rect 111614 92384 111670 92440
rect 111706 91160 111762 91216
rect 111062 78376 111118 78432
rect 113454 92384 113510 92440
rect 115478 92384 115534 92440
rect 118054 92384 118110 92440
rect 112626 91704 112682 91760
rect 113362 91160 113418 91216
rect 112626 89392 112682 89448
rect 114282 91160 114338 91216
rect 115570 91704 115626 91760
rect 113362 87896 113418 87952
rect 117134 91296 117190 91352
rect 115662 91160 115718 91216
rect 115202 83952 115258 84008
rect 117042 80824 117098 80880
rect 108946 51856 109002 51912
rect 117226 91160 117282 91216
rect 121182 91704 121238 91760
rect 119710 91296 119766 91352
rect 118514 91160 118570 91216
rect 119894 91160 119950 91216
rect 121366 91160 121422 91216
rect 120078 64232 120134 64288
rect 136086 92420 136088 92440
rect 136088 92420 136140 92440
rect 136140 92420 136142 92440
rect 136086 92384 136142 92420
rect 152094 92404 152150 92440
rect 152094 92384 152096 92404
rect 152096 92384 152148 92404
rect 152148 92384 152150 92404
rect 124862 91976 124918 92032
rect 124034 91432 124090 91488
rect 122746 91160 122802 91216
rect 124126 91160 124182 91216
rect 124770 91160 124826 91216
rect 120078 58656 120134 58712
rect 124770 86536 124826 86592
rect 151542 91432 151598 91488
rect 126518 91160 126574 91216
rect 126886 91160 126942 91216
rect 129646 91160 129702 91216
rect 131026 91160 131082 91216
rect 126886 82592 126942 82648
rect 133786 91160 133842 91216
rect 134522 91160 134578 91216
rect 134522 85176 134578 85232
rect 151726 91296 151782 91352
rect 151634 91160 151690 91216
rect 135902 84088 135958 84144
rect 164974 85176 165030 85232
rect 167642 135224 167698 135280
rect 168286 111732 168288 111752
rect 168288 111732 168340 111752
rect 168340 111732 168342 111752
rect 168286 111696 168342 111732
rect 167826 110064 167882 110120
rect 167734 108704 167790 108760
rect 167642 93608 167698 93664
rect 166538 92112 166594 92168
rect 167918 89528 167974 89584
rect 169022 87896 169078 87952
rect 169574 96600 169630 96656
rect 169298 94832 169354 94888
rect 169206 93064 169262 93120
rect 169114 82728 169170 82784
rect 191102 445848 191158 445904
rect 171230 299376 171286 299432
rect 171138 221992 171194 222048
rect 173162 360848 173218 360904
rect 174542 329976 174598 330032
rect 172426 299376 172482 299432
rect 172426 298696 172482 298752
rect 171874 232872 171930 232928
rect 173162 232736 173218 232792
rect 171874 204992 171930 205048
rect 173806 233008 173862 233064
rect 173346 198056 173402 198112
rect 171966 175344 172022 175400
rect 170402 140800 170458 140856
rect 170402 93472 170458 93528
rect 171874 116456 171930 116512
rect 171782 85312 171838 85368
rect 171874 82592 171930 82648
rect 171966 74432 172022 74488
rect 173254 91024 173310 91080
rect 177394 346568 177450 346624
rect 176014 342488 176070 342544
rect 174634 291352 174690 291408
rect 174726 287272 174782 287328
rect 174634 264152 174690 264208
rect 174634 262520 174690 262576
rect 175922 270544 175978 270600
rect 174726 243888 174782 243944
rect 176106 302232 176162 302288
rect 176566 302232 176622 302288
rect 175922 82184 175978 82240
rect 160742 67088 160798 67144
rect 135258 43424 135314 43480
rect 176198 90888 176254 90944
rect 132958 12960 133014 13016
rect 124862 3440 124918 3496
rect 125874 3440 125930 3496
rect 177578 297472 177634 297528
rect 177486 293936 177542 293992
rect 178774 341128 178830 341184
rect 178866 285776 178922 285832
rect 178682 254496 178738 254552
rect 180154 347928 180210 347984
rect 178958 249872 179014 249928
rect 178866 240216 178922 240272
rect 178682 235728 178738 235784
rect 178682 209072 178738 209128
rect 177486 178200 177542 178256
rect 180062 257216 180118 257272
rect 179050 241440 179106 241496
rect 178958 236816 179014 236872
rect 180062 213288 180118 213344
rect 178866 182144 178922 182200
rect 178774 175208 178830 175264
rect 177578 78376 177634 78432
rect 178958 93064 179014 93120
rect 180246 327528 180302 327584
rect 181442 324400 181498 324456
rect 180246 283192 180302 283248
rect 181626 335552 181682 335608
rect 181534 288632 181590 288688
rect 181442 234504 181498 234560
rect 182178 256672 182234 256728
rect 180338 193976 180394 194032
rect 180246 188400 180302 188456
rect 180154 108296 180210 108352
rect 180062 46144 180118 46200
rect 180062 43424 180118 43480
rect 181442 189896 181498 189952
rect 180338 187584 180394 187640
rect 180338 183640 180394 183696
rect 180246 37848 180302 37904
rect 181626 179288 181682 179344
rect 181534 176840 181590 176896
rect 184202 349288 184258 349344
rect 183466 257216 183522 257272
rect 183466 256672 183522 256728
rect 183466 178608 183522 178664
rect 182914 109112 182970 109168
rect 182822 35128 182878 35184
rect 184386 295296 184442 295352
rect 184754 188400 184810 188456
rect 185766 336776 185822 336832
rect 185674 323584 185730 323640
rect 185766 284824 185822 284880
rect 186318 273400 186374 273456
rect 185766 230424 185822 230480
rect 188526 351872 188582 351928
rect 582654 471416 582710 471472
rect 582470 458088 582526 458144
rect 582378 431568 582434 431624
rect 582470 418240 582526 418296
rect 202142 358944 202198 359000
rect 193862 357448 193918 357504
rect 191102 349016 191158 349072
rect 191746 349016 191802 349072
rect 189722 320728 189778 320784
rect 188434 286320 188490 286376
rect 188434 279384 188490 279440
rect 187054 247288 187110 247344
rect 185674 179424 185730 179480
rect 184478 86672 184534 86728
rect 187698 230460 187700 230480
rect 187700 230460 187752 230480
rect 187752 230460 187754 230480
rect 187698 230424 187754 230460
rect 187698 221992 187754 222048
rect 188986 278840 189042 278896
rect 185582 88984 185638 89040
rect 184662 86536 184718 86592
rect 185766 80008 185822 80064
rect 187974 88168 188030 88224
rect 188434 89664 188490 89720
rect 191102 311072 191158 311128
rect 190366 286048 190422 286104
rect 189906 255856 189962 255912
rect 189814 231512 189870 231568
rect 191194 292576 191250 292632
rect 191746 292576 191802 292632
rect 191194 253136 191250 253192
rect 191102 221584 191158 221640
rect 189814 88032 189870 88088
rect 189722 42064 189778 42120
rect 191654 242528 191710 242584
rect 191654 241576 191710 241632
rect 192850 326304 192906 326360
rect 200762 356088 200818 356144
rect 198002 353504 198058 353560
rect 193954 326984 194010 327040
rect 191746 226888 191802 226944
rect 191286 225936 191342 225992
rect 192482 220224 192538 220280
rect 191194 214648 191250 214704
rect 193954 291080 194010 291136
rect 194506 291080 194562 291136
rect 194506 289992 194562 290048
rect 193034 184320 193090 184376
rect 191286 180784 191342 180840
rect 191194 118224 191250 118280
rect 191194 73072 191250 73128
rect 192574 92248 192630 92304
rect 192482 28192 192538 28248
rect 195334 334192 195390 334248
rect 195978 305632 196034 305688
rect 195978 304952 196034 305008
rect 195334 285640 195390 285696
rect 195150 233824 195206 233880
rect 194690 232872 194746 232928
rect 195150 232872 195206 232928
rect 194506 209072 194562 209128
rect 197266 304952 197322 305008
rect 197266 292576 197322 292632
rect 197082 288768 197138 288824
rect 197358 282376 197414 282432
rect 198002 281560 198058 281616
rect 197358 280744 197414 280800
rect 197358 280200 197414 280256
rect 196898 279248 196954 279304
rect 196622 265784 196678 265840
rect 196622 262248 196678 262304
rect 196622 246200 196678 246256
rect 198186 287408 198242 287464
rect 198094 278704 198150 278760
rect 197358 278024 197414 278080
rect 197358 276700 197360 276720
rect 197360 276700 197412 276720
rect 197412 276700 197414 276720
rect 197082 245112 197138 245168
rect 195518 234368 195574 234424
rect 195426 222944 195482 223000
rect 196622 221448 196678 221504
rect 195426 216552 195482 216608
rect 195426 189896 195482 189952
rect 195334 177384 195390 177440
rect 195518 177112 195574 177168
rect 193954 118768 194010 118824
rect 195242 91704 195298 91760
rect 193954 89392 194010 89448
rect 193862 10240 193918 10296
rect 191102 3440 191158 3496
rect 196714 189760 196770 189816
rect 197174 216008 197230 216064
rect 196806 183096 196862 183152
rect 197358 276664 197414 276700
rect 197358 275032 197414 275088
rect 197358 272856 197414 272912
rect 197450 272312 197506 272368
rect 197450 271496 197506 271552
rect 197358 269320 197414 269376
rect 197358 268776 197414 268832
rect 197358 267960 197414 268016
rect 197358 267144 197414 267200
rect 198738 284280 198794 284336
rect 198646 278704 198702 278760
rect 198554 270952 198610 271008
rect 198186 267008 198242 267064
rect 197450 266600 197506 266656
rect 197358 265240 197414 265296
rect 197450 264424 197506 264480
rect 197358 263628 197414 263664
rect 197358 263608 197360 263628
rect 197360 263608 197412 263628
rect 197412 263608 197414 263628
rect 197358 261432 197414 261488
rect 198002 260888 198058 260944
rect 197358 260072 197414 260128
rect 197358 259256 197414 259312
rect 197450 258712 197506 258768
rect 197450 257896 197506 257952
rect 197358 255720 197414 255776
rect 197358 255176 197414 255232
rect 198554 259392 198610 259448
rect 197450 253544 197506 253600
rect 197358 253000 197414 253056
rect 198002 252184 198058 252240
rect 197358 251640 197414 251696
rect 197358 250824 197414 250880
rect 197358 249464 197414 249520
rect 197358 248684 197360 248704
rect 197360 248684 197412 248704
rect 197412 248684 197414 248704
rect 197358 248648 197414 248684
rect 197358 247832 197414 247888
rect 197358 246472 197414 246528
rect 197450 244296 197506 244352
rect 197358 242936 197414 242992
rect 198002 242528 198058 242584
rect 197542 242120 197598 242176
rect 197358 241576 197414 241632
rect 197358 240760 197414 240816
rect 200026 284552 200082 284608
rect 203062 346568 203118 346624
rect 200762 291080 200818 291136
rect 200762 285640 200818 285696
rect 201406 285640 201462 285696
rect 200762 284552 200818 284608
rect 202234 288496 202290 288552
rect 201958 284008 202014 284064
rect 203154 289992 203210 290048
rect 203706 285776 203762 285832
rect 204258 284416 204314 284472
rect 206282 349424 206338 349480
rect 209042 339632 209098 339688
rect 207662 331200 207718 331256
rect 206282 298152 206338 298208
rect 204994 284824 205050 284880
rect 206098 285640 206154 285696
rect 208490 310528 208546 310584
rect 209134 310528 209190 310584
rect 209962 292576 210018 292632
rect 210514 292848 210570 292904
rect 210882 284280 210938 284336
rect 200026 282920 200082 282976
rect 205362 283872 205418 283928
rect 321558 371320 321614 371376
rect 212906 363568 212962 363624
rect 211986 287544 212042 287600
rect 212354 284416 212410 284472
rect 213642 298696 213698 298752
rect 213458 291352 213514 291408
rect 213826 291760 213882 291816
rect 213826 291352 213882 291408
rect 213642 290400 213698 290456
rect 218242 361800 218298 361856
rect 215298 294072 215354 294128
rect 215298 293120 215354 293176
rect 215298 292576 215354 292632
rect 215206 286592 215262 286648
rect 214746 284280 214802 284336
rect 216954 292848 217010 292904
rect 215942 292576 215998 292632
rect 216954 292576 217010 292632
rect 217322 288632 217378 288688
rect 216770 284552 216826 284608
rect 222842 361664 222898 361720
rect 220082 342352 220138 342408
rect 218702 320184 218758 320240
rect 219162 286048 219218 286104
rect 220174 338408 220230 338464
rect 220174 295432 220230 295488
rect 220726 295432 220782 295488
rect 220082 285776 220138 285832
rect 220726 284008 220782 284064
rect 211618 283872 211674 283928
rect 214470 283872 214526 283928
rect 215942 283872 215998 283928
rect 217414 283872 217470 283928
rect 222934 332560 222990 332616
rect 223026 319368 223082 319424
rect 221554 286592 221610 286648
rect 223486 285776 223542 285832
rect 224314 295296 224370 295352
rect 223946 285640 224002 285696
rect 224314 285640 224370 285696
rect 223762 284008 223818 284064
rect 221278 283872 221334 283928
rect 224682 283872 224738 283928
rect 225602 298696 225658 298752
rect 225418 285640 225474 285696
rect 227442 352008 227498 352064
rect 226982 288632 227038 288688
rect 226522 285776 226578 285832
rect 227902 290400 227958 290456
rect 230478 326304 230534 326360
rect 228362 286592 228418 286648
rect 225234 283872 225290 283928
rect 229742 294072 229798 294128
rect 229742 287000 229798 287056
rect 230386 286592 230442 286648
rect 233974 332696 234030 332752
rect 230754 288768 230810 288824
rect 230110 283872 230166 283928
rect 233698 295296 233754 295352
rect 232778 291488 232834 291544
rect 232502 285640 232558 285696
rect 233974 302776 234030 302832
rect 233974 295296 234030 295352
rect 235538 298696 235594 298752
rect 235262 298016 235318 298072
rect 234618 285640 234674 285696
rect 236182 298016 236238 298072
rect 236182 296792 236238 296848
rect 235998 285640 236054 285696
rect 238114 287408 238170 287464
rect 236734 286320 236790 286376
rect 241242 330112 241298 330168
rect 240782 315288 240838 315344
rect 240782 299512 240838 299568
rect 240230 294480 240286 294536
rect 239034 294072 239090 294128
rect 240230 294072 240286 294128
rect 239954 287272 240010 287328
rect 239586 285776 239642 285832
rect 240782 285640 240838 285696
rect 248418 368464 248474 368520
rect 246302 354728 246358 354784
rect 242254 346704 242310 346760
rect 244094 328480 244150 328536
rect 242254 294616 242310 294672
rect 242162 285504 242218 285560
rect 242622 285504 242678 285560
rect 243818 285640 243874 285696
rect 243634 284008 243690 284064
rect 231582 283872 231638 283928
rect 236734 283872 236790 283928
rect 238666 283872 238722 283928
rect 199474 282784 199530 282840
rect 200026 274524 200028 274544
rect 200028 274524 200080 274544
rect 200080 274524 200082 274544
rect 200026 274488 200082 274524
rect 199382 270136 199438 270192
rect 198738 241440 198794 241496
rect 198830 240216 198886 240272
rect 199566 256536 199622 256592
rect 199474 219272 199530 219328
rect 198002 212608 198058 212664
rect 198278 211112 198334 211168
rect 198002 184184 198058 184240
rect 196898 181464 196954 181520
rect 196714 87488 196770 87544
rect 198094 133048 198150 133104
rect 196622 3440 196678 3496
rect 244094 284008 244150 284064
rect 244094 282920 244150 282976
rect 244278 274488 244334 274544
rect 244002 259256 244058 259312
rect 244554 280200 244610 280256
rect 245474 280220 245530 280256
rect 245474 280200 245476 280220
rect 245476 280200 245528 280220
rect 245528 280200 245530 280220
rect 245658 278840 245714 278896
rect 245750 276684 245806 276720
rect 245750 276664 245752 276684
rect 245752 276664 245804 276684
rect 245804 276664 245806 276684
rect 245658 273672 245714 273728
rect 245934 281560 245990 281616
rect 245934 281016 245990 281072
rect 245934 279420 245936 279440
rect 245936 279420 245988 279440
rect 245988 279420 245990 279440
rect 245934 279384 245990 279420
rect 245934 278060 245936 278080
rect 245936 278060 245988 278080
rect 245988 278060 245990 278080
rect 245934 278024 245990 278060
rect 246026 277480 246082 277536
rect 246302 283212 246358 283248
rect 246302 283192 246304 283212
rect 246304 283192 246356 283212
rect 246356 283192 246358 283212
rect 245934 275848 245990 275904
rect 245842 273128 245898 273184
rect 245842 271496 245898 271552
rect 245750 267960 245806 268016
rect 245934 269592 245990 269648
rect 245934 267416 245990 267472
rect 245934 265784 245990 265840
rect 245750 265240 245806 265296
rect 244554 264424 244610 264480
rect 244462 259528 244518 259584
rect 244370 253000 244426 253056
rect 244002 248376 244058 248432
rect 243910 240488 243966 240544
rect 200118 240352 200174 240408
rect 200946 240080 201002 240136
rect 200578 239672 200634 239728
rect 200302 229744 200358 229800
rect 200210 222944 200266 223000
rect 202050 238584 202106 238640
rect 201590 233824 201646 233880
rect 202234 238176 202290 238232
rect 201498 228656 201554 228712
rect 202142 199416 202198 199472
rect 199382 134136 199438 134192
rect 198278 123392 198334 123448
rect 200762 89120 200818 89176
rect 198186 30912 198242 30968
rect 202786 222808 202842 222864
rect 204902 239672 204958 239728
rect 203522 234368 203578 234424
rect 204074 234368 204130 234424
rect 203062 222808 203118 222864
rect 203338 212472 203394 212528
rect 204810 220768 204866 220824
rect 204810 219408 204866 219464
rect 204810 218728 204866 218784
rect 204994 226072 205050 226128
rect 205362 220768 205418 220824
rect 204994 216144 205050 216200
rect 204994 198600 205050 198656
rect 203522 187176 203578 187232
rect 207938 239536 207994 239592
rect 207386 218048 207442 218104
rect 205914 207032 205970 207088
rect 205914 202272 205970 202328
rect 207754 220224 207810 220280
rect 207754 204992 207810 205048
rect 210330 235456 210386 235512
rect 211066 235592 211122 235648
rect 212170 224984 212226 225040
rect 210422 205536 210478 205592
rect 210698 205536 210754 205592
rect 209778 187584 209834 187640
rect 211066 187584 211122 187640
rect 211066 186904 211122 186960
rect 210422 184184 210478 184240
rect 213642 238584 213698 238640
rect 213090 212608 213146 212664
rect 213734 212608 213790 212664
rect 213182 210432 213238 210488
rect 213734 210432 213790 210488
rect 212722 193160 212778 193216
rect 202234 142704 202290 142760
rect 202234 84768 202290 84824
rect 203522 93744 203578 93800
rect 204994 138080 205050 138136
rect 204902 86128 204958 86184
rect 203706 84088 203762 84144
rect 207754 116456 207810 116512
rect 209134 93880 209190 93936
rect 209226 91568 209282 91624
rect 209226 90344 209282 90400
rect 211894 78512 211950 78568
rect 206282 8880 206338 8936
rect 214194 238448 214250 238504
rect 215206 238584 215262 238640
rect 214562 237224 214618 237280
rect 214102 222128 214158 222184
rect 214470 211112 214526 211168
rect 213826 199416 213882 199472
rect 213918 175616 213974 175672
rect 214102 175208 214158 175264
rect 213918 174936 213974 174992
rect 214010 174256 214066 174312
rect 213918 173576 213974 173632
rect 214010 172896 214066 172952
rect 213918 172216 213974 172272
rect 214010 171536 214066 171592
rect 213918 170312 213974 170368
rect 213918 169652 213974 169688
rect 213918 169632 213920 169652
rect 213920 169632 213972 169652
rect 213972 169632 213974 169652
rect 214010 168952 214066 169008
rect 213918 168292 213974 168328
rect 213918 168272 213920 168292
rect 213920 168272 213972 168292
rect 213972 168272 213974 168292
rect 214010 167592 214066 167648
rect 213918 166948 213920 166968
rect 213920 166948 213972 166968
rect 213972 166948 213974 166968
rect 213918 166912 213974 166948
rect 214010 165688 214066 165744
rect 213918 165008 213974 165064
rect 214010 164328 214066 164384
rect 213918 163648 213974 163704
rect 214010 162968 214066 163024
rect 213918 162288 213974 162344
rect 214010 161744 214066 161800
rect 213918 161064 213974 161120
rect 214010 160384 214066 160440
rect 213918 159704 213974 159760
rect 214010 159024 214066 159080
rect 213918 158344 213974 158400
rect 214010 157664 214066 157720
rect 213918 157120 213974 157176
rect 214010 156440 214066 156496
rect 213918 155760 213974 155816
rect 213918 153720 213974 153776
rect 213918 153040 213974 153096
rect 214010 152496 214066 152552
rect 214010 151136 214066 151192
rect 213918 150476 213974 150512
rect 213918 150456 213920 150476
rect 213920 150456 213972 150476
rect 213972 150456 213974 150476
rect 215390 224984 215446 225040
rect 216586 237224 216642 237280
rect 216034 236000 216090 236056
rect 216586 236000 216642 236056
rect 216034 227432 216090 227488
rect 215942 226344 215998 226400
rect 215390 202816 215446 202872
rect 217414 213832 217470 213888
rect 219530 240080 219586 240136
rect 219438 239400 219494 239456
rect 219530 238856 219586 238912
rect 220174 237360 220230 237416
rect 218702 209616 218758 209672
rect 218702 192616 218758 192672
rect 221370 237360 221426 237416
rect 222290 239944 222346 240000
rect 222290 239672 222346 239728
rect 221922 213832 221978 213888
rect 221002 204176 221058 204232
rect 221462 204176 221518 204232
rect 220174 197240 220230 197296
rect 221554 189080 221610 189136
rect 221462 180104 221518 180160
rect 221554 179288 221610 179344
rect 215298 178064 215354 178120
rect 214930 175888 214986 175944
rect 214654 170992 214710 171048
rect 222934 218184 222990 218240
rect 224222 233824 224278 233880
rect 224866 225936 224922 225992
rect 226706 238312 226762 238368
rect 226890 237088 226946 237144
rect 223394 219272 223450 219328
rect 223394 218184 223450 218240
rect 225602 217912 225658 217968
rect 228362 239672 228418 239728
rect 228178 234504 228234 234560
rect 227718 233824 227774 233880
rect 227718 231648 227774 231704
rect 227626 226208 227682 226264
rect 226982 224576 227038 224632
rect 227718 222808 227774 222864
rect 226338 215192 226394 215248
rect 226338 214784 226394 214840
rect 226982 214784 227038 214840
rect 225694 196288 225750 196344
rect 226982 181600 227038 181656
rect 226338 180648 226394 180704
rect 222842 177928 222898 177984
rect 226338 178608 226394 178664
rect 226338 178472 226394 178528
rect 223486 178200 223542 178256
rect 223394 177248 223450 177304
rect 229098 234504 229154 234560
rect 230570 240080 230626 240136
rect 231122 233960 231178 234016
rect 230202 232872 230258 232928
rect 228638 196288 228694 196344
rect 227810 176704 227866 176760
rect 227718 176160 227774 176216
rect 223670 175888 223726 175944
rect 228362 175888 228418 175944
rect 228546 175888 228602 175944
rect 214930 166368 214986 166424
rect 214838 154400 214894 154456
rect 214562 149776 214618 149832
rect 214010 149096 214066 149152
rect 213918 148416 213974 148472
rect 213918 147872 213974 147928
rect 213918 147192 213974 147248
rect 213918 145832 213974 145888
rect 214470 145152 214526 145208
rect 214010 144472 214066 144528
rect 213918 143792 213974 143848
rect 213918 143248 213974 143304
rect 214010 142568 214066 142624
rect 213274 141888 213330 141944
rect 214010 140528 214066 140584
rect 213918 139848 213974 139904
rect 213918 139168 213974 139224
rect 215942 151816 215998 151872
rect 213918 137264 213974 137320
rect 214010 136584 214066 136640
rect 213918 135904 213974 135960
rect 213918 133900 213920 133920
rect 213920 133900 213972 133920
rect 213972 133900 213974 133920
rect 213918 133864 213974 133900
rect 213918 132640 213974 132696
rect 213918 131960 213974 132016
rect 214746 137944 214802 138000
rect 231490 231784 231546 231840
rect 229282 181328 229338 181384
rect 229374 177928 229430 177984
rect 229190 176840 229246 176896
rect 229190 176568 229246 176624
rect 229282 174548 229338 174584
rect 229282 174528 229284 174548
rect 229284 174528 229336 174548
rect 229336 174528 229338 174548
rect 229190 173304 229246 173360
rect 230018 164872 230074 164928
rect 229742 158072 229798 158128
rect 229742 153720 229798 153776
rect 229374 150592 229430 150648
rect 229098 146784 229154 146840
rect 216034 146512 216090 146568
rect 214562 131280 214618 131336
rect 214010 130600 214066 130656
rect 213918 129920 213974 129976
rect 214010 129240 214066 129296
rect 213918 128696 213974 128752
rect 214010 128016 214066 128072
rect 213918 127336 213974 127392
rect 214010 126656 214066 126712
rect 213918 125976 213974 126032
rect 213918 125296 213974 125352
rect 213918 124072 213974 124128
rect 213366 123392 213422 123448
rect 214010 123392 214066 123448
rect 214010 122712 214066 122768
rect 213918 122032 213974 122088
rect 213918 121352 213974 121408
rect 214010 119992 214066 120048
rect 213918 119448 213974 119504
rect 214010 118088 214066 118144
rect 213918 117428 213974 117464
rect 213918 117408 213920 117428
rect 213920 117408 213972 117428
rect 213972 117408 213974 117428
rect 214010 116728 214066 116784
rect 213918 116048 213974 116104
rect 213918 114824 213974 114880
rect 214010 114144 214066 114200
rect 213918 113464 213974 113520
rect 213918 112104 213974 112160
rect 214010 111424 214066 111480
rect 213918 110744 213974 110800
rect 213918 110200 213974 110256
rect 214010 108840 214066 108896
rect 213918 108160 213974 108216
rect 214930 124616 214986 124672
rect 214838 115368 214894 115424
rect 214746 112784 214802 112840
rect 214562 108296 214618 108352
rect 214010 107480 214066 107536
rect 213918 106800 213974 106856
rect 214010 106120 214066 106176
rect 213918 104932 213920 104952
rect 213920 104932 213972 104952
rect 213972 104932 213974 104952
rect 213918 104896 213974 104932
rect 214378 105576 214434 105632
rect 213918 103556 213974 103592
rect 213918 103536 213920 103556
rect 213920 103536 213972 103556
rect 213972 103536 213974 103556
rect 214010 102856 214066 102912
rect 213918 102212 213920 102232
rect 213920 102212 213972 102232
rect 213972 102212 213974 102232
rect 213918 102176 213974 102212
rect 213918 101496 213974 101552
rect 214378 101360 214434 101416
rect 214010 100272 214066 100328
rect 213918 99592 213974 99648
rect 214010 98912 214066 98968
rect 213918 98232 213974 98288
rect 214838 100952 214894 101008
rect 213458 97552 213514 97608
rect 213918 96328 213974 96384
rect 213458 85448 213514 85504
rect 214838 96872 214894 96928
rect 214838 86808 214894 86864
rect 214746 67088 214802 67144
rect 229926 148280 229982 148336
rect 229742 141072 229798 141128
rect 229742 137128 229798 137184
rect 216126 120672 216182 120728
rect 217230 118360 217286 118416
rect 229098 97824 229154 97880
rect 223670 95920 223726 95976
rect 200762 3304 200818 3360
rect 213182 3304 213238 3360
rect 224222 89120 224278 89176
rect 229098 95260 229154 95296
rect 229098 95240 229100 95260
rect 229100 95240 229152 95260
rect 229152 95240 229154 95260
rect 225602 64232 225658 64288
rect 228362 93064 228418 93120
rect 227074 43424 227130 43480
rect 229834 131960 229890 132016
rect 232594 235592 232650 235648
rect 234066 237496 234122 237552
rect 233514 228928 233570 228984
rect 232962 228792 233018 228848
rect 233882 228248 233938 228304
rect 231858 216688 231914 216744
rect 233330 205672 233386 205728
rect 232042 196696 232098 196752
rect 231766 182008 231822 182064
rect 231766 178200 231822 178256
rect 231490 176568 231546 176624
rect 230846 173848 230902 173904
rect 230754 173712 230810 173768
rect 230662 170448 230718 170504
rect 231766 175228 231822 175264
rect 231766 175208 231768 175228
rect 231768 175208 231820 175228
rect 231820 175208 231822 175228
rect 231490 174664 231546 174720
rect 231582 172760 231638 172816
rect 231766 171844 231768 171864
rect 231768 171844 231820 171864
rect 231820 171844 231822 171864
rect 231766 171808 231822 171844
rect 231122 171400 231178 171456
rect 231214 169904 231270 169960
rect 230938 169496 230994 169552
rect 231674 168952 231730 169008
rect 230938 167592 230994 167648
rect 231674 167048 231730 167104
rect 231306 166096 231362 166152
rect 231674 165688 231730 165744
rect 231122 164328 231178 164384
rect 231490 163784 231546 163840
rect 231582 162832 231638 162888
rect 231766 161880 231822 161936
rect 231766 160928 231822 160984
rect 231582 160656 231638 160712
rect 231306 160520 231362 160576
rect 231766 160012 231768 160032
rect 231768 160012 231820 160032
rect 231820 160012 231822 160032
rect 231766 159976 231822 160012
rect 231674 159568 231730 159624
rect 231582 159024 231638 159080
rect 230938 158616 230994 158672
rect 231490 157664 231546 157720
rect 231122 157392 231178 157448
rect 230754 155216 230810 155272
rect 230662 152496 230718 152552
rect 230754 148688 230810 148744
rect 231766 156712 231822 156768
rect 231490 155760 231546 155816
rect 231674 154300 231676 154320
rect 231676 154300 231728 154320
rect 231728 154300 231730 154320
rect 231674 154264 231730 154300
rect 231766 153856 231822 153912
rect 231582 153312 231638 153368
rect 231766 153040 231822 153096
rect 232042 174528 232098 174584
rect 231950 164736 232006 164792
rect 233422 182960 233478 183016
rect 232502 165552 232558 165608
rect 232042 163376 232098 163432
rect 231858 152904 231914 152960
rect 231766 151952 231822 152008
rect 231122 151544 231178 151600
rect 231766 151000 231822 151056
rect 231674 150864 231730 150920
rect 231490 149096 231546 149152
rect 230846 147736 230902 147792
rect 230754 145832 230810 145888
rect 230754 144608 230810 144664
rect 230754 143928 230810 143984
rect 230294 143384 230350 143440
rect 230662 140664 230718 140720
rect 230018 137264 230074 137320
rect 230938 135360 230994 135416
rect 231766 150048 231822 150104
rect 231766 148144 231822 148200
rect 231674 147192 231730 147248
rect 231398 146920 231454 146976
rect 231306 144336 231362 144392
rect 231766 146240 231822 146296
rect 232686 154944 232742 155000
rect 231766 144744 231822 144800
rect 231766 142976 231822 143032
rect 231306 141616 231362 141672
rect 231122 131144 231178 131200
rect 230570 129784 230626 129840
rect 230754 128832 230810 128888
rect 231306 139712 231362 139768
rect 231766 138216 231822 138272
rect 231582 136856 231638 136912
rect 231214 130600 231270 130656
rect 231398 135904 231454 135960
rect 231766 134952 231822 135008
rect 231674 134408 231730 134464
rect 231490 134000 231546 134056
rect 231674 132504 231730 132560
rect 231766 132096 231822 132152
rect 231766 130192 231822 130248
rect 231766 129240 231822 129296
rect 231122 127336 231178 127392
rect 230938 126384 230994 126440
rect 231306 128968 231362 129024
rect 231214 125976 231270 126032
rect 231766 127880 231822 127936
rect 231766 126948 231822 126984
rect 231766 126928 231768 126948
rect 231768 126928 231820 126948
rect 231820 126928 231822 126948
rect 231306 125432 231362 125488
rect 230478 124480 230534 124536
rect 230018 121760 230074 121816
rect 229926 105576 229982 105632
rect 231122 124752 231178 124808
rect 230662 120264 230718 120320
rect 230938 117952 230994 118008
rect 230754 116048 230810 116104
rect 230938 114552 230994 114608
rect 230570 113600 230626 113656
rect 230570 102720 230626 102776
rect 231766 124108 231768 124128
rect 231768 124108 231820 124128
rect 231820 124108 231822 124128
rect 231766 124072 231822 124108
rect 231398 123120 231454 123176
rect 231766 122168 231822 122224
rect 231490 121624 231546 121680
rect 231766 121216 231822 121272
rect 231214 120672 231270 120728
rect 231306 112240 231362 112296
rect 231766 119992 231822 120048
rect 231766 119312 231822 119368
rect 231490 118904 231546 118960
rect 231674 117952 231730 118008
rect 231582 117408 231638 117464
rect 231490 116456 231546 116512
rect 231490 115096 231546 115152
rect 231766 117000 231822 117056
rect 231398 111288 231454 111344
rect 231306 111016 231362 111072
rect 231214 109792 231270 109848
rect 231214 107072 231270 107128
rect 231398 107888 231454 107944
rect 231122 104624 231178 104680
rect 231306 104216 231362 104272
rect 231306 103672 231362 103728
rect 231674 113192 231730 113248
rect 231766 112648 231822 112704
rect 231674 111716 231730 111752
rect 231674 111696 231676 111716
rect 231676 111696 231728 111716
rect 231728 111696 231730 111716
rect 231766 110744 231822 110800
rect 231766 109384 231822 109440
rect 231766 108432 231822 108488
rect 231766 106528 231822 106584
rect 231766 105168 231822 105224
rect 231490 103264 231546 103320
rect 231306 102856 231362 102912
rect 231214 101768 231270 101824
rect 231214 98912 231270 98968
rect 231122 98776 231178 98832
rect 230754 96600 230810 96656
rect 230478 96192 230534 96248
rect 231214 97552 231270 97608
rect 231214 96464 231270 96520
rect 231582 102312 231638 102368
rect 231398 101360 231454 101416
rect 231582 101360 231638 101416
rect 231674 100816 231730 100872
rect 231766 100408 231822 100464
rect 231674 99864 231730 99920
rect 231582 99456 231638 99512
rect 231398 98504 231454 98560
rect 235262 237360 235318 237416
rect 234986 233144 235042 233200
rect 234618 225120 234674 225176
rect 233882 206896 233938 206952
rect 233882 205672 233938 205728
rect 233882 194112 233938 194168
rect 233882 182960 233938 183016
rect 233882 179968 233938 180024
rect 233882 154808 233938 154864
rect 234066 166912 234122 166968
rect 236458 240080 236514 240136
rect 235906 238584 235962 238640
rect 237930 240080 237986 240136
rect 237378 237360 237434 237416
rect 235446 207848 235502 207904
rect 236182 181600 236238 181656
rect 235354 181328 235410 181384
rect 236090 178336 236146 178392
rect 235998 170312 236054 170368
rect 234618 157120 234674 157176
rect 232870 133456 232926 133512
rect 232778 116456 232834 116512
rect 232686 98640 232742 98696
rect 232594 53080 232650 53136
rect 232870 102720 232926 102776
rect 234250 123392 234306 123448
rect 235538 163104 235594 163160
rect 235446 153176 235502 153232
rect 234158 75112 234214 75168
rect 236366 166640 236422 166696
rect 236826 157528 236882 157584
rect 236734 136856 236790 136912
rect 236642 125024 236698 125080
rect 235538 122576 235594 122632
rect 235538 120672 235594 120728
rect 236642 120128 236698 120184
rect 239218 239944 239274 240000
rect 238942 238756 238944 238776
rect 238944 238756 238996 238776
rect 238996 238756 238998 238776
rect 238942 238720 238998 238756
rect 238850 233008 238906 233064
rect 240690 236952 240746 237008
rect 239770 224712 239826 224768
rect 239402 199552 239458 199608
rect 238850 187176 238906 187232
rect 238298 173984 238354 174040
rect 238114 130056 238170 130112
rect 238022 116864 238078 116920
rect 237010 98640 237066 98696
rect 241794 238584 241850 238640
rect 241794 237496 241850 237552
rect 241518 209072 241574 209128
rect 239402 167048 239458 167104
rect 238942 165552 238998 165608
rect 238758 144880 238814 144936
rect 239402 124480 239458 124536
rect 238114 76472 238170 76528
rect 238022 50224 238078 50280
rect 238022 46144 238078 46200
rect 240874 152360 240930 152416
rect 240874 149368 240930 149424
rect 239678 103944 239734 104000
rect 239494 98640 239550 98696
rect 240138 42064 240194 42120
rect 236642 4800 236698 4856
rect 195242 1944 195298 2000
rect 239310 2080 239366 2136
rect 240874 107480 240930 107536
rect 241610 198192 241666 198248
rect 242714 235728 242770 235784
rect 243634 238856 243690 238912
rect 244370 245112 244426 245168
rect 244094 241304 244150 241360
rect 243266 228248 243322 228304
rect 244278 224712 244334 224768
rect 242254 216144 242310 216200
rect 242162 186360 242218 186416
rect 241702 184320 241758 184376
rect 241610 168544 241666 168600
rect 241518 146920 241574 146976
rect 242254 156576 242310 156632
rect 241058 106256 241114 106312
rect 241058 75248 241114 75304
rect 242346 145288 242402 145344
rect 242346 117952 242402 118008
rect 242254 109384 242310 109440
rect 245842 263880 245898 263936
rect 245658 263064 245714 263120
rect 245750 260072 245806 260128
rect 245658 257352 245714 257408
rect 245658 253000 245714 253056
rect 245106 250280 245162 250336
rect 244646 243752 244702 243808
rect 245842 258712 245898 258768
rect 245934 258168 245990 258224
rect 245934 256572 245936 256592
rect 245936 256572 245988 256592
rect 245988 256572 245990 256592
rect 245934 256536 245990 256572
rect 245934 255196 245990 255232
rect 245934 255176 245936 255196
rect 245936 255176 245988 255196
rect 245988 255176 245990 255196
rect 245842 254360 245898 254416
rect 245934 253852 245936 253872
rect 245936 253852 245988 253872
rect 245988 253852 245990 253872
rect 245934 253816 245990 253852
rect 245934 252184 245990 252240
rect 245842 251640 245898 251696
rect 245934 249464 245990 249520
rect 245934 248104 245990 248160
rect 245842 246472 245898 246528
rect 245934 244568 245990 244624
rect 245934 242392 245990 242448
rect 245842 235864 245898 235920
rect 245750 221584 245806 221640
rect 242990 205128 243046 205184
rect 243634 160384 243690 160440
rect 245842 204176 245898 204232
rect 244370 172352 244426 172408
rect 244554 178064 244610 178120
rect 243634 119720 243690 119776
rect 243726 107888 243782 107944
rect 243634 102176 243690 102232
rect 242346 69536 242402 69592
rect 245014 142432 245070 142488
rect 244278 96464 244334 96520
rect 247222 290128 247278 290184
rect 246486 274488 246542 274544
rect 246118 272176 246174 272232
rect 246394 272176 246450 272232
rect 246118 270952 246174 271008
rect 246302 270136 246358 270192
rect 246394 260888 246450 260944
rect 246394 245928 246450 245984
rect 246394 204176 246450 204232
rect 247130 262248 247186 262304
rect 247222 255992 247278 256048
rect 247222 231512 247278 231568
rect 246026 164872 246082 164928
rect 245934 161472 245990 161528
rect 245750 144744 245806 144800
rect 245198 142704 245254 142760
rect 245106 103672 245162 103728
rect 245014 98776 245070 98832
rect 247682 178744 247738 178800
rect 246578 134408 246634 134464
rect 246394 119992 246450 120048
rect 246302 59880 246358 59936
rect 246486 95240 246542 95296
rect 246486 79464 246542 79520
rect 248694 294616 248750 294672
rect 249982 291216 250038 291272
rect 251362 338272 251418 338328
rect 251270 283464 251326 283520
rect 248602 195880 248658 195936
rect 248510 189080 248566 189136
rect 248510 156168 248566 156224
rect 248602 151000 248658 151056
rect 249154 150728 249210 150784
rect 249062 132504 249118 132560
rect 247958 123528 248014 123584
rect 247774 110744 247830 110800
rect 247682 65592 247738 65648
rect 248418 71032 248474 71088
rect 247774 51856 247830 51912
rect 246394 3576 246450 3632
rect 247590 3440 247646 3496
rect 249154 108976 249210 109032
rect 251270 278840 251326 278896
rect 250534 133592 250590 133648
rect 251454 293936 251510 293992
rect 252558 292712 252614 292768
rect 251546 292576 251602 292632
rect 251546 170312 251602 170368
rect 251822 165688 251878 165744
rect 250442 115776 250498 115832
rect 250442 108024 250498 108080
rect 249338 90344 249394 90400
rect 249246 73752 249302 73808
rect 249062 68312 249118 68368
rect 252926 235900 252928 235920
rect 252928 235900 252980 235920
rect 252980 235900 252982 235920
rect 252926 235864 252982 235900
rect 252558 157936 252614 157992
rect 251822 128968 251878 129024
rect 251822 117544 251878 117600
rect 250810 102856 250866 102912
rect 250626 93064 250682 93120
rect 250534 66952 250590 67008
rect 254030 176568 254086 176624
rect 253202 168408 253258 168464
rect 253202 128288 253258 128344
rect 252098 86128 252154 86184
rect 254674 172760 254730 172816
rect 254582 170176 254638 170232
rect 254582 123392 254638 123448
rect 254582 114824 254638 114880
rect 256790 297336 256846 297392
rect 256790 261160 256846 261216
rect 262218 357992 262274 358048
rect 258078 240080 258134 240136
rect 258170 238584 258226 238640
rect 256698 174256 256754 174312
rect 257434 171536 257490 171592
rect 256790 162424 256846 162480
rect 254766 111968 254822 112024
rect 256146 80688 256202 80744
rect 256238 68176 256294 68232
rect 260102 287408 260158 287464
rect 260102 174392 260158 174448
rect 259458 153040 259514 153096
rect 258814 151952 258870 152008
rect 257526 146512 257582 146568
rect 257526 124752 257582 124808
rect 257342 64096 257398 64152
rect 257526 76608 257582 76664
rect 258078 35128 258134 35184
rect 255318 19896 255374 19952
rect 259090 148280 259146 148336
rect 259090 147872 259146 147928
rect 258906 113328 258962 113384
rect 258814 110336 258870 110392
rect 260102 121624 260158 121680
rect 258906 77832 258962 77888
rect 251178 11600 251234 11656
rect 252374 3440 252430 3496
rect 260286 101360 260342 101416
rect 263690 349152 263746 349208
rect 262862 285776 262918 285832
rect 304998 335416 305054 335472
rect 267002 310528 267058 310584
rect 264242 284416 264298 284472
rect 263690 266464 263746 266520
rect 263598 224848 263654 224904
rect 263598 224440 263654 224496
rect 264242 224440 264298 224496
rect 268382 295432 268438 295488
rect 267002 193976 267058 194032
rect 269762 181464 269818 181520
rect 272522 304952 272578 305008
rect 271142 185680 271198 185736
rect 272522 177384 272578 177440
rect 276754 216008 276810 216064
rect 278042 179424 278098 179480
rect 276754 178880 276810 178936
rect 278778 176976 278834 177032
rect 264978 175616 265034 175672
rect 265070 175208 265126 175264
rect 264978 174800 265034 174856
rect 265070 173576 265126 173632
rect 264978 172644 265034 172680
rect 264978 172624 264980 172644
rect 264980 172624 265032 172644
rect 265032 172624 265034 172644
rect 265070 172216 265126 172272
rect 264978 171400 265034 171456
rect 265070 170992 265126 171048
rect 264978 170040 265034 170096
rect 264978 169632 265034 169688
rect 264242 169224 264298 169280
rect 261758 164464 261814 164520
rect 260378 83408 260434 83464
rect 263046 162832 263102 162888
rect 262862 138216 262918 138272
rect 262126 120672 262182 120728
rect 262310 119448 262366 119504
rect 262310 119040 262366 119096
rect 262218 116864 262274 116920
rect 262218 116048 262274 116104
rect 262770 108296 262826 108352
rect 262770 107888 262826 107944
rect 261758 100816 261814 100872
rect 262678 96328 262734 96384
rect 261758 73888 261814 73944
rect 262218 69672 262274 69728
rect 261574 54440 261630 54496
rect 262954 135632 263010 135688
rect 265162 168816 265218 168872
rect 264978 167864 265034 167920
rect 265070 167456 265126 167512
rect 265070 166640 265126 166696
rect 264978 166232 265034 166288
rect 264978 165280 265034 165336
rect 267830 164600 267886 164656
rect 265622 164328 265678 164384
rect 267830 164328 267886 164384
rect 265070 164056 265126 164112
rect 264978 163648 265034 163704
rect 265162 162288 265218 162344
rect 265070 161880 265126 161936
rect 264978 161508 264980 161528
rect 264980 161508 265032 161528
rect 265032 161508 265034 161528
rect 264978 161472 265034 161508
rect 265070 161064 265126 161120
rect 264978 160248 265034 160304
rect 265070 159704 265126 159760
rect 264978 158888 265034 158944
rect 264978 158480 265034 158536
rect 265162 158072 265218 158128
rect 265070 157120 265126 157176
rect 264978 156712 265034 156768
rect 265162 156576 265218 156632
rect 265162 155896 265218 155952
rect 264978 154536 265034 154592
rect 265714 156304 265770 156360
rect 265254 153720 265310 153776
rect 265070 152904 265126 152960
rect 264978 152496 265034 152552
rect 264242 118904 264298 118960
rect 263046 102584 263102 102640
rect 263230 97824 263286 97880
rect 263138 88984 263194 89040
rect 263046 82048 263102 82104
rect 262954 58520 263010 58576
rect 263598 30912 263654 30968
rect 261758 12960 261814 13016
rect 259458 10240 259514 10296
rect 264978 151544 265034 151600
rect 264426 114416 264482 114472
rect 265070 151136 265126 151192
rect 264978 150320 265034 150376
rect 265162 149912 265218 149968
rect 264978 148960 265034 149016
rect 265622 148552 265678 148608
rect 265162 146376 265218 146432
rect 265070 145968 265126 146024
rect 264978 145152 265034 145208
rect 264978 144744 265034 144800
rect 265254 143792 265310 143848
rect 264978 143384 265034 143440
rect 265162 142976 265218 143032
rect 265070 142196 265072 142216
rect 265072 142196 265124 142216
rect 265124 142196 265126 142216
rect 265070 142160 265126 142196
rect 264978 140820 265034 140856
rect 264978 140800 264980 140820
rect 264980 140800 265032 140820
rect 265032 140800 265034 140820
rect 264978 139576 265034 139632
rect 264978 138624 265034 138680
rect 264978 137400 265034 137456
rect 265070 136584 265126 136640
rect 265346 141752 265402 141808
rect 265806 155488 265862 155544
rect 266266 154128 266322 154184
rect 279146 188536 279202 188592
rect 279422 179016 279478 179072
rect 279238 176704 279294 176760
rect 279330 175208 279386 175264
rect 279422 174392 279478 174448
rect 279330 165824 279386 165880
rect 279330 150592 279386 150648
rect 265898 147328 265954 147384
rect 265806 139984 265862 140040
rect 265346 134408 265402 134464
rect 265622 134408 265678 134464
rect 264978 134000 265034 134056
rect 265070 133592 265126 133648
rect 264978 133048 265034 133104
rect 264978 131824 265034 131880
rect 265070 131416 265126 131472
rect 264978 130464 265034 130520
rect 264978 129648 265034 129704
rect 264978 127472 265034 127528
rect 264978 126248 265034 126304
rect 264610 125296 264666 125352
rect 264978 124888 265034 124944
rect 264978 124072 265034 124128
rect 265070 123256 265126 123312
rect 264978 122304 265034 122360
rect 264978 121080 265034 121136
rect 265070 118496 265126 118552
rect 264978 118088 265034 118144
rect 264978 117136 265034 117192
rect 265070 116320 265126 116376
rect 264978 115504 265034 115560
rect 265070 114144 265126 114200
rect 264978 113736 265034 113792
rect 264978 112512 265034 112568
rect 265070 111560 265126 111616
rect 264978 111152 265034 111208
rect 264426 110336 264482 110392
rect 264334 80824 264390 80880
rect 264978 109928 265034 109984
rect 265070 108976 265126 109032
rect 264978 107772 265034 107808
rect 264978 107752 264980 107772
rect 264980 107752 265032 107772
rect 265032 107752 265034 107772
rect 265070 107344 265126 107400
rect 264978 106936 265034 106992
rect 264978 105984 265034 106040
rect 265070 105576 265126 105632
rect 264978 104760 265034 104816
rect 264978 103400 265034 103456
rect 264794 102992 264850 103048
rect 264978 101768 265034 101824
rect 265070 101224 265126 101280
rect 264978 99592 265034 99648
rect 264794 98640 264850 98696
rect 264978 98640 265034 98696
rect 264978 97416 265034 97472
rect 265070 96600 265126 96656
rect 264426 71168 264482 71224
rect 265714 125840 265770 125896
rect 279422 147056 279478 147112
rect 280158 145832 280214 145888
rect 267094 136176 267150 136232
rect 265898 135224 265954 135280
rect 267002 122848 267058 122904
rect 265898 97008 265954 97064
rect 265898 79328 265954 79384
rect 265622 61376 265678 61432
rect 264978 28192 265034 28248
rect 267278 120672 267334 120728
rect 267186 105168 267242 105224
rect 280434 179424 280490 179480
rect 280342 174664 280398 174720
rect 281538 171672 281594 171728
rect 280434 170176 280490 170232
rect 281538 169360 281594 169416
rect 281722 181328 281778 181384
rect 281814 168680 281870 168736
rect 282274 226888 282330 226944
rect 282182 202272 282238 202328
rect 282826 172488 282882 172544
rect 283010 218048 283066 218104
rect 282826 166404 282828 166424
rect 282828 166404 282880 166424
rect 282880 166404 282882 166424
rect 282826 166368 282882 166404
rect 282826 164872 282882 164928
rect 282826 164056 282882 164112
rect 282826 163240 282882 163296
rect 282826 162560 282882 162616
rect 282734 161744 282790 161800
rect 282826 161064 282882 161120
rect 282734 160248 282790 160304
rect 282550 159432 282606 159488
rect 282458 158752 282514 158808
rect 282090 157936 282146 157992
rect 281906 157256 281962 157312
rect 282182 154944 282238 155000
rect 282090 154128 282146 154184
rect 281722 152632 281778 152688
rect 281630 151816 281686 151872
rect 281538 148860 281540 148880
rect 281540 148860 281592 148880
rect 281592 148860 281594 148880
rect 281538 148824 281594 148860
rect 282826 155624 282882 155680
rect 282366 153448 282422 153504
rect 282826 151136 282882 151192
rect 282826 148008 282882 148064
rect 282826 147328 282882 147384
rect 282274 145016 282330 145072
rect 281906 144200 281962 144256
rect 282458 143520 282514 143576
rect 282090 142704 282146 142760
rect 283102 180104 283158 180160
rect 281906 142060 281908 142080
rect 281908 142060 281960 142080
rect 281960 142060 281962 142080
rect 281906 142024 281962 142060
rect 282274 141208 282330 141264
rect 281722 140392 281778 140448
rect 282274 139712 282330 139768
rect 282274 138896 282330 138952
rect 282826 138216 282882 138272
rect 281722 137400 281778 137456
rect 282826 136584 282882 136640
rect 281906 135904 281962 135960
rect 282090 134408 282146 134464
rect 282826 133592 282882 133648
rect 282274 132776 282330 132832
rect 282826 132096 282882 132152
rect 282734 131280 282790 131336
rect 282274 130600 282330 130656
rect 281538 129784 281594 129840
rect 282090 128968 282146 129024
rect 282826 128308 282882 128344
rect 282826 128288 282828 128308
rect 282828 128288 282880 128308
rect 282880 128288 282882 128308
rect 282734 127472 282790 127528
rect 282274 125976 282330 126032
rect 282090 125160 282146 125216
rect 282826 124480 282882 124536
rect 282274 123664 282330 123720
rect 282826 122984 282882 123040
rect 282458 122168 282514 122224
rect 282826 121388 282828 121408
rect 282828 121388 282880 121408
rect 282880 121388 282882 121408
rect 282826 121352 282882 121388
rect 282642 119856 282698 119912
rect 282090 119176 282146 119232
rect 281814 118396 281816 118416
rect 281816 118396 281868 118416
rect 281868 118396 281870 118416
rect 281814 118360 281870 118396
rect 280250 117544 280306 117600
rect 281998 112240 282054 112296
rect 281722 108432 281778 108488
rect 282826 116864 282882 116920
rect 282366 116048 282422 116104
rect 282826 115368 282882 115424
rect 282274 114552 282330 114608
rect 282826 113736 282882 113792
rect 282826 113092 282828 113112
rect 282828 113092 282880 113112
rect 282880 113092 282882 113112
rect 282826 113056 282882 113092
rect 282826 110744 282882 110800
rect 282274 109928 282330 109984
rect 282826 109248 282882 109304
rect 287242 233824 287298 233880
rect 298742 302232 298798 302288
rect 288438 287272 288494 287328
rect 282182 107752 282238 107808
rect 281998 103944 282054 104000
rect 281538 100816 281594 100872
rect 279422 98776 279478 98832
rect 267738 98232 267794 98288
rect 279330 98096 279386 98152
rect 269118 94832 269174 94888
rect 279330 95104 279386 95160
rect 280066 95784 280122 95840
rect 279422 94968 279478 95024
rect 281722 100136 281778 100192
rect 282826 105440 282882 105496
rect 282826 104624 282882 104680
rect 282826 103128 282882 103184
rect 288714 178880 288770 178936
rect 289910 210432 289966 210488
rect 290002 198056 290058 198112
rect 293958 187040 294014 187096
rect 292762 178744 292818 178800
rect 282734 102312 282790 102368
rect 282826 101632 282882 101688
rect 282274 97824 282330 97880
rect 281722 97008 281778 97064
rect 280066 93608 280122 93664
rect 277398 91704 277454 91760
rect 270498 84768 270554 84824
rect 273258 82184 273314 82240
rect 268382 14456 268438 14512
rect 266542 3576 266598 3632
rect 276018 65456 276074 65512
rect 280158 87488 280214 87544
rect 280802 22752 280858 22808
rect 274822 3440 274878 3496
rect 276018 3304 276074 3360
rect 284298 72392 284354 72448
rect 292578 37848 292634 37904
rect 286598 3440 286654 3496
rect 287794 3440 287850 3496
rect 288990 3440 289046 3496
rect 291382 3440 291438 3496
rect 298098 220088 298154 220144
rect 294878 3848 294934 3904
rect 299478 202136 299534 202192
rect 298374 177248 298430 177304
rect 300858 189896 300914 189952
rect 301134 204992 301190 205048
rect 302422 222944 302478 223000
rect 304262 284280 304318 284336
rect 303710 229744 303766 229800
rect 304262 211928 304318 211984
rect 298466 3984 298522 4040
rect 300766 3440 300822 3496
rect 305090 188264 305146 188320
rect 304906 3440 304962 3496
rect 305550 3440 305606 3496
rect 306470 218592 306526 218648
rect 307758 273264 307814 273320
rect 307850 237360 307906 237416
rect 307850 22616 307906 22672
rect 310518 285640 310574 285696
rect 309230 270544 309286 270600
rect 311898 199280 311954 199336
rect 313830 4800 313886 4856
rect 318062 306448 318118 306504
rect 316682 300872 316738 300928
rect 314658 282920 314714 282976
rect 316038 206352 316094 206408
rect 316130 195200 316186 195256
rect 317418 17176 317474 17232
rect 318798 190984 318854 191040
rect 324318 342216 324374 342272
rect 323582 322088 323638 322144
rect 322938 210296 322994 210352
rect 582378 365064 582434 365120
rect 331218 353368 331274 353424
rect 329838 185544 329894 185600
rect 580170 351872 580226 351928
rect 580170 349016 580226 349072
rect 357438 345072 357494 345128
rect 336002 340856 336058 340912
rect 333978 313928 334034 313984
rect 332690 196560 332746 196616
rect 335358 189624 335414 189680
rect 339498 338136 339554 338192
rect 338118 308352 338174 308408
rect 342258 217232 342314 217288
rect 340878 213152 340934 213208
rect 345018 207576 345074 207632
rect 347042 57160 347098 57216
rect 344558 3304 344614 3360
rect 356058 215872 356114 215928
rect 351918 211792 351974 211848
rect 351642 3576 351698 3632
rect 348054 3440 348110 3496
rect 353298 208936 353354 208992
rect 582378 343712 582434 343768
rect 574742 296792 574798 296848
rect 358818 197920 358874 197976
rect 579802 258848 579858 258904
rect 580170 245520 580226 245576
rect 580170 240080 580226 240136
rect 580170 219000 580226 219056
rect 580354 272176 580410 272232
rect 580262 192480 580318 192536
rect 580262 186904 580318 186960
rect 580170 179152 580226 179208
rect 580906 125976 580962 126032
rect 580262 59608 580318 59664
rect 582562 404912 582618 404968
rect 582470 291760 582526 291816
rect 582562 291080 582618 291136
rect 582746 378392 582802 378448
rect 582838 325216 582894 325272
rect 583022 312024 583078 312080
rect 582930 298152 582986 298208
rect 582654 232328 582710 232384
rect 582654 224984 582710 225040
rect 582470 86128 582526 86184
rect 358818 3576 358874 3632
rect 357438 3440 357494 3496
rect 356058 3304 356114 3360
rect 583114 299512 583170 299568
rect 582930 112784 582986 112840
rect 583390 298696 583446 298752
rect 583666 295296 583722 295352
rect 583482 237224 583538 237280
rect 583390 205672 583446 205728
rect 583390 204856 583446 204912
rect 583298 152632 583354 152688
rect 583114 139304 583170 139360
rect 583022 99456 583078 99512
rect 582838 46280 582894 46336
rect 582746 33088 582802 33144
rect 582654 6568 582710 6624
rect 583482 200640 583538 200696
rect 583574 166368 583630 166424
rect 583758 294480 583814 294536
rect 583758 73208 583814 73264
rect 583666 20304 583722 20360
<< metal3 >>
rect 69606 702476 69612 702540
rect 69676 702538 69682 702540
rect 154113 702538 154179 702541
rect 69676 702536 154179 702538
rect 69676 702480 154118 702536
rect 154174 702480 154179 702536
rect 69676 702478 154179 702480
rect 69676 702476 69682 702478
rect 154113 702475 154179 702478
rect 72969 699546 73035 699549
rect 76046 699546 76052 699548
rect 72969 699544 76052 699546
rect 72969 699488 72974 699544
rect 73030 699488 76052 699544
rect 72969 699486 76052 699488
rect 72969 699483 73035 699486
rect 76046 699484 76052 699486
rect 76116 699484 76122 699548
rect -960 697220 480 697460
rect 582373 697234 582439 697237
rect 583520 697234 584960 697324
rect 582373 697232 584960 697234
rect 582373 697176 582378 697232
rect 582434 697176 584960 697232
rect 582373 697174 584960 697176
rect 582373 697171 582439 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 582465 683906 582531 683909
rect 583520 683906 584960 683996
rect 582465 683904 584960 683906
rect 582465 683848 582470 683904
rect 582526 683848 584960 683904
rect 582465 683846 584960 683848
rect 582465 683843 582531 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580257 670714 580323 670717
rect 583520 670714 584960 670804
rect 580257 670712 584960 670714
rect 580257 670656 580262 670712
rect 580318 670656 584960 670712
rect 580257 670654 584960 670656
rect 580257 670651 580323 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 582557 644058 582623 644061
rect 583520 644058 584960 644148
rect 582557 644056 584960 644058
rect 582557 644000 582562 644056
rect 582618 644000 584960 644056
rect 582557 643998 584960 644000
rect 582557 643995 582623 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 582649 630866 582715 630869
rect 583520 630866 584960 630956
rect 582649 630864 584960 630866
rect 582649 630808 582654 630864
rect 582710 630808 584960 630864
rect 582649 630806 584960 630808
rect 582649 630803 582715 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 2773 619170 2839 619173
rect -960 619168 2839 619170
rect -960 619112 2778 619168
rect 2834 619112 2839 619168
rect -960 619110 2839 619112
rect -960 619020 480 619110
rect 2773 619107 2839 619110
rect 582741 617538 582807 617541
rect 583520 617538 584960 617628
rect 582741 617536 584960 617538
rect 582741 617480 582746 617536
rect 582802 617480 584960 617536
rect 582741 617478 584960 617480
rect 582741 617475 582807 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect 89161 593466 89227 593469
rect 582741 593466 582807 593469
rect 89161 593464 582807 593466
rect 89161 593408 89166 593464
rect 89222 593408 582746 593464
rect 582802 593408 582807 593464
rect 89161 593406 582807 593408
rect 89161 593403 89227 593406
rect 582741 593403 582807 593406
rect -960 592908 480 593148
rect 77937 592106 78003 592109
rect 98637 592106 98703 592109
rect 77937 592104 98703 592106
rect 77937 592048 77942 592104
rect 77998 592048 98642 592104
rect 98698 592048 98703 592104
rect 77937 592046 98703 592048
rect 77937 592043 78003 592046
rect 98637 592043 98703 592046
rect 83733 591970 83799 591973
rect 84326 591970 84332 591972
rect 83733 591968 84332 591970
rect 83733 591912 83738 591968
rect 83794 591912 84332 591968
rect 83733 591910 84332 591912
rect 83733 591907 83799 591910
rect 84326 591908 84332 591910
rect 84396 591908 84402 591972
rect 82537 591018 82603 591021
rect 107101 591018 107167 591021
rect 82537 591016 107167 591018
rect 82537 590960 82542 591016
rect 82598 590960 107106 591016
rect 107162 590960 107167 591016
rect 82537 590958 107167 590960
rect 82537 590955 82603 590958
rect 107101 590955 107167 590958
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 72417 590882 72483 590885
rect 84326 590882 84332 590884
rect 72417 590880 84332 590882
rect 72417 590824 72422 590880
rect 72478 590824 84332 590880
rect 72417 590822 84332 590824
rect 72417 590819 72483 590822
rect 84326 590820 84332 590822
rect 84396 590820 84402 590884
rect 86861 590882 86927 590885
rect 95877 590882 95943 590885
rect 86861 590880 95943 590882
rect 86861 590824 86866 590880
rect 86922 590824 95882 590880
rect 95938 590824 95943 590880
rect 583520 590868 584960 590958
rect 86861 590822 95943 590824
rect 86861 590819 86927 590822
rect 95877 590819 95943 590822
rect 52269 590746 52335 590749
rect 73613 590746 73679 590749
rect 52269 590744 73679 590746
rect 52269 590688 52274 590744
rect 52330 590688 73618 590744
rect 73674 590688 73679 590744
rect 52269 590686 73679 590688
rect 52269 590683 52335 590686
rect 73613 590683 73679 590686
rect 84101 590746 84167 590749
rect 88190 590746 88196 590748
rect 84101 590744 88196 590746
rect 84101 590688 84106 590744
rect 84162 590688 88196 590744
rect 84101 590686 88196 590688
rect 84101 590683 84167 590686
rect 88190 590684 88196 590686
rect 88260 590684 88266 590748
rect 73153 590066 73219 590069
rect 93894 590066 93900 590068
rect 73153 590064 93900 590066
rect 73153 590008 73158 590064
rect 73214 590008 93900 590064
rect 73153 590006 93900 590008
rect 73153 590003 73219 590006
rect 93894 590004 93900 590006
rect 93964 590004 93970 590068
rect 67725 589930 67791 589933
rect 580165 589930 580231 589933
rect 67725 589928 580231 589930
rect 67725 589872 67730 589928
rect 67786 589872 580170 589928
rect 580226 589872 580231 589928
rect 67725 589870 580231 589872
rect 67725 589867 67791 589870
rect 580165 589867 580231 589870
rect 75637 588842 75703 588845
rect 75637 588840 93870 588842
rect 75637 588784 75642 588840
rect 75698 588784 93870 588840
rect 75637 588782 93870 588784
rect 75637 588779 75703 588782
rect 84377 588708 84443 588709
rect 87873 588708 87939 588709
rect 84326 588706 84332 588708
rect 84286 588646 84332 588706
rect 84396 588704 84443 588708
rect 87822 588706 87828 588708
rect 84438 588648 84443 588704
rect 84326 588644 84332 588646
rect 84396 588644 84443 588648
rect 87782 588646 87828 588706
rect 87892 588704 87939 588708
rect 87934 588648 87939 588704
rect 87822 588644 87828 588646
rect 87892 588644 87939 588648
rect 93810 588706 93870 588782
rect 98729 588706 98795 588709
rect 93810 588704 98795 588706
rect 93810 588648 98734 588704
rect 98790 588648 98795 588704
rect 93810 588646 98795 588648
rect 84377 588643 84443 588644
rect 87873 588643 87939 588644
rect 98729 588643 98795 588646
rect 66805 588298 66871 588301
rect 68878 588298 68938 588472
rect 88885 588436 88951 588437
rect 88885 588432 88932 588436
rect 88996 588434 89002 588436
rect 88885 588376 88890 588432
rect 88885 588372 88932 588376
rect 88996 588374 89042 588434
rect 88996 588372 89002 588374
rect 88885 588371 88951 588372
rect 66805 588296 68938 588298
rect 66805 588240 66810 588296
rect 66866 588240 68938 588296
rect 66805 588238 68938 588240
rect 66805 588235 66871 588238
rect 66253 586530 66319 586533
rect 66253 586528 66362 586530
rect 66253 586472 66258 586528
rect 66314 586472 66362 586528
rect 66253 586467 66362 586472
rect 66302 586394 66362 586467
rect 68878 586394 68938 587112
rect 88566 586938 88626 587656
rect 88566 586878 96630 586938
rect 66302 586334 68938 586394
rect 96570 586394 96630 586878
rect 169702 586468 169708 586532
rect 169772 586468 169778 586532
rect 169710 586394 169770 586468
rect 96570 586334 169770 586394
rect 67725 585850 67791 585853
rect 67725 585848 68938 585850
rect 67725 585792 67730 585848
rect 67786 585792 68938 585848
rect 67725 585790 68938 585792
rect 67725 585787 67791 585790
rect 68878 585752 68938 585790
rect 88566 585714 88626 586296
rect 89897 585714 89963 585717
rect 88566 585712 89963 585714
rect 88566 585656 89902 585712
rect 89958 585656 89963 585712
rect 88566 585654 89963 585656
rect 89897 585651 89963 585654
rect 88190 585516 88196 585580
rect 88260 585578 88266 585580
rect 88260 585518 93870 585578
rect 88260 585516 88266 585518
rect 93810 585442 93870 585518
rect 112437 585442 112503 585445
rect 93810 585440 112503 585442
rect 93810 585384 112442 585440
rect 112498 585384 112503 585440
rect 93810 585382 112503 585384
rect 112437 585379 112503 585382
rect 88566 584626 88626 584936
rect 91921 584626 91987 584629
rect 88566 584624 91987 584626
rect 88566 584568 91926 584624
rect 91982 584568 91987 584624
rect 88566 584566 91987 584568
rect 91921 584563 91987 584566
rect 67725 583810 67791 583813
rect 68878 583810 68938 584392
rect 67725 583808 68938 583810
rect 67725 583752 67730 583808
rect 67786 583752 68938 583808
rect 67725 583750 68938 583752
rect 67725 583747 67791 583750
rect 91921 583674 91987 583677
rect 88566 583672 91987 583674
rect 88566 583616 91926 583672
rect 91982 583616 91987 583672
rect 88566 583614 91987 583616
rect 88566 583576 88626 583614
rect 91921 583611 91987 583614
rect 66805 582450 66871 582453
rect 68878 582450 68938 583032
rect 88926 582932 88932 582996
rect 88996 582994 89002 582996
rect 132493 582994 132559 582997
rect 88996 582992 132559 582994
rect 88996 582936 132498 582992
rect 132554 582936 132559 582992
rect 88996 582934 132559 582936
rect 88996 582932 89002 582934
rect 132493 582931 132559 582934
rect 66805 582448 68938 582450
rect 66805 582392 66810 582448
rect 66866 582392 68938 582448
rect 66805 582390 68938 582392
rect 66805 582387 66871 582390
rect 69422 582252 69428 582316
rect 69492 582252 69498 582316
rect 66989 581090 67055 581093
rect 69430 581090 69490 582252
rect 88566 581634 88626 582216
rect 91093 581634 91159 581637
rect 88566 581632 91159 581634
rect 88566 581576 91098 581632
rect 91154 581576 91159 581632
rect 88566 581574 91159 581576
rect 91093 581571 91159 581574
rect 93761 581634 93827 581637
rect 122598 581634 122604 581636
rect 93761 581632 122604 581634
rect 93761 581576 93766 581632
rect 93822 581576 122604 581632
rect 93761 581574 122604 581576
rect 93761 581571 93827 581574
rect 122598 581572 122604 581574
rect 122668 581572 122674 581636
rect 66989 581088 69490 581090
rect 66989 581032 66994 581088
rect 67050 581032 69490 581088
rect 66989 581030 69490 581032
rect 66989 581027 67055 581030
rect 97901 580954 97967 580957
rect 88566 580952 97967 580954
rect 88566 580896 97906 580952
rect 97962 580896 97967 580952
rect 88566 580894 97967 580896
rect 88566 580856 88626 580894
rect 97901 580891 97967 580894
rect -960 580002 480 580092
rect 3417 580002 3483 580005
rect -960 580000 3483 580002
rect -960 579944 3422 580000
rect 3478 579944 3483 580000
rect -960 579942 3483 579944
rect -960 579852 480 579942
rect 3417 579939 3483 579942
rect 66069 579730 66135 579733
rect 68878 579730 68938 580312
rect 97901 580274 97967 580277
rect 119470 580274 119476 580276
rect 97901 580272 119476 580274
rect 97901 580216 97906 580272
rect 97962 580216 119476 580272
rect 97901 580214 119476 580216
rect 97901 580211 97967 580214
rect 119470 580212 119476 580214
rect 119540 580212 119546 580276
rect 66069 579728 68938 579730
rect 66069 579672 66074 579728
rect 66130 579672 68938 579728
rect 66069 579670 68938 579672
rect 66069 579667 66135 579670
rect 67766 578308 67772 578372
rect 67836 578370 67842 578372
rect 68878 578370 68938 578952
rect 88566 578914 88626 579496
rect 91093 578914 91159 578917
rect 88566 578912 91159 578914
rect 88566 578856 91098 578912
rect 91154 578856 91159 578912
rect 88566 578854 91159 578856
rect 91093 578851 91159 578854
rect 67836 578310 68938 578370
rect 67836 578308 67842 578310
rect 67817 577010 67883 577013
rect 68878 577010 68938 577592
rect 88566 577554 88626 578136
rect 580257 577690 580323 577693
rect 583520 577690 584960 577780
rect 580257 577688 584960 577690
rect 580257 577632 580262 577688
rect 580318 577632 584960 577688
rect 580257 577630 584960 577632
rect 580257 577627 580323 577630
rect 91093 577554 91159 577557
rect 88566 577552 91159 577554
rect 88566 577496 91098 577552
rect 91154 577496 91159 577552
rect 583520 577540 584960 577630
rect 88566 577494 91159 577496
rect 91093 577491 91159 577494
rect 67817 577008 68938 577010
rect 67817 576952 67822 577008
rect 67878 576952 68938 577008
rect 67817 576950 68938 576952
rect 67817 576947 67883 576950
rect 88566 576738 88626 576776
rect 91185 576738 91251 576741
rect 88566 576736 91251 576738
rect 88566 576680 91190 576736
rect 91246 576680 91251 576736
rect 88566 576678 91251 576680
rect 91185 576675 91251 576678
rect 66897 575650 66963 575653
rect 68878 575650 68938 576232
rect 66897 575648 68938 575650
rect 66897 575592 66902 575648
rect 66958 575592 68938 575648
rect 66897 575590 68938 575592
rect 66897 575587 66963 575590
rect 67449 575378 67515 575381
rect 67449 575376 68938 575378
rect 67449 575320 67454 575376
rect 67510 575320 68938 575376
rect 67449 575318 68938 575320
rect 67449 575315 67515 575318
rect 68878 574872 68938 575318
rect 88566 574834 88626 575416
rect 91921 574834 91987 574837
rect 88566 574832 91987 574834
rect 88566 574776 91926 574832
rect 91982 574776 91987 574832
rect 88566 574774 91987 574776
rect 91921 574771 91987 574774
rect 66437 573202 66503 573205
rect 68878 573202 68938 573512
rect 88566 573474 88626 574056
rect 91093 573474 91159 573477
rect 88566 573472 91159 573474
rect 88566 573416 91098 573472
rect 91154 573416 91159 573472
rect 88566 573414 91159 573416
rect 91093 573411 91159 573414
rect 66437 573200 68938 573202
rect 66437 573144 66442 573200
rect 66498 573144 68938 573200
rect 66437 573142 68938 573144
rect 66437 573139 66503 573142
rect 66437 571842 66503 571845
rect 68878 571842 68938 572152
rect 88566 572114 88626 572696
rect 91185 572114 91251 572117
rect 88566 572112 91251 572114
rect 88566 572056 91190 572112
rect 91246 572056 91251 572112
rect 88566 572054 91251 572056
rect 91185 572051 91251 572054
rect 66437 571840 68938 571842
rect 66437 571784 66442 571840
rect 66498 571784 68938 571840
rect 66437 571782 68938 571784
rect 66437 571779 66503 571782
rect 91093 571434 91159 571437
rect 88566 571432 91159 571434
rect 88566 571376 91098 571432
rect 91154 571376 91159 571432
rect 88566 571374 91159 571376
rect 88566 571336 88626 571374
rect 91093 571371 91159 571374
rect 67265 570210 67331 570213
rect 68878 570210 68938 570792
rect 67265 570208 68938 570210
rect 67265 570152 67270 570208
rect 67326 570152 68938 570208
rect 67265 570150 68938 570152
rect 67265 570147 67331 570150
rect 91093 570074 91159 570077
rect 88566 570072 91159 570074
rect 88566 570016 91098 570072
rect 91154 570016 91159 570072
rect 88566 570014 91159 570016
rect 88566 569976 88626 570014
rect 91093 570011 91159 570014
rect 66805 568850 66871 568853
rect 68878 568850 68938 569432
rect 66805 568848 68938 568850
rect 66805 568792 66810 568848
rect 66866 568792 68938 568848
rect 66805 568790 68938 568792
rect 66805 568787 66871 568790
rect 91737 568714 91803 568717
rect 88566 568712 91803 568714
rect 88566 568656 91742 568712
rect 91798 568656 91803 568712
rect 88566 568654 91803 568656
rect 88566 568616 88626 568654
rect 91737 568651 91803 568654
rect 66897 567490 66963 567493
rect 68878 567490 68938 568072
rect 91277 567898 91343 567901
rect 66897 567488 68938 567490
rect 66897 567432 66902 567488
rect 66958 567432 68938 567488
rect 66897 567430 68938 567432
rect 88566 567896 91343 567898
rect 88566 567840 91282 567896
rect 91338 567840 91343 567896
rect 88566 567838 91343 567840
rect 66897 567427 66963 567430
rect 88566 567256 88626 567838
rect 91277 567835 91343 567838
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 67541 566810 67607 566813
rect 67541 566808 68938 566810
rect 67541 566752 67546 566808
rect 67602 566752 68938 566808
rect 67541 566750 68938 566752
rect 67541 566747 67607 566750
rect 68878 566712 68938 566750
rect 88566 565858 88626 565896
rect 91093 565858 91159 565861
rect 88566 565856 91159 565858
rect 88566 565800 91098 565856
rect 91154 565800 91159 565856
rect 88566 565798 91159 565800
rect 91093 565795 91159 565798
rect 66621 564634 66687 564637
rect 68878 564634 68938 565080
rect 66621 564632 68938 564634
rect 66621 564576 66626 564632
rect 66682 564576 68938 564632
rect 66621 564574 68938 564576
rect 66621 564571 66687 564574
rect 88566 564498 88626 564536
rect 91093 564498 91159 564501
rect 88566 564496 91159 564498
rect 88566 564440 91098 564496
rect 91154 564440 91159 564496
rect 88566 564438 91159 564440
rect 91093 564435 91159 564438
rect 582741 564362 582807 564365
rect 583520 564362 584960 564452
rect 582741 564360 584960 564362
rect 582741 564304 582746 564360
rect 582802 564304 584960 564360
rect 582741 564302 584960 564304
rect 582741 564299 582807 564302
rect 583520 564212 584960 564302
rect 66437 564090 66503 564093
rect 66437 564088 68938 564090
rect 66437 564032 66442 564088
rect 66498 564032 68938 564088
rect 66437 564030 68938 564032
rect 66437 564027 66503 564030
rect 68878 563720 68938 564030
rect 88566 563138 88626 563176
rect 91093 563138 91159 563141
rect 88566 563136 91159 563138
rect 88566 563080 91098 563136
rect 91154 563080 91159 563136
rect 88566 563078 91159 563080
rect 91093 563075 91159 563078
rect 66437 562050 66503 562053
rect 68878 562050 68938 562360
rect 66437 562048 68938 562050
rect 66437 561992 66442 562048
rect 66498 561992 68938 562048
rect 66437 561990 68938 561992
rect 66437 561987 66503 561990
rect 66621 560418 66687 560421
rect 68878 560418 68938 561000
rect 88566 560962 88626 561544
rect 91093 560962 91159 560965
rect 88566 560960 91159 560962
rect 88566 560904 91098 560960
rect 91154 560904 91159 560960
rect 88566 560902 91159 560904
rect 91093 560899 91159 560902
rect 66621 560416 68938 560418
rect 66621 560360 66626 560416
rect 66682 560360 68938 560416
rect 66621 560358 68938 560360
rect 66621 560355 66687 560358
rect 88566 560146 88626 560184
rect 89805 560146 89871 560149
rect 91829 560146 91895 560149
rect 88566 560144 91895 560146
rect 88566 560088 89810 560144
rect 89866 560088 91834 560144
rect 91890 560088 91895 560144
rect 88566 560086 91895 560088
rect 89805 560083 89871 560086
rect 91829 560083 91895 560086
rect 66621 559058 66687 559061
rect 68878 559058 68938 559640
rect 66621 559056 68938 559058
rect 66621 559000 66626 559056
rect 66682 559000 68938 559056
rect 66621 558998 68938 559000
rect 66621 558995 66687 558998
rect 67633 558922 67699 558925
rect 67633 558920 68938 558922
rect 67633 558864 67638 558920
rect 67694 558864 68938 558920
rect 67633 558862 68938 558864
rect 67633 558859 67699 558862
rect 68878 558280 68938 558862
rect 88566 558242 88626 558824
rect 91185 558242 91251 558245
rect 88566 558240 91251 558242
rect 88566 558184 91190 558240
rect 91246 558184 91251 558240
rect 88566 558182 91251 558184
rect 91185 558179 91251 558182
rect 67357 556338 67423 556341
rect 68878 556338 68938 556920
rect 88566 556882 88626 557464
rect 91185 556882 91251 556885
rect 88566 556880 91251 556882
rect 88566 556824 91190 556880
rect 91246 556824 91251 556880
rect 88566 556822 91251 556824
rect 91185 556819 91251 556822
rect 67357 556336 68938 556338
rect 67357 556280 67362 556336
rect 67418 556280 68938 556336
rect 67357 556278 68938 556280
rect 67357 556275 67423 556278
rect 66345 555250 66411 555253
rect 68878 555250 68938 555560
rect 88566 555522 88626 556104
rect 91185 555522 91251 555525
rect 88566 555520 91251 555522
rect 88566 555464 91190 555520
rect 91246 555464 91251 555520
rect 88566 555462 91251 555464
rect 91185 555459 91251 555462
rect 66345 555248 68938 555250
rect 66345 555192 66350 555248
rect 66406 555192 68938 555248
rect 66345 555190 68938 555192
rect 66345 555187 66411 555190
rect 66253 554706 66319 554709
rect 66253 554704 68938 554706
rect 66253 554648 66258 554704
rect 66314 554648 68938 554704
rect 66253 554646 68938 554648
rect 66253 554643 66319 554646
rect 68878 554200 68938 554646
rect 88566 554026 88626 554744
rect -960 553890 480 553980
rect 88566 553966 93870 554026
rect 3325 553890 3391 553893
rect -960 553888 3391 553890
rect -960 553832 3330 553888
rect 3386 553832 3391 553888
rect -960 553830 3391 553832
rect -960 553740 480 553830
rect 3325 553827 3391 553830
rect 93810 553482 93870 553966
rect 111006 553482 111012 553484
rect 93810 553422 111012 553482
rect 111006 553420 111012 553422
rect 111076 553420 111082 553484
rect 67449 552258 67515 552261
rect 68878 552258 68938 552840
rect 88566 552802 88626 553384
rect 91277 552802 91343 552805
rect 88566 552800 91343 552802
rect 88566 552744 91282 552800
rect 91338 552744 91343 552800
rect 88566 552742 91343 552744
rect 91277 552739 91343 552742
rect 67449 552256 68938 552258
rect 67449 552200 67454 552256
rect 67510 552200 68938 552256
rect 67449 552198 68938 552200
rect 67449 552195 67515 552198
rect 91185 552122 91251 552125
rect 88566 552120 91251 552122
rect 88566 552064 91190 552120
rect 91246 552064 91251 552120
rect 88566 552062 91251 552064
rect 88566 552024 88626 552062
rect 91185 552059 91251 552062
rect 66662 550836 66668 550900
rect 66732 550898 66738 550900
rect 68878 550898 68938 551480
rect 583520 551020 584960 551260
rect 66732 550838 68938 550898
rect 66732 550836 66738 550838
rect 99966 550762 99972 550764
rect 88566 550702 99972 550762
rect 88566 550664 88626 550702
rect 99966 550700 99972 550702
rect 100036 550700 100042 550764
rect 66529 549674 66595 549677
rect 68878 549674 68938 550120
rect 66529 549672 68938 549674
rect 66529 549616 66534 549672
rect 66590 549616 68938 549672
rect 66529 549614 68938 549616
rect 66529 549611 66595 549614
rect 91185 549402 91251 549405
rect 88566 549400 91251 549402
rect 88566 549344 91190 549400
rect 91246 549344 91251 549400
rect 88566 549342 91251 549344
rect 88566 549304 88626 549342
rect 91185 549339 91251 549342
rect 66529 548314 66595 548317
rect 68878 548314 68938 548760
rect 66529 548312 68938 548314
rect 66529 548256 66534 548312
rect 66590 548256 68938 548312
rect 66529 548254 68938 548256
rect 66529 548251 66595 548254
rect 88566 547906 88626 547944
rect 91185 547906 91251 547909
rect 88566 547904 91251 547906
rect 88566 547848 91190 547904
rect 91246 547848 91251 547904
rect 88566 547846 91251 547848
rect 91185 547843 91251 547846
rect 66805 547634 66871 547637
rect 66805 547632 68938 547634
rect 66805 547576 66810 547632
rect 66866 547576 68938 547632
rect 66805 547574 68938 547576
rect 66805 547571 66871 547574
rect 68878 547400 68938 547574
rect 88566 546546 88626 546584
rect 91277 546546 91343 546549
rect 88566 546544 91343 546546
rect 88566 546488 91282 546544
rect 91338 546488 91343 546544
rect 88566 546486 91343 546488
rect 91277 546483 91343 546486
rect 66161 546410 66227 546413
rect 66161 546408 68938 546410
rect 66161 546352 66166 546408
rect 66222 546352 68938 546408
rect 66161 546350 68938 546352
rect 66161 546347 66227 546350
rect 68878 546040 68938 546350
rect 91277 545458 91343 545461
rect 88566 545456 91343 545458
rect 88566 545400 91282 545456
rect 91338 545400 91343 545456
rect 88566 545398 91343 545400
rect 88566 545224 88626 545398
rect 91277 545395 91343 545398
rect 66805 544914 66871 544917
rect 66805 544912 68938 544914
rect 66805 544856 66810 544912
rect 66866 544856 68938 544912
rect 66805 544854 68938 544856
rect 66805 544851 66871 544854
rect 68878 544680 68938 544854
rect 91277 544098 91343 544101
rect 88566 544096 91343 544098
rect 88566 544040 91282 544096
rect 91338 544040 91343 544096
rect 88566 544038 91343 544040
rect 88566 543864 88626 544038
rect 91277 544035 91343 544038
rect 66805 542738 66871 542741
rect 68878 542738 68938 543320
rect 66805 542736 68938 542738
rect 66805 542680 66810 542736
rect 66866 542680 68938 542736
rect 66805 542678 68938 542680
rect 66805 542675 66871 542678
rect 88566 542466 88626 542504
rect 91277 542466 91343 542469
rect 88566 542464 91343 542466
rect 88566 542408 91282 542464
rect 91338 542408 91343 542464
rect 88566 542406 91343 542408
rect 91277 542403 91343 542406
rect 67081 541786 67147 541789
rect 68878 541786 68938 541960
rect 67081 541784 68938 541786
rect 67081 541728 67086 541784
rect 67142 541728 68938 541784
rect 67081 541726 68938 541728
rect 67081 541723 67147 541726
rect 91277 541378 91343 541381
rect 88566 541376 91343 541378
rect 88566 541320 91282 541376
rect 91338 541320 91343 541376
rect 88566 541318 91343 541320
rect 88566 541144 88626 541318
rect 91277 541315 91343 541318
rect -960 540684 480 540924
rect 68645 540834 68711 540837
rect 68645 540832 68938 540834
rect 68645 540776 68650 540832
rect 68706 540776 68938 540832
rect 68645 540774 68938 540776
rect 68645 540771 68711 540774
rect 68878 540600 68938 540774
rect 88566 539746 88626 539784
rect 91277 539746 91343 539749
rect 88566 539744 91343 539746
rect 88566 539688 91282 539744
rect 91338 539688 91343 539744
rect 88566 539686 91343 539688
rect 91277 539683 91343 539686
rect 76046 538052 76052 538116
rect 76116 538114 76122 538116
rect 76741 538114 76807 538117
rect 76116 538112 76807 538114
rect 76116 538056 76746 538112
rect 76802 538056 76807 538112
rect 76116 538054 76807 538056
rect 76116 538052 76122 538054
rect 76741 538051 76807 538054
rect 579797 537842 579863 537845
rect 583520 537842 584960 537932
rect 579797 537840 584960 537842
rect 579797 537784 579802 537840
rect 579858 537784 584960 537840
rect 579797 537782 584960 537784
rect 579797 537779 579863 537782
rect 583520 537692 584960 537782
rect 82721 536754 82787 536757
rect 130377 536754 130443 536757
rect 82721 536752 130443 536754
rect 82721 536696 82726 536752
rect 82782 536696 130382 536752
rect 130438 536696 130443 536752
rect 82721 536694 130443 536696
rect 82721 536691 82787 536694
rect 130377 536691 130443 536694
rect 84745 536074 84811 536077
rect 128997 536074 129063 536077
rect 582373 536074 582439 536077
rect 84745 536072 582439 536074
rect 84745 536016 84750 536072
rect 84806 536016 129002 536072
rect 129058 536016 582378 536072
rect 582434 536016 582439 536072
rect 84745 536014 582439 536016
rect 84745 536011 84811 536014
rect 128997 536011 129063 536014
rect 582373 536011 582439 536014
rect 68134 535468 68140 535532
rect 68204 535530 68210 535532
rect 68461 535530 68527 535533
rect 69657 535532 69723 535533
rect 69606 535530 69612 535532
rect 68204 535528 68527 535530
rect 68204 535472 68466 535528
rect 68522 535472 68527 535528
rect 68204 535470 68527 535472
rect 69566 535470 69612 535530
rect 69676 535528 69723 535532
rect 69718 535472 69723 535528
rect 68204 535468 68210 535470
rect 68461 535467 68527 535470
rect 69606 535468 69612 535470
rect 69676 535468 69723 535472
rect 69657 535467 69723 535468
rect 70669 535530 70735 535533
rect 71814 535530 71820 535532
rect 70669 535528 71820 535530
rect 70669 535472 70674 535528
rect 70730 535472 71820 535528
rect 70669 535470 71820 535472
rect 70669 535467 70735 535470
rect 71814 535468 71820 535470
rect 71884 535468 71890 535532
rect 75913 535530 75979 535533
rect 76741 535530 76807 535533
rect 75913 535528 76807 535530
rect 75913 535472 75918 535528
rect 75974 535472 76746 535528
rect 76802 535472 76807 535528
rect 75913 535470 76807 535472
rect 75913 535467 75979 535470
rect 76741 535467 76807 535470
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 582465 524514 582531 524517
rect 583520 524514 584960 524604
rect 582465 524512 584960 524514
rect 582465 524456 582470 524512
rect 582526 524456 584960 524512
rect 582465 524454 584960 524456
rect 582465 524451 582531 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3509 514858 3575 514861
rect -960 514856 3575 514858
rect -960 514800 3514 514856
rect 3570 514800 3575 514856
rect -960 514798 3575 514800
rect -960 514708 480 514798
rect 3509 514795 3575 514798
rect 93117 512682 93183 512685
rect 102174 512682 102180 512684
rect 93117 512680 102180 512682
rect 93117 512624 93122 512680
rect 93178 512624 102180 512680
rect 93117 512622 102180 512624
rect 93117 512619 93183 512622
rect 102174 512620 102180 512622
rect 102244 512620 102250 512684
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3325 501802 3391 501805
rect -960 501800 3391 501802
rect -960 501744 3330 501800
rect 3386 501744 3391 501800
rect -960 501742 3391 501744
rect -960 501652 480 501742
rect 3325 501739 3391 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 582373 484666 582439 484669
rect 583520 484666 584960 484756
rect 582373 484664 584960 484666
rect 582373 484608 582378 484664
rect 582434 484608 584960 484664
rect 582373 484606 584960 484608
rect 582373 484603 582439 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 4061 475690 4127 475693
rect -960 475688 4127 475690
rect -960 475632 4066 475688
rect 4122 475632 4127 475688
rect -960 475630 4127 475632
rect -960 475540 480 475630
rect 4061 475627 4127 475630
rect 582649 471474 582715 471477
rect 583520 471474 584960 471564
rect 582649 471472 584960 471474
rect 582649 471416 582654 471472
rect 582710 471416 584960 471472
rect 582649 471414 584960 471416
rect 582649 471411 582715 471414
rect 583520 471324 584960 471414
rect 67766 467740 67772 467804
rect 67836 467802 67842 467804
rect 76557 467802 76623 467805
rect 67836 467800 76623 467802
rect 67836 467744 76562 467800
rect 76618 467744 76623 467800
rect 67836 467742 76623 467744
rect 67836 467740 67842 467742
rect 76557 467739 76623 467742
rect 96429 467122 96495 467125
rect 107694 467122 107700 467124
rect 96429 467120 107700 467122
rect 96429 467064 96434 467120
rect 96490 467064 107700 467120
rect 96429 467062 107700 467064
rect 96429 467059 96495 467062
rect 107694 467060 107700 467062
rect 107764 467060 107770 467124
rect 96521 464402 96587 464405
rect 106406 464402 106412 464404
rect 96521 464400 106412 464402
rect 96521 464344 96526 464400
rect 96582 464344 106412 464400
rect 96521 464342 106412 464344
rect 96521 464339 96587 464342
rect 106406 464340 106412 464342
rect 106476 464340 106482 464404
rect 104249 463586 104315 463589
rect 111742 463586 111748 463588
rect 104249 463584 111748 463586
rect 104249 463528 104254 463584
rect 104310 463528 111748 463584
rect 104249 463526 111748 463528
rect 104249 463523 104315 463526
rect 111742 463524 111748 463526
rect 111812 463524 111818 463588
rect 81433 462906 81499 462909
rect 89662 462906 89668 462908
rect 81433 462904 89668 462906
rect 81433 462848 81438 462904
rect 81494 462848 89668 462904
rect 81433 462846 89668 462848
rect 81433 462843 81499 462846
rect 89662 462844 89668 462846
rect 89732 462844 89738 462908
rect -960 462634 480 462724
rect 2773 462634 2839 462637
rect -960 462632 2839 462634
rect -960 462576 2778 462632
rect 2834 462576 2839 462632
rect -960 462574 2839 462576
rect -960 462484 480 462574
rect 2773 462571 2839 462574
rect 86953 461546 87019 461549
rect 98126 461546 98132 461548
rect 86953 461544 98132 461546
rect 86953 461488 86958 461544
rect 87014 461488 98132 461544
rect 86953 461486 98132 461488
rect 86953 461483 87019 461486
rect 98126 461484 98132 461486
rect 98196 461484 98202 461548
rect 107009 461546 107075 461549
rect 115974 461546 115980 461548
rect 107009 461544 115980 461546
rect 107009 461488 107014 461544
rect 107070 461488 115980 461544
rect 107009 461486 115980 461488
rect 107009 461483 107075 461486
rect 115974 461484 115980 461486
rect 116044 461484 116050 461548
rect 88190 460124 88196 460188
rect 88260 460186 88266 460188
rect 118693 460186 118759 460189
rect 88260 460184 118759 460186
rect 88260 460128 118698 460184
rect 118754 460128 118759 460184
rect 88260 460126 118759 460128
rect 88260 460124 88266 460126
rect 118693 460123 118759 460126
rect 104157 458282 104223 458285
rect 109166 458282 109172 458284
rect 104157 458280 109172 458282
rect 104157 458224 104162 458280
rect 104218 458224 109172 458280
rect 104157 458222 109172 458224
rect 104157 458219 104223 458222
rect 109166 458220 109172 458222
rect 109236 458220 109242 458284
rect 97257 458146 97323 458149
rect 104934 458146 104940 458148
rect 97257 458144 104940 458146
rect 97257 458088 97262 458144
rect 97318 458088 104940 458144
rect 97257 458086 104940 458088
rect 97257 458083 97323 458086
rect 104934 458084 104940 458086
rect 105004 458084 105010 458148
rect 582465 458146 582531 458149
rect 583520 458146 584960 458236
rect 582465 458144 584960 458146
rect 582465 458088 582470 458144
rect 582526 458088 584960 458144
rect 582465 458086 584960 458088
rect 582465 458083 582531 458086
rect 583520 457996 584960 458086
rect 86861 457466 86927 457469
rect 96654 457466 96660 457468
rect 86861 457464 96660 457466
rect 86861 457408 86866 457464
rect 86922 457408 96660 457464
rect 86861 457406 96660 457408
rect 86861 457403 86927 457406
rect 96654 457404 96660 457406
rect 96724 457404 96730 457468
rect 88333 456106 88399 456109
rect 100702 456106 100708 456108
rect 88333 456104 100708 456106
rect 88333 456048 88338 456104
rect 88394 456048 100708 456104
rect 88333 456046 100708 456048
rect 88333 456043 88399 456046
rect 100702 456044 100708 456046
rect 100772 456044 100778 456108
rect 84101 454746 84167 454749
rect 92790 454746 92796 454748
rect 84101 454744 92796 454746
rect 84101 454688 84106 454744
rect 84162 454688 92796 454744
rect 84101 454686 92796 454688
rect 84101 454683 84167 454686
rect 92790 454684 92796 454686
rect 92860 454684 92866 454748
rect 82721 453250 82787 453253
rect 91134 453250 91140 453252
rect 82721 453248 91140 453250
rect 82721 453192 82726 453248
rect 82782 453192 91140 453248
rect 82721 453190 91140 453192
rect 82721 453187 82787 453190
rect 91134 453188 91140 453190
rect 91204 453188 91210 453252
rect 83457 451346 83523 451349
rect 160134 451346 160140 451348
rect 83457 451344 160140 451346
rect 83457 451288 83462 451344
rect 83518 451288 160140 451344
rect 83457 451286 160140 451288
rect 83457 451283 83523 451286
rect 160134 451284 160140 451286
rect 160204 451284 160210 451348
rect 108297 449986 108363 449989
rect 132534 449986 132540 449988
rect 108297 449984 132540 449986
rect 108297 449928 108302 449984
rect 108358 449928 132540 449984
rect 108297 449926 132540 449928
rect 108297 449923 108363 449926
rect 132534 449924 132540 449926
rect 132604 449924 132610 449988
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 41321 449170 41387 449173
rect 70301 449170 70367 449173
rect 41321 449168 74550 449170
rect 41321 449112 41326 449168
rect 41382 449112 70306 449168
rect 70362 449112 74550 449168
rect 41321 449110 74550 449112
rect 41321 449107 41387 449110
rect 70301 449107 70367 449110
rect 74490 448626 74550 449110
rect 142797 448626 142863 448629
rect 74490 448624 142863 448626
rect 74490 448568 142802 448624
rect 142858 448568 142863 448624
rect 74490 448566 142863 448568
rect 142797 448563 142863 448566
rect 108941 447946 109007 447949
rect 120022 447946 120028 447948
rect 108941 447944 120028 447946
rect 108941 447888 108946 447944
rect 109002 447888 120028 447944
rect 108941 447886 120028 447888
rect 108941 447883 109007 447886
rect 120022 447884 120028 447886
rect 120092 447884 120098 447948
rect 65977 447810 66043 447813
rect 78765 447810 78831 447813
rect 65977 447808 78831 447810
rect 65977 447752 65982 447808
rect 66038 447752 78770 447808
rect 78826 447752 78831 447808
rect 65977 447750 78831 447752
rect 65977 447747 66043 447750
rect 78765 447747 78831 447750
rect 86217 447810 86283 447813
rect 95182 447810 95188 447812
rect 86217 447808 95188 447810
rect 86217 447752 86222 447808
rect 86278 447752 95188 447808
rect 86217 447750 95188 447752
rect 86217 447747 86283 447750
rect 95182 447748 95188 447750
rect 95252 447748 95258 447812
rect 100661 447810 100727 447813
rect 122966 447810 122972 447812
rect 100661 447808 122972 447810
rect 100661 447752 100666 447808
rect 100722 447752 122972 447808
rect 100661 447750 122972 447752
rect 100661 447747 100727 447750
rect 122966 447748 122972 447750
rect 123036 447748 123042 447812
rect 59169 445906 59235 445909
rect 85573 445906 85639 445909
rect 59169 445904 85639 445906
rect 59169 445848 59174 445904
rect 59230 445848 85578 445904
rect 85634 445848 85639 445904
rect 59169 445846 85639 445848
rect 59169 445843 59235 445846
rect 85573 445843 85639 445846
rect 105537 445906 105603 445909
rect 191097 445906 191163 445909
rect 105537 445904 191163 445906
rect 105537 445848 105542 445904
rect 105598 445848 191102 445904
rect 191158 445848 191163 445904
rect 105537 445846 191163 445848
rect 105537 445843 105603 445846
rect 191097 445843 191163 445846
rect 88793 445770 88859 445773
rect 92606 445770 92612 445772
rect 88793 445768 92612 445770
rect 88793 445712 88798 445768
rect 88854 445712 92612 445768
rect 88793 445710 92612 445712
rect 88793 445707 88859 445710
rect 92606 445708 92612 445710
rect 92676 445708 92682 445772
rect 93894 445708 93900 445772
rect 93964 445770 93970 445772
rect 94405 445770 94471 445773
rect 93964 445768 94471 445770
rect 93964 445712 94410 445768
rect 94466 445712 94471 445768
rect 93964 445710 94471 445712
rect 93964 445708 93970 445710
rect 94405 445707 94471 445710
rect 96470 445708 96476 445772
rect 96540 445770 96546 445772
rect 96613 445770 96679 445773
rect 97349 445770 97415 445773
rect 96540 445768 97415 445770
rect 96540 445712 96618 445768
rect 96674 445712 97354 445768
rect 97410 445712 97415 445768
rect 96540 445710 97415 445712
rect 96540 445708 96546 445710
rect 96613 445707 96679 445710
rect 97349 445707 97415 445710
rect 98637 445770 98703 445773
rect 102133 445770 102199 445773
rect 102358 445770 102364 445772
rect 98637 445768 102364 445770
rect 98637 445712 98642 445768
rect 98698 445712 102138 445768
rect 102194 445712 102364 445768
rect 98637 445710 102364 445712
rect 98637 445707 98703 445710
rect 102133 445707 102199 445710
rect 102358 445708 102364 445710
rect 102428 445708 102434 445772
rect 110413 445770 110479 445773
rect 111425 445770 111491 445773
rect 111558 445770 111564 445772
rect 110413 445768 111564 445770
rect 110413 445712 110418 445768
rect 110474 445712 111430 445768
rect 111486 445712 111564 445768
rect 110413 445710 111564 445712
rect 110413 445707 110479 445710
rect 111425 445707 111491 445710
rect 111558 445708 111564 445710
rect 111628 445708 111634 445772
rect 117313 445770 117379 445773
rect 118550 445770 118556 445772
rect 117313 445768 118556 445770
rect 117313 445712 117318 445768
rect 117374 445712 118556 445768
rect 117313 445710 118556 445712
rect 117313 445707 117379 445710
rect 118550 445708 118556 445710
rect 118620 445708 118626 445772
rect 68737 444818 68803 444821
rect 68870 444818 68876 444820
rect 68737 444816 68876 444818
rect 68737 444760 68742 444816
rect 68798 444760 68876 444816
rect 68737 444758 68876 444760
rect 68737 444755 68803 444758
rect 68870 444756 68876 444758
rect 68940 444756 68946 444820
rect 114318 444756 114324 444820
rect 114388 444818 114394 444820
rect 114461 444818 114527 444821
rect 114388 444816 114527 444818
rect 114388 444760 114466 444816
rect 114522 444760 114527 444816
rect 114388 444758 114527 444760
rect 114388 444756 114394 444758
rect 114461 444755 114527 444758
rect 109493 444684 109559 444685
rect 109493 444680 109540 444684
rect 109604 444682 109610 444684
rect 119015 444682 119081 444685
rect 143574 444682 143580 444684
rect 109493 444624 109498 444680
rect 109493 444620 109540 444624
rect 109604 444622 109650 444682
rect 119015 444680 143580 444682
rect 119015 444624 119020 444680
rect 119076 444624 143580 444680
rect 119015 444622 143580 444624
rect 109604 444620 109610 444622
rect 109493 444619 109559 444620
rect 119015 444619 119081 444622
rect 143574 444620 143580 444622
rect 143644 444620 143650 444684
rect 583520 444668 584960 444908
rect 90127 444546 90193 444549
rect 137277 444546 137343 444549
rect 90127 444544 137343 444546
rect 90127 444488 90132 444544
rect 90188 444488 137282 444544
rect 137338 444488 137343 444544
rect 90127 444486 137343 444488
rect 90127 444483 90193 444486
rect 137277 444483 137343 444486
rect 124121 444274 124187 444277
rect 120612 444272 124187 444274
rect 120612 444216 124126 444272
rect 124182 444216 124187 444272
rect 120612 444214 124187 444216
rect 124121 444211 124187 444214
rect 67725 442098 67791 442101
rect 124121 442098 124187 442101
rect 67725 442096 68908 442098
rect 67725 442040 67730 442096
rect 67786 442040 68908 442096
rect 67725 442038 68908 442040
rect 120612 442096 124187 442098
rect 120612 442040 124126 442096
rect 124182 442040 124187 442096
rect 120612 442038 124187 442040
rect 67725 442035 67791 442038
rect 124121 442035 124187 442038
rect 66989 439922 67055 439925
rect 120809 439922 120875 439925
rect 124121 439922 124187 439925
rect 66989 439920 68908 439922
rect 66989 439864 66994 439920
rect 67050 439864 68908 439920
rect 66989 439862 68908 439864
rect 120612 439920 124187 439922
rect 120612 439864 120814 439920
rect 120870 439864 124126 439920
rect 124182 439864 124187 439920
rect 120612 439862 124187 439864
rect 66989 439859 67055 439862
rect 120809 439859 120875 439862
rect 124121 439859 124187 439862
rect 66805 437746 66871 437749
rect 124121 437746 124187 437749
rect 66805 437744 68908 437746
rect 66805 437688 66810 437744
rect 66866 437688 68908 437744
rect 66805 437686 68908 437688
rect 120612 437744 124187 437746
rect 120612 437688 124126 437744
rect 124182 437688 124187 437744
rect 120612 437686 124187 437688
rect 66805 437683 66871 437686
rect 124121 437683 124187 437686
rect -960 436508 480 436748
rect 122598 435842 122604 435844
rect 120582 435782 122604 435842
rect 66805 435298 66871 435301
rect 120582 435298 120642 435782
rect 122598 435780 122604 435782
rect 122668 435780 122674 435844
rect 120809 435298 120875 435301
rect 66805 435296 68908 435298
rect 66805 435240 66810 435296
rect 66866 435240 68908 435296
rect 120582 435296 120875 435298
rect 120582 435268 120814 435296
rect 66805 435238 68908 435240
rect 120612 435240 120814 435268
rect 120870 435240 120875 435296
rect 120612 435238 120875 435240
rect 66805 435235 66871 435238
rect 120809 435235 120875 435238
rect 66897 433122 66963 433125
rect 122925 433122 122991 433125
rect 124121 433122 124187 433125
rect 66897 433120 68908 433122
rect 66897 433064 66902 433120
rect 66958 433064 68908 433120
rect 66897 433062 68908 433064
rect 120612 433120 124187 433122
rect 120612 433064 122930 433120
rect 122986 433064 124126 433120
rect 124182 433064 124187 433120
rect 120612 433062 124187 433064
rect 66897 433059 66963 433062
rect 122925 433059 122991 433062
rect 124121 433059 124187 433062
rect 582373 431626 582439 431629
rect 583520 431626 584960 431716
rect 582373 431624 584960 431626
rect 582373 431568 582378 431624
rect 582434 431568 584960 431624
rect 582373 431566 584960 431568
rect 582373 431563 582439 431566
rect 120022 431428 120028 431492
rect 120092 431428 120098 431492
rect 583520 431476 584960 431566
rect 66897 430946 66963 430949
rect 120030 430946 120090 431428
rect 122598 430946 122604 430948
rect 66897 430944 68908 430946
rect 66897 430888 66902 430944
rect 66958 430888 68908 430944
rect 120030 430916 122604 430946
rect 66897 430886 68908 430888
rect 120060 430886 122604 430916
rect 66897 430883 66963 430886
rect 122598 430884 122604 430886
rect 122668 430884 122674 430948
rect 66805 428498 66871 428501
rect 121545 428498 121611 428501
rect 122833 428498 122899 428501
rect 66805 428496 68908 428498
rect 66805 428440 66810 428496
rect 66866 428440 68908 428496
rect 66805 428438 68908 428440
rect 120612 428496 122899 428498
rect 120612 428440 121550 428496
rect 121606 428440 122838 428496
rect 122894 428440 122899 428496
rect 120612 428438 122899 428440
rect 66805 428435 66871 428438
rect 121545 428435 121611 428438
rect 122833 428435 122899 428438
rect 66253 426322 66319 426325
rect 122966 426322 122972 426324
rect 66253 426320 68908 426322
rect 66253 426264 66258 426320
rect 66314 426264 68908 426320
rect 66253 426262 68908 426264
rect 120612 426262 122972 426322
rect 66253 426259 66319 426262
rect 122966 426260 122972 426262
rect 123036 426260 123042 426324
rect 66253 424146 66319 424149
rect 123017 424146 123083 424149
rect 66253 424144 68908 424146
rect 66253 424088 66258 424144
rect 66314 424088 68908 424144
rect 66253 424086 68908 424088
rect 120612 424144 123083 424146
rect 120612 424088 123022 424144
rect 123078 424088 123083 424144
rect 120612 424086 123083 424088
rect 66253 424083 66319 424086
rect 123017 424083 123083 424086
rect -960 423602 480 423692
rect 3141 423602 3207 423605
rect -960 423600 3207 423602
rect -960 423544 3146 423600
rect 3202 423544 3207 423600
rect -960 423542 3207 423544
rect -960 423452 480 423542
rect 3141 423539 3207 423542
rect 66253 421970 66319 421973
rect 123017 421970 123083 421973
rect 66253 421968 68908 421970
rect 66253 421912 66258 421968
rect 66314 421912 68908 421968
rect 66253 421910 68908 421912
rect 120612 421968 123083 421970
rect 120612 421912 123022 421968
rect 123078 421912 123083 421968
rect 120612 421910 123083 421912
rect 66253 421907 66319 421910
rect 123017 421907 123083 421910
rect 67357 419522 67423 419525
rect 67357 419520 69276 419522
rect 67357 419464 67362 419520
rect 67418 419492 69276 419520
rect 67418 419464 69306 419492
rect 67357 419462 69306 419464
rect 67357 419459 67423 419462
rect 69246 419388 69306 419462
rect 69238 419324 69244 419388
rect 69308 419324 69314 419388
rect 120582 418978 120642 419492
rect 120717 418978 120783 418981
rect 120582 418976 120783 418978
rect 120582 418920 120722 418976
rect 120778 418920 120783 418976
rect 120582 418918 120783 418920
rect 120717 418915 120783 418918
rect 582465 418298 582531 418301
rect 583520 418298 584960 418388
rect 582465 418296 584960 418298
rect 582465 418240 582470 418296
rect 582526 418240 584960 418296
rect 582465 418238 584960 418240
rect 582465 418235 582531 418238
rect 583520 418148 584960 418238
rect 66897 417346 66963 417349
rect 121545 417346 121611 417349
rect 66897 417344 68908 417346
rect 66897 417288 66902 417344
rect 66958 417288 68908 417344
rect 66897 417286 68908 417288
rect 120612 417344 121611 417346
rect 120612 417288 121550 417344
rect 121606 417288 121611 417344
rect 120612 417286 121611 417288
rect 66897 417283 66963 417286
rect 121545 417283 121611 417286
rect 66437 415170 66503 415173
rect 124121 415170 124187 415173
rect 66437 415168 68908 415170
rect 66437 415112 66442 415168
rect 66498 415112 68908 415168
rect 66437 415110 68908 415112
rect 120612 415168 124187 415170
rect 120612 415112 124126 415168
rect 124182 415112 124187 415168
rect 120612 415110 124187 415112
rect 66437 415107 66503 415110
rect 124121 415107 124187 415110
rect 67449 412722 67515 412725
rect 123109 412722 123175 412725
rect 67449 412720 68908 412722
rect 67449 412664 67454 412720
rect 67510 412664 68908 412720
rect 67449 412662 68908 412664
rect 120612 412720 123175 412722
rect 120612 412664 123114 412720
rect 123170 412664 123175 412720
rect 120612 412662 123175 412664
rect 67449 412659 67515 412662
rect 123109 412659 123175 412662
rect 59261 411362 59327 411365
rect 66662 411362 66668 411364
rect 59261 411360 66668 411362
rect 59261 411304 59266 411360
rect 59322 411304 66668 411360
rect 59261 411302 66668 411304
rect 59261 411299 59327 411302
rect 66662 411300 66668 411302
rect 66732 411362 66738 411364
rect 66732 411302 66914 411362
rect 66732 411300 66738 411302
rect 66854 411226 66914 411302
rect 66854 411166 68938 411226
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect 68878 410516 68938 411166
rect 121637 410546 121703 410549
rect 120612 410544 121703 410546
rect -960 410486 3483 410488
rect 120612 410488 121642 410544
rect 121698 410488 121703 410544
rect 120612 410486 121703 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 121637 410483 121703 410486
rect 66529 408370 66595 408373
rect 124121 408370 124187 408373
rect 66529 408368 68908 408370
rect 66529 408312 66534 408368
rect 66590 408312 68908 408368
rect 66529 408310 68908 408312
rect 120612 408368 124187 408370
rect 120612 408312 124126 408368
rect 124182 408312 124187 408368
rect 120612 408310 124187 408312
rect 66529 408307 66595 408310
rect 124121 408307 124187 408310
rect 124949 406330 125015 406333
rect 146886 406330 146892 406332
rect 124949 406328 146892 406330
rect 124949 406272 124954 406328
rect 125010 406272 146892 406328
rect 124949 406270 146892 406272
rect 124949 406267 125015 406270
rect 146886 406268 146892 406270
rect 146956 406268 146962 406332
rect 66621 406194 66687 406197
rect 123201 406194 123267 406197
rect 66621 406192 68908 406194
rect 66621 406136 66626 406192
rect 66682 406136 68908 406192
rect 66621 406134 68908 406136
rect 120612 406192 123267 406194
rect 120612 406136 123206 406192
rect 123262 406136 123267 406192
rect 120612 406134 123267 406136
rect 66621 406131 66687 406134
rect 123201 406131 123267 406134
rect 582557 404970 582623 404973
rect 583520 404970 584960 405060
rect 582557 404968 584960 404970
rect 582557 404912 582562 404968
rect 582618 404912 584960 404968
rect 582557 404910 584960 404912
rect 582557 404907 582623 404910
rect 583520 404820 584960 404910
rect 120625 404290 120691 404293
rect 120582 404288 120691 404290
rect 120582 404232 120630 404288
rect 120686 404232 120691 404288
rect 120582 404227 120691 404232
rect 66345 403746 66411 403749
rect 66345 403744 68908 403746
rect 66345 403688 66350 403744
rect 66406 403688 68908 403744
rect 120582 403716 120642 404227
rect 66345 403686 68908 403688
rect 66345 403683 66411 403686
rect 66805 401570 66871 401573
rect 124121 401570 124187 401573
rect 66805 401568 68908 401570
rect 66805 401512 66810 401568
rect 66866 401512 68908 401568
rect 66805 401510 68908 401512
rect 120612 401568 124187 401570
rect 120612 401512 124126 401568
rect 124182 401512 124187 401568
rect 120612 401510 124187 401512
rect 66805 401507 66871 401510
rect 124121 401507 124187 401510
rect 66345 399394 66411 399397
rect 123477 399394 123543 399397
rect 66345 399392 68908 399394
rect 66345 399336 66350 399392
rect 66406 399336 68908 399392
rect 66345 399334 68908 399336
rect 120612 399392 123543 399394
rect 120612 399336 123482 399392
rect 123538 399336 123543 399392
rect 120612 399334 123543 399336
rect 66345 399331 66411 399334
rect 123477 399331 123543 399334
rect -960 397490 480 397580
rect 2773 397490 2839 397493
rect -960 397488 2839 397490
rect -960 397432 2778 397488
rect 2834 397432 2839 397488
rect -960 397430 2839 397432
rect -960 397340 480 397430
rect 2773 397427 2839 397430
rect 66989 396946 67055 396949
rect 67357 396946 67423 396949
rect 121453 396946 121519 396949
rect 66989 396944 68908 396946
rect 66989 396888 66994 396944
rect 67050 396888 67362 396944
rect 67418 396888 68908 396944
rect 66989 396886 68908 396888
rect 120612 396944 121519 396946
rect 120612 396888 121458 396944
rect 121514 396888 121519 396944
rect 120612 396886 121519 396888
rect 66989 396883 67055 396886
rect 67357 396883 67423 396886
rect 121453 396883 121519 396886
rect 67541 394770 67607 394773
rect 122966 394770 122972 394772
rect 67541 394768 68908 394770
rect 67541 394712 67546 394768
rect 67602 394712 68908 394768
rect 67541 394710 68908 394712
rect 120612 394710 122972 394770
rect 67541 394707 67607 394710
rect 122966 394708 122972 394710
rect 123036 394770 123042 394772
rect 123661 394770 123727 394773
rect 123036 394768 123727 394770
rect 123036 394712 123666 394768
rect 123722 394712 123727 394768
rect 123036 394710 123727 394712
rect 123036 394708 123042 394710
rect 123661 394707 123727 394710
rect 122649 393274 122715 393277
rect 122782 393274 122788 393276
rect 122649 393272 122788 393274
rect 122649 393216 122654 393272
rect 122710 393216 122788 393272
rect 122649 393214 122788 393216
rect 122649 393211 122715 393214
rect 122782 393212 122788 393214
rect 122852 393212 122858 393276
rect 66110 392532 66116 392596
rect 66180 392594 66186 392596
rect 66253 392594 66319 392597
rect 122741 392594 122807 392597
rect 122925 392594 122991 392597
rect 66180 392592 68908 392594
rect 66180 392536 66258 392592
rect 66314 392536 68908 392592
rect 66180 392534 68908 392536
rect 120612 392592 122991 392594
rect 120612 392536 122746 392592
rect 122802 392536 122930 392592
rect 122986 392536 122991 392592
rect 120612 392534 122991 392536
rect 66180 392532 66186 392534
rect 66253 392531 66319 392534
rect 122741 392531 122807 392534
rect 122925 392531 122991 392534
rect 583520 391628 584960 391868
rect 68645 391234 68711 391237
rect 72366 391234 72372 391236
rect 68645 391232 72372 391234
rect 68645 391176 68650 391232
rect 68706 391176 72372 391232
rect 68645 391174 72372 391176
rect 68645 391171 68711 391174
rect 72366 391172 72372 391174
rect 72436 391172 72442 391236
rect 65885 390962 65951 390965
rect 86309 390962 86375 390965
rect 92841 390964 92907 390965
rect 65885 390960 86375 390962
rect 65885 390904 65890 390960
rect 65946 390904 86314 390960
rect 86370 390904 86375 390960
rect 65885 390902 86375 390904
rect 65885 390899 65951 390902
rect 86309 390899 86375 390902
rect 92790 390900 92796 390964
rect 92860 390962 92907 390964
rect 102133 390964 102199 390965
rect 102133 390962 102180 390964
rect 92860 390960 92952 390962
rect 92902 390904 92952 390960
rect 92860 390902 92952 390904
rect 102088 390960 102180 390962
rect 102088 390904 102138 390960
rect 102088 390902 102180 390904
rect 92860 390900 92907 390902
rect 92841 390899 92907 390900
rect 102133 390900 102180 390902
rect 102244 390900 102250 390964
rect 111006 390900 111012 390964
rect 111076 390962 111082 390964
rect 118693 390962 118759 390965
rect 111076 390960 118759 390962
rect 111076 390904 118698 390960
rect 118754 390904 118759 390960
rect 111076 390902 118759 390904
rect 111076 390900 111082 390902
rect 102133 390899 102199 390900
rect 118693 390899 118759 390902
rect 115749 390690 115815 390693
rect 120717 390690 120783 390693
rect 115749 390688 120783 390690
rect 115749 390632 115754 390688
rect 115810 390632 120722 390688
rect 120778 390632 120783 390688
rect 115749 390630 120783 390632
rect 115749 390627 115815 390630
rect 120717 390627 120783 390630
rect 69606 390356 69612 390420
rect 69676 390418 69682 390420
rect 69933 390418 69999 390421
rect 71865 390420 71931 390421
rect 71814 390418 71820 390420
rect 69676 390416 69999 390418
rect 69676 390360 69938 390416
rect 69994 390360 69999 390416
rect 69676 390358 69999 390360
rect 71774 390358 71820 390418
rect 71884 390416 71931 390420
rect 71926 390360 71931 390416
rect 69676 390356 69682 390358
rect 69933 390355 69999 390358
rect 71814 390356 71820 390358
rect 71884 390356 71931 390360
rect 71865 390355 71931 390356
rect 80053 390418 80119 390421
rect 80605 390418 80671 390421
rect 80053 390416 80671 390418
rect 80053 390360 80058 390416
rect 80114 390360 80610 390416
rect 80666 390360 80671 390416
rect 80053 390358 80671 390360
rect 80053 390355 80119 390358
rect 80605 390355 80671 390358
rect 89662 390356 89668 390420
rect 89732 390418 89738 390420
rect 89805 390418 89871 390421
rect 89732 390416 89871 390418
rect 89732 390360 89810 390416
rect 89866 390360 89871 390416
rect 89732 390358 89871 390360
rect 89732 390356 89738 390358
rect 89805 390355 89871 390358
rect 91134 390356 91140 390420
rect 91204 390418 91210 390420
rect 91277 390418 91343 390421
rect 91204 390416 91343 390418
rect 91204 390360 91282 390416
rect 91338 390360 91343 390416
rect 91204 390358 91343 390360
rect 91204 390356 91210 390358
rect 91277 390355 91343 390358
rect 96654 390356 96660 390420
rect 96724 390418 96730 390420
rect 97349 390418 97415 390421
rect 96724 390416 97415 390418
rect 96724 390360 97354 390416
rect 97410 390360 97415 390416
rect 96724 390358 97415 390360
rect 96724 390356 96730 390358
rect 97349 390355 97415 390358
rect 98126 390356 98132 390420
rect 98196 390418 98202 390420
rect 98821 390418 98887 390421
rect 98196 390416 98887 390418
rect 98196 390360 98826 390416
rect 98882 390360 98887 390416
rect 98196 390358 98887 390360
rect 98196 390356 98202 390358
rect 98821 390355 98887 390358
rect 100661 390420 100727 390421
rect 100661 390416 100708 390420
rect 100772 390418 100778 390420
rect 100661 390360 100666 390416
rect 100661 390356 100708 390360
rect 100772 390358 100818 390418
rect 100772 390356 100778 390358
rect 104934 390356 104940 390420
rect 105004 390418 105010 390420
rect 105077 390418 105143 390421
rect 105004 390416 105143 390418
rect 105004 390360 105082 390416
rect 105138 390360 105143 390416
rect 105004 390358 105143 390360
rect 105004 390356 105010 390358
rect 100661 390355 100727 390356
rect 105077 390355 105143 390358
rect 106406 390356 106412 390420
rect 106476 390418 106482 390420
rect 106549 390418 106615 390421
rect 106476 390416 106615 390418
rect 106476 390360 106554 390416
rect 106610 390360 106615 390416
rect 106476 390358 106615 390360
rect 106476 390356 106482 390358
rect 106549 390355 106615 390358
rect 107694 390356 107700 390420
rect 107764 390418 107770 390420
rect 108021 390418 108087 390421
rect 107764 390416 108087 390418
rect 107764 390360 108026 390416
rect 108082 390360 108087 390416
rect 107764 390358 108087 390360
rect 107764 390356 107770 390358
rect 108021 390355 108087 390358
rect 109166 390356 109172 390420
rect 109236 390418 109242 390420
rect 109493 390418 109559 390421
rect 109236 390416 109559 390418
rect 109236 390360 109498 390416
rect 109554 390360 109559 390416
rect 109236 390358 109559 390360
rect 109236 390356 109242 390358
rect 109493 390355 109559 390358
rect 115933 390420 115999 390421
rect 115933 390416 115980 390420
rect 116044 390418 116050 390420
rect 115933 390360 115938 390416
rect 115933 390356 115980 390360
rect 116044 390358 116090 390418
rect 116044 390356 116050 390358
rect 120022 390356 120028 390420
rect 120092 390418 120098 390420
rect 120165 390418 120231 390421
rect 120092 390416 120231 390418
rect 120092 390360 120170 390416
rect 120226 390360 120231 390416
rect 120092 390358 120231 390360
rect 120092 390356 120098 390358
rect 115933 390355 115999 390356
rect 120165 390355 120231 390358
rect 66161 389194 66227 389197
rect 80053 389194 80119 389197
rect 66161 389192 80119 389194
rect 66161 389136 66166 389192
rect 66222 389136 80058 389192
rect 80114 389136 80119 389192
rect 66161 389134 80119 389136
rect 66161 389131 66227 389134
rect 80053 389131 80119 389134
rect 67766 388996 67772 389060
rect 67836 389058 67842 389060
rect 68134 389058 68140 389060
rect 67836 388998 68140 389058
rect 67836 388996 67842 388998
rect 68134 388996 68140 388998
rect 68204 389058 68210 389060
rect 68461 389058 68527 389061
rect 68204 389056 68527 389058
rect 68204 389000 68466 389056
rect 68522 389000 68527 389056
rect 68204 388998 68527 389000
rect 68204 388996 68210 388998
rect 68461 388995 68527 388998
rect 72049 389058 72115 389061
rect 73061 389058 73127 389061
rect 72049 389056 73127 389058
rect 72049 389000 72054 389056
rect 72110 389000 73066 389056
rect 73122 389000 73127 389056
rect 72049 388998 73127 389000
rect 72049 388995 72115 388998
rect 73061 388995 73127 388998
rect 89713 389058 89779 389061
rect 95182 389058 95188 389060
rect 89713 389056 95188 389058
rect 89713 389000 89718 389056
rect 89774 389000 95188 389056
rect 89713 388998 95188 389000
rect 89713 388995 89779 388998
rect 95182 388996 95188 388998
rect 95252 389058 95258 389060
rect 95877 389058 95943 389061
rect 95252 389056 95943 389058
rect 95252 389000 95882 389056
rect 95938 389000 95943 389056
rect 95252 388998 95943 389000
rect 95252 388996 95258 388998
rect 95877 388995 95943 388998
rect 101121 389058 101187 389061
rect 101949 389058 102015 389061
rect 111793 389060 111859 389061
rect 111742 389058 111748 389060
rect 101121 389056 102015 389058
rect 101121 389000 101126 389056
rect 101182 389000 101954 389056
rect 102010 389000 102015 389056
rect 101121 388998 102015 389000
rect 111666 388998 111748 389058
rect 111812 389058 111859 389060
rect 112621 389058 112687 389061
rect 111812 389056 112687 389058
rect 111854 389000 112626 389056
rect 112682 389000 112687 389056
rect 101121 388995 101187 388998
rect 101949 388995 102015 388998
rect 111742 388996 111748 388998
rect 111812 388998 112687 389000
rect 111812 388996 111859 388998
rect 111793 388995 111859 388996
rect 112621 388995 112687 388998
rect 59077 388922 59143 388925
rect 88885 388922 88951 388925
rect 59077 388920 88951 388922
rect 59077 388864 59082 388920
rect 59138 388864 88890 388920
rect 88946 388864 88951 388920
rect 59077 388862 88951 388864
rect 59077 388859 59143 388862
rect 88885 388859 88951 388862
rect 99966 388860 99972 388924
rect 100036 388922 100042 388924
rect 100036 388862 103530 388922
rect 100036 388860 100042 388862
rect 3417 388786 3483 388789
rect 90357 388786 90423 388789
rect 3417 388784 90423 388786
rect 3417 388728 3422 388784
rect 3478 388728 90362 388784
rect 90418 388728 90423 388784
rect 3417 388726 90423 388728
rect 3417 388723 3483 388726
rect 90357 388723 90423 388726
rect 103470 388650 103530 388862
rect 113173 388650 113239 388653
rect 114093 388650 114159 388653
rect 103470 388648 114159 388650
rect 103470 388592 113178 388648
rect 113234 388592 114098 388648
rect 114154 388592 114159 388648
rect 103470 388590 114159 388592
rect 113173 388587 113239 388590
rect 114093 388587 114159 388590
rect 64597 387698 64663 387701
rect 79317 387698 79383 387701
rect 64597 387696 79383 387698
rect 64597 387640 64602 387696
rect 64658 387640 79322 387696
rect 79378 387640 79383 387696
rect 64597 387638 79383 387640
rect 64597 387635 64663 387638
rect 79317 387635 79383 387638
rect 52361 385658 52427 385661
rect 122649 385658 122715 385661
rect 52361 385656 122715 385658
rect 52361 385600 52366 385656
rect 52422 385600 122654 385656
rect 122710 385600 122715 385656
rect 52361 385598 122715 385600
rect 52361 385595 52427 385598
rect 122649 385595 122715 385598
rect -960 384284 480 384524
rect 67633 380218 67699 380221
rect 123017 380218 123083 380221
rect 67633 380216 123083 380218
rect 67633 380160 67638 380216
rect 67694 380160 123022 380216
rect 123078 380160 123083 380216
rect 67633 380158 123083 380160
rect 67633 380155 67699 380158
rect 123017 380155 123083 380158
rect 582741 378450 582807 378453
rect 583520 378450 584960 378540
rect 582741 378448 584960 378450
rect 582741 378392 582746 378448
rect 582802 378392 584960 378448
rect 582741 378390 584960 378392
rect 582741 378387 582807 378390
rect 583520 378300 584960 378390
rect 133137 377362 133203 377365
rect 166942 377362 166948 377364
rect 133137 377360 166948 377362
rect 133137 377304 133142 377360
rect 133198 377304 166948 377360
rect 133137 377302 166948 377304
rect 133137 377299 133203 377302
rect 166942 377300 166948 377302
rect 167012 377300 167018 377364
rect 68870 375940 68876 376004
rect 68940 376002 68946 376004
rect 145557 376002 145623 376005
rect 68940 376000 145623 376002
rect 68940 375944 145562 376000
rect 145618 375944 145623 376000
rect 68940 375942 145623 375944
rect 68940 375940 68946 375942
rect 145557 375939 145623 375942
rect 120809 375458 120875 375461
rect 244222 375458 244228 375460
rect 120809 375456 244228 375458
rect 120809 375400 120814 375456
rect 120870 375400 244228 375456
rect 120809 375398 244228 375400
rect 120809 375395 120875 375398
rect 244222 375396 244228 375398
rect 244292 375396 244298 375460
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 102041 371378 102107 371381
rect 321553 371378 321619 371381
rect 102041 371376 321619 371378
rect 102041 371320 102046 371376
rect 102102 371320 321558 371376
rect 321614 371320 321619 371376
rect 102041 371318 321619 371320
rect 102041 371315 102107 371318
rect 321553 371315 321619 371318
rect 108849 370698 108915 370701
rect 161473 370698 161539 370701
rect 108849 370696 161539 370698
rect 108849 370640 108854 370696
rect 108910 370640 161478 370696
rect 161534 370640 161539 370696
rect 108849 370638 161539 370640
rect 108849 370635 108915 370638
rect 161473 370635 161539 370638
rect 70158 370500 70164 370564
rect 70228 370562 70234 370564
rect 122833 370562 122899 370565
rect 70228 370560 122899 370562
rect 70228 370504 122838 370560
rect 122894 370504 122899 370560
rect 70228 370502 122899 370504
rect 70228 370500 70234 370502
rect 122833 370499 122899 370502
rect 96429 369612 96495 369613
rect 96429 369608 96476 369612
rect 96540 369610 96546 369612
rect 96429 369552 96434 369608
rect 96429 369548 96476 369552
rect 96540 369550 96586 369610
rect 96540 369548 96546 369550
rect 96429 369547 96495 369548
rect 96429 368522 96495 368525
rect 248413 368522 248479 368525
rect 96429 368520 248479 368522
rect 96429 368464 96434 368520
rect 96490 368464 248418 368520
rect 248474 368464 248479 368520
rect 96429 368462 248479 368464
rect 96429 368459 96495 368462
rect 248413 368459 248479 368462
rect 114318 368324 114324 368388
rect 114388 368386 114394 368388
rect 119337 368386 119403 368389
rect 114388 368384 119403 368386
rect 114388 368328 119342 368384
rect 119398 368328 119403 368384
rect 114388 368326 119403 368328
rect 114388 368324 114394 368326
rect 119337 368323 119403 368326
rect 69790 367644 69796 367708
rect 69860 367706 69866 367708
rect 122925 367706 122991 367709
rect 69860 367704 122991 367706
rect 69860 367648 122930 367704
rect 122986 367648 122991 367704
rect 69860 367646 122991 367648
rect 69860 367644 69866 367646
rect 122925 367643 122991 367646
rect 127617 367162 127683 367165
rect 208894 367162 208900 367164
rect 127617 367160 208900 367162
rect 127617 367104 127622 367160
rect 127678 367104 208900 367160
rect 127617 367102 208900 367104
rect 127617 367099 127683 367102
rect 208894 367100 208900 367102
rect 208964 367100 208970 367164
rect 135897 367026 135963 367029
rect 136541 367026 136607 367029
rect 135897 367024 136607 367026
rect 135897 366968 135902 367024
rect 135958 366968 136546 367024
rect 136602 366968 136607 367024
rect 135897 366966 136607 366968
rect 135897 366963 135963 366966
rect 136541 366963 136607 366966
rect 57697 366346 57763 366349
rect 160093 366346 160159 366349
rect 57697 366344 160159 366346
rect 57697 366288 57702 366344
rect 57758 366288 160098 366344
rect 160154 366288 160159 366344
rect 57697 366286 160159 366288
rect 57697 366283 57763 366286
rect 160093 366283 160159 366286
rect 136541 365802 136607 365805
rect 218646 365802 218652 365804
rect 136541 365800 218652 365802
rect 136541 365744 136546 365800
rect 136602 365744 218652 365800
rect 136541 365742 218652 365744
rect 136541 365739 136607 365742
rect 218646 365740 218652 365742
rect 218716 365740 218722 365804
rect 582373 365122 582439 365125
rect 583520 365122 584960 365212
rect 582373 365120 584960 365122
rect 582373 365064 582378 365120
rect 582434 365064 584960 365120
rect 582373 365062 584960 365064
rect 582373 365059 582439 365062
rect 80053 364986 80119 364989
rect 157333 364986 157399 364989
rect 80053 364984 157399 364986
rect 80053 364928 80058 364984
rect 80114 364928 157338 364984
rect 157394 364928 157399 364984
rect 583520 364972 584960 365062
rect 80053 364926 157399 364928
rect 80053 364923 80119 364926
rect 157333 364923 157399 364926
rect 99281 364442 99347 364445
rect 184054 364442 184060 364444
rect 99281 364440 184060 364442
rect 99281 364384 99286 364440
rect 99342 364384 184060 364440
rect 99281 364382 184060 364384
rect 99281 364379 99347 364382
rect 184054 364380 184060 364382
rect 184124 364380 184130 364444
rect 93761 364306 93827 364309
rect 128997 364306 129063 364309
rect 93761 364304 129063 364306
rect 93761 364248 93766 364304
rect 93822 364248 129002 364304
rect 129058 364248 129063 364304
rect 93761 364246 129063 364248
rect 93761 364243 93827 364246
rect 128997 364243 129063 364246
rect 100017 363762 100083 363765
rect 151721 363762 151787 363765
rect 100017 363760 151787 363762
rect 100017 363704 100022 363760
rect 100078 363704 151726 363760
rect 151782 363704 151787 363760
rect 100017 363702 151787 363704
rect 100017 363699 100083 363702
rect 151721 363699 151787 363702
rect 128997 363626 129063 363629
rect 212901 363626 212967 363629
rect 128997 363624 212967 363626
rect 128997 363568 129002 363624
rect 129058 363568 212906 363624
rect 212962 363568 212967 363624
rect 128997 363566 212967 363568
rect 128997 363563 129063 363566
rect 212901 363563 212967 363566
rect 93117 363082 93183 363085
rect 93761 363082 93827 363085
rect 93117 363080 93827 363082
rect 93117 363024 93122 363080
rect 93178 363024 93766 363080
rect 93822 363024 93827 363080
rect 93117 363022 93827 363024
rect 93117 363019 93183 363022
rect 93761 363019 93827 363022
rect 76557 362266 76623 362269
rect 138054 362266 138060 362268
rect 76557 362264 138060 362266
rect 76557 362208 76562 362264
rect 76618 362208 138060 362264
rect 76557 362206 138060 362208
rect 76557 362203 76623 362206
rect 138054 362204 138060 362206
rect 138124 362204 138130 362268
rect 147438 361796 147444 361860
rect 147508 361858 147514 361860
rect 218237 361858 218303 361861
rect 147508 361856 218303 361858
rect 147508 361800 218242 361856
rect 218298 361800 218303 361856
rect 147508 361798 218303 361800
rect 147508 361796 147514 361798
rect 218237 361795 218303 361798
rect 121453 361722 121519 361725
rect 122598 361722 122604 361724
rect 121453 361720 122604 361722
rect 121453 361664 121458 361720
rect 121514 361664 122604 361720
rect 121453 361662 122604 361664
rect 121453 361659 121519 361662
rect 122598 361660 122604 361662
rect 122668 361722 122674 361724
rect 222837 361722 222903 361725
rect 122668 361720 222903 361722
rect 122668 361664 222842 361720
rect 222898 361664 222903 361720
rect 122668 361662 222903 361664
rect 122668 361660 122674 361662
rect 222837 361659 222903 361662
rect 84101 360906 84167 360909
rect 101397 360906 101463 360909
rect 84101 360904 101463 360906
rect 84101 360848 84106 360904
rect 84162 360848 101402 360904
rect 101458 360848 101463 360904
rect 84101 360846 101463 360848
rect 84101 360843 84167 360846
rect 101397 360843 101463 360846
rect 151077 360906 151143 360909
rect 173157 360906 173223 360909
rect 151077 360904 173223 360906
rect 151077 360848 151082 360904
rect 151138 360848 173162 360904
rect 173218 360848 173223 360904
rect 151077 360846 173223 360848
rect 151077 360843 151143 360846
rect 173157 360843 173223 360846
rect 123293 360228 123359 360229
rect 123293 360224 123340 360228
rect 123404 360226 123410 360228
rect 248454 360226 248460 360228
rect 123293 360168 123298 360224
rect 123293 360164 123340 360168
rect 123404 360166 248460 360226
rect 123404 360164 123410 360166
rect 248454 360164 248460 360166
rect 248524 360164 248530 360228
rect 123293 360163 123359 360164
rect 76557 359274 76623 359277
rect 77201 359274 77267 359277
rect 76557 359272 77267 359274
rect 76557 359216 76562 359272
rect 76618 359216 77206 359272
rect 77262 359216 77267 359272
rect 76557 359214 77267 359216
rect 76557 359211 76623 359214
rect 77201 359211 77267 359214
rect 101397 359002 101463 359005
rect 101949 359002 102015 359005
rect 202137 359002 202203 359005
rect 101397 359000 202203 359002
rect 101397 358944 101402 359000
rect 101458 358944 101954 359000
rect 102010 358944 202142 359000
rect 202198 358944 202203 359000
rect 101397 358942 202203 358944
rect 101397 358939 101463 358942
rect 101949 358939 102015 358942
rect 202137 358939 202203 358942
rect 77201 358866 77267 358869
rect 252502 358866 252508 358868
rect 77201 358864 252508 358866
rect 77201 358808 77206 358864
rect 77262 358808 252508 358864
rect 77201 358806 252508 358808
rect 77201 358803 77267 358806
rect 252502 358804 252508 358806
rect 252572 358804 252578 358868
rect 109534 358668 109540 358732
rect 109604 358730 109610 358732
rect 109677 358730 109743 358733
rect 109604 358728 109743 358730
rect 109604 358672 109682 358728
rect 109738 358672 109743 358728
rect 109604 358670 109743 358672
rect 109604 358668 109610 358670
rect 109677 358667 109743 358670
rect -960 358458 480 358548
rect 3509 358458 3575 358461
rect -960 358456 3575 358458
rect -960 358400 3514 358456
rect 3570 358400 3575 358456
rect -960 358398 3575 358400
rect -960 358308 480 358398
rect 3509 358395 3575 358398
rect 130377 358186 130443 358189
rect 158069 358186 158135 358189
rect 130377 358184 158135 358186
rect 130377 358128 130382 358184
rect 130438 358128 158074 358184
rect 158130 358128 158135 358184
rect 130377 358126 158135 358128
rect 130377 358123 130443 358126
rect 158069 358123 158135 358126
rect 96521 358050 96587 358053
rect 125685 358050 125751 358053
rect 262213 358050 262279 358053
rect 96521 358048 262279 358050
rect 96521 357992 96526 358048
rect 96582 357992 125690 358048
rect 125746 357992 262218 358048
rect 262274 357992 262279 358048
rect 96521 357990 262279 357992
rect 96521 357987 96587 357990
rect 125685 357987 125751 357990
rect 262213 357987 262279 357990
rect 109677 357506 109743 357509
rect 193857 357506 193923 357509
rect 109677 357504 193923 357506
rect 109677 357448 109682 357504
rect 109738 357448 193862 357504
rect 193918 357448 193923 357504
rect 109677 357446 193923 357448
rect 109677 357443 109743 357446
rect 193857 357443 193923 357446
rect 151169 357370 151235 357373
rect 151721 357370 151787 357373
rect 160737 357370 160803 357373
rect 151169 357368 160803 357370
rect 151169 357312 151174 357368
rect 151230 357312 151726 357368
rect 151782 357312 160742 357368
rect 160798 357312 160803 357368
rect 151169 357310 160803 357312
rect 151169 357307 151235 357310
rect 151721 357307 151787 357310
rect 160737 357307 160803 357310
rect 92381 356690 92447 356693
rect 121453 356690 121519 356693
rect 92381 356688 121519 356690
rect 92381 356632 92386 356688
rect 92442 356632 121458 356688
rect 121514 356632 121519 356688
rect 92381 356630 121519 356632
rect 92381 356627 92447 356630
rect 121453 356627 121519 356630
rect 129089 356690 129155 356693
rect 151854 356690 151860 356692
rect 129089 356688 151860 356690
rect 129089 356632 129094 356688
rect 129150 356632 151860 356688
rect 129089 356630 151860 356632
rect 129089 356627 129155 356630
rect 151854 356628 151860 356630
rect 151924 356628 151930 356692
rect 111333 356146 111399 356149
rect 111558 356146 111564 356148
rect 111333 356144 111564 356146
rect 111333 356088 111338 356144
rect 111394 356088 111564 356144
rect 111333 356086 111564 356088
rect 111333 356083 111399 356086
rect 111558 356084 111564 356086
rect 111628 356146 111634 356148
rect 200757 356146 200823 356149
rect 111628 356144 200823 356146
rect 111628 356088 200762 356144
rect 200818 356088 200823 356144
rect 111628 356086 200823 356088
rect 111628 356084 111634 356086
rect 200757 356083 200823 356086
rect 110413 355874 110479 355877
rect 111701 355874 111767 355877
rect 110413 355872 111767 355874
rect 110413 355816 110418 355872
rect 110474 355816 111706 355872
rect 111762 355816 111767 355872
rect 110413 355814 111767 355816
rect 110413 355811 110479 355814
rect 111701 355811 111767 355814
rect 71037 355330 71103 355333
rect 123293 355330 123359 355333
rect 71037 355328 123359 355330
rect 71037 355272 71042 355328
rect 71098 355272 123298 355328
rect 123354 355272 123359 355328
rect 71037 355270 123359 355272
rect 71037 355267 71103 355270
rect 123293 355267 123359 355270
rect 129641 354922 129707 354925
rect 232446 354922 232452 354924
rect 129641 354920 232452 354922
rect 129641 354864 129646 354920
rect 129702 354864 232452 354920
rect 129641 354862 232452 354864
rect 129641 354859 129707 354862
rect 232446 354860 232452 354862
rect 232516 354860 232522 354924
rect 111701 354786 111767 354789
rect 246297 354786 246363 354789
rect 111701 354784 246363 354786
rect 111701 354728 111706 354784
rect 111762 354728 246302 354784
rect 246358 354728 246363 354784
rect 111701 354726 246363 354728
rect 111701 354723 111767 354726
rect 246297 354723 246363 354726
rect 60549 353970 60615 353973
rect 156689 353970 156755 353973
rect 60549 353968 156755 353970
rect 60549 353912 60554 353968
rect 60610 353912 156694 353968
rect 156750 353912 156755 353968
rect 60549 353910 156755 353912
rect 60549 353907 60615 353910
rect 156689 353907 156755 353910
rect 93853 353562 93919 353565
rect 197997 353562 198063 353565
rect 93853 353560 198063 353562
rect 93853 353504 93858 353560
rect 93914 353504 198002 353560
rect 198058 353504 198063 353560
rect 93853 353502 198063 353504
rect 93853 353499 93919 353502
rect 197997 353499 198063 353502
rect 142061 353426 142127 353429
rect 331213 353426 331279 353429
rect 142061 353424 331279 353426
rect 142061 353368 142066 353424
rect 142122 353368 331218 353424
rect 331274 353368 331279 353424
rect 142061 353366 331279 353368
rect 142061 353363 142127 353366
rect 331213 353363 331279 353366
rect 92657 353292 92723 353293
rect 92606 353290 92612 353292
rect 92566 353230 92612 353290
rect 92676 353288 92723 353292
rect 92718 353232 92723 353288
rect 92606 353228 92612 353230
rect 92676 353228 92723 353232
rect 92657 353227 92723 353228
rect 114553 352066 114619 352069
rect 115841 352066 115907 352069
rect 227437 352066 227503 352069
rect 114553 352064 227503 352066
rect 114553 352008 114558 352064
rect 114614 352008 115846 352064
rect 115902 352008 227442 352064
rect 227498 352008 227503 352064
rect 114553 352006 227503 352008
rect 114553 352003 114619 352006
rect 115841 352003 115907 352006
rect 227437 352003 227503 352006
rect 59169 351930 59235 351933
rect 188521 351930 188587 351933
rect 59169 351928 188587 351930
rect 59169 351872 59174 351928
rect 59230 351872 188526 351928
rect 188582 351872 188587 351928
rect 59169 351870 188587 351872
rect 59169 351867 59235 351870
rect 188521 351867 188587 351870
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect 69606 351052 69612 351116
rect 69676 351114 69682 351116
rect 86217 351114 86283 351117
rect 69676 351112 86283 351114
rect 69676 351056 86222 351112
rect 86278 351056 86283 351112
rect 69676 351054 86283 351056
rect 69676 351052 69682 351054
rect 86217 351051 86283 351054
rect 86861 351114 86927 351117
rect 102358 351114 102364 351116
rect 86861 351112 102364 351114
rect 86861 351056 86866 351112
rect 86922 351056 102364 351112
rect 86861 351054 102364 351056
rect 86861 351051 86927 351054
rect 102358 351052 102364 351054
rect 102428 351052 102434 351116
rect 107469 351114 107535 351117
rect 155166 351114 155172 351116
rect 107469 351112 155172 351114
rect 107469 351056 107474 351112
rect 107530 351056 155172 351112
rect 107469 351054 155172 351056
rect 107469 351051 107535 351054
rect 155166 351052 155172 351054
rect 155236 351052 155242 351116
rect 99189 350706 99255 350709
rect 178534 350706 178540 350708
rect 99189 350704 178540 350706
rect 99189 350648 99194 350704
rect 99250 350648 178540 350704
rect 99189 350646 178540 350648
rect 99189 350643 99255 350646
rect 178534 350644 178540 350646
rect 178604 350644 178610 350708
rect 126973 350570 127039 350573
rect 127709 350570 127775 350573
rect 233734 350570 233740 350572
rect 126973 350568 233740 350570
rect 126973 350512 126978 350568
rect 127034 350512 127714 350568
rect 127770 350512 233740 350568
rect 126973 350510 233740 350512
rect 126973 350507 127039 350510
rect 127709 350507 127775 350510
rect 233734 350508 233740 350510
rect 233804 350508 233810 350572
rect 136541 349890 136607 349893
rect 138013 349890 138079 349893
rect 136541 349888 138079 349890
rect 136541 349832 136546 349888
rect 136602 349832 138018 349888
rect 138074 349832 138079 349888
rect 136541 349830 138079 349832
rect 136541 349827 136607 349830
rect 138013 349827 138079 349830
rect 77293 349754 77359 349757
rect 136030 349754 136036 349756
rect 77293 349752 136036 349754
rect 77293 349696 77298 349752
rect 77354 349696 136036 349752
rect 77293 349694 136036 349696
rect 77293 349691 77359 349694
rect 136030 349692 136036 349694
rect 136100 349692 136106 349756
rect 144913 349754 144979 349757
rect 145557 349754 145623 349757
rect 144913 349752 151830 349754
rect 144913 349696 144918 349752
rect 144974 349696 145562 349752
rect 145618 349696 151830 349752
rect 144913 349694 151830 349696
rect 144913 349691 144979 349694
rect 145557 349691 145623 349694
rect 151770 349482 151830 349694
rect 206277 349482 206343 349485
rect 151770 349480 206343 349482
rect 151770 349424 206282 349480
rect 206338 349424 206343 349480
rect 151770 349422 206343 349424
rect 206277 349419 206343 349422
rect 108941 349346 109007 349349
rect 184197 349346 184263 349349
rect 108941 349344 184263 349346
rect 108941 349288 108946 349344
rect 109002 349288 184202 349344
rect 184258 349288 184263 349344
rect 108941 349286 184263 349288
rect 108941 349283 109007 349286
rect 184197 349283 184263 349286
rect 117313 349210 117379 349213
rect 118550 349210 118556 349212
rect 117313 349208 118556 349210
rect 117313 349152 117318 349208
rect 117374 349152 118556 349208
rect 117313 349150 118556 349152
rect 117313 349147 117379 349150
rect 118550 349148 118556 349150
rect 118620 349210 118626 349212
rect 263685 349210 263751 349213
rect 118620 349208 263751 349210
rect 118620 349152 263690 349208
rect 263746 349152 263751 349208
rect 118620 349150 263751 349152
rect 118620 349148 118626 349150
rect 263685 349147 263751 349150
rect 191097 349074 191163 349077
rect 191741 349074 191807 349077
rect 580165 349074 580231 349077
rect 191097 349072 580231 349074
rect 191097 349016 191102 349072
rect 191158 349016 191746 349072
rect 191802 349016 580170 349072
rect 580226 349016 580231 349072
rect 191097 349014 580231 349016
rect 191097 349011 191163 349014
rect 191741 349011 191807 349014
rect 580165 349011 580231 349014
rect 113081 347986 113147 347989
rect 180149 347986 180215 347989
rect 113081 347984 180215 347986
rect 113081 347928 113086 347984
rect 113142 347928 180154 347984
rect 180210 347928 180215 347984
rect 113081 347926 180215 347928
rect 113081 347923 113147 347926
rect 180149 347923 180215 347926
rect 70158 347788 70164 347852
rect 70228 347850 70234 347852
rect 223614 347850 223620 347852
rect 70228 347790 223620 347850
rect 70228 347788 70234 347790
rect 223614 347788 223620 347790
rect 223684 347788 223690 347852
rect 66662 347652 66668 347716
rect 66732 347714 66738 347716
rect 67357 347714 67423 347717
rect 66732 347712 67423 347714
rect 66732 347656 67362 347712
rect 67418 347656 67423 347712
rect 66732 347654 67423 347656
rect 66732 347652 66738 347654
rect 67357 347651 67423 347654
rect 135161 347034 135227 347037
rect 156454 347034 156460 347036
rect 135161 347032 156460 347034
rect 135161 346976 135166 347032
rect 135222 346976 156460 347032
rect 135161 346974 156460 346976
rect 135161 346971 135227 346974
rect 156454 346972 156460 346974
rect 156524 346972 156530 347036
rect 66662 346700 66668 346764
rect 66732 346762 66738 346764
rect 242249 346762 242315 346765
rect 66732 346760 242315 346762
rect 66732 346704 242254 346760
rect 242310 346704 242315 346760
rect 66732 346702 242315 346704
rect 66732 346700 66738 346702
rect 242249 346699 242315 346702
rect 115054 346564 115060 346628
rect 115124 346626 115130 346628
rect 177389 346626 177455 346629
rect 203057 346628 203123 346629
rect 203006 346626 203012 346628
rect 115124 346624 177455 346626
rect 115124 346568 177394 346624
rect 177450 346568 177455 346624
rect 115124 346566 177455 346568
rect 202966 346566 203012 346626
rect 203076 346624 203123 346628
rect 203118 346568 203123 346624
rect 115124 346564 115130 346566
rect 177389 346563 177455 346566
rect 203006 346564 203012 346566
rect 203076 346564 203123 346568
rect 203057 346563 203123 346564
rect 65977 346354 66043 346357
rect 67766 346354 67772 346356
rect 65977 346352 67772 346354
rect 65977 346296 65982 346352
rect 66038 346296 67772 346352
rect 65977 346294 67772 346296
rect 65977 346291 66043 346294
rect 67766 346292 67772 346294
rect 67836 346292 67842 346356
rect 67950 345748 67956 345812
rect 68020 345810 68026 345812
rect 115933 345810 115999 345813
rect 68020 345808 115999 345810
rect 68020 345752 115938 345808
rect 115994 345752 115999 345808
rect 68020 345750 115999 345752
rect 68020 345748 68026 345750
rect 115933 345747 115999 345750
rect 105537 345674 105603 345677
rect 153837 345674 153903 345677
rect 105537 345672 153903 345674
rect 105537 345616 105542 345672
rect 105598 345616 153842 345672
rect 153898 345616 153903 345672
rect 105537 345614 153903 345616
rect 105537 345611 105603 345614
rect 153837 345611 153903 345614
rect -960 345402 480 345492
rect 2773 345402 2839 345405
rect -960 345400 2839 345402
rect -960 345344 2778 345400
rect 2834 345344 2839 345400
rect -960 345342 2839 345344
rect -960 345252 480 345342
rect 2773 345339 2839 345342
rect 137277 345266 137343 345269
rect 186814 345266 186820 345268
rect 137277 345264 186820 345266
rect 137277 345208 137282 345264
rect 137338 345208 186820 345264
rect 137277 345206 186820 345208
rect 137277 345203 137343 345206
rect 186814 345204 186820 345206
rect 186884 345204 186890 345268
rect 118601 345130 118667 345133
rect 357433 345130 357499 345133
rect 118601 345128 357499 345130
rect 118601 345072 118606 345128
rect 118662 345072 357438 345128
rect 357494 345072 357499 345128
rect 118601 345070 357499 345072
rect 118601 345067 118667 345070
rect 357433 345067 357499 345070
rect 119337 343906 119403 343909
rect 164969 343906 165035 343909
rect 119337 343904 165035 343906
rect 119337 343848 119342 343904
rect 119398 343848 164974 343904
rect 165030 343848 165035 343904
rect 119337 343846 165035 343848
rect 119337 343843 119403 343846
rect 164969 343843 165035 343846
rect 108849 343770 108915 343773
rect 582373 343770 582439 343773
rect 108849 343768 582439 343770
rect 108849 343712 108854 343768
rect 108910 343712 582378 343768
rect 582434 343712 582439 343768
rect 108849 343710 582439 343712
rect 108849 343707 108915 343710
rect 582373 343707 582439 343710
rect 135161 342546 135227 342549
rect 176009 342546 176075 342549
rect 135161 342544 176075 342546
rect 135161 342488 135166 342544
rect 135222 342488 176014 342544
rect 176070 342488 176075 342544
rect 135161 342486 176075 342488
rect 135161 342483 135227 342486
rect 176009 342483 176075 342486
rect 105537 342410 105603 342413
rect 220077 342410 220143 342413
rect 105537 342408 220143 342410
rect 105537 342352 105542 342408
rect 105598 342352 220082 342408
rect 220138 342352 220143 342408
rect 105537 342350 220143 342352
rect 105537 342347 105603 342350
rect 220077 342347 220143 342350
rect 78581 342274 78647 342277
rect 324313 342274 324379 342277
rect 78581 342272 324379 342274
rect 78581 342216 78586 342272
rect 78642 342216 324318 342272
rect 324374 342216 324379 342272
rect 78581 342214 324379 342216
rect 78581 342211 78647 342214
rect 324313 342211 324379 342214
rect 67173 341186 67239 341189
rect 178769 341186 178835 341189
rect 67173 341184 178835 341186
rect 67173 341128 67178 341184
rect 67234 341128 178774 341184
rect 178830 341128 178835 341184
rect 67173 341126 178835 341128
rect 67173 341123 67239 341126
rect 178769 341123 178835 341126
rect 80789 341050 80855 341053
rect 228214 341050 228220 341052
rect 80789 341048 228220 341050
rect 80789 340992 80794 341048
rect 80850 340992 228220 341048
rect 80789 340990 228220 340992
rect 80789 340987 80855 340990
rect 228214 340988 228220 340990
rect 228284 340988 228290 341052
rect 111701 340914 111767 340917
rect 335997 340914 336063 340917
rect 111701 340912 336063 340914
rect 111701 340856 111706 340912
rect 111762 340856 336002 340912
rect 336058 340856 336063 340912
rect 111701 340854 336063 340856
rect 111701 340851 111767 340854
rect 335997 340851 336063 340854
rect 107837 339826 107903 339829
rect 169201 339826 169267 339829
rect 107837 339824 169267 339826
rect 107837 339768 107842 339824
rect 107898 339768 169206 339824
rect 169262 339768 169267 339824
rect 107837 339766 169267 339768
rect 107837 339763 107903 339766
rect 169201 339763 169267 339766
rect 73061 339690 73127 339693
rect 209037 339690 209103 339693
rect 73061 339688 209103 339690
rect 73061 339632 73066 339688
rect 73122 339632 209042 339688
rect 209098 339632 209103 339688
rect 73061 339630 209103 339632
rect 73061 339627 73127 339630
rect 209037 339627 209103 339630
rect 97901 339554 97967 339557
rect 291142 339554 291148 339556
rect 97901 339552 291148 339554
rect 97901 339496 97906 339552
rect 97962 339496 291148 339552
rect 97901 339494 291148 339496
rect 97901 339491 97967 339494
rect 291142 339492 291148 339494
rect 291212 339492 291218 339556
rect 89437 338466 89503 338469
rect 220169 338466 220235 338469
rect 89437 338464 220235 338466
rect 89437 338408 89442 338464
rect 89498 338408 220174 338464
rect 220230 338408 220235 338464
rect 583520 338452 584960 338692
rect 89437 338406 220235 338408
rect 89437 338403 89503 338406
rect 220169 338403 220235 338406
rect 85665 338330 85731 338333
rect 251357 338330 251423 338333
rect 85665 338328 251423 338330
rect 85665 338272 85670 338328
rect 85726 338272 251362 338328
rect 251418 338272 251423 338328
rect 85665 338270 251423 338272
rect 85665 338267 85731 338270
rect 251357 338267 251423 338270
rect 125501 338194 125567 338197
rect 339493 338194 339559 338197
rect 125501 338192 339559 338194
rect 125501 338136 125506 338192
rect 125562 338136 339498 338192
rect 339554 338136 339559 338192
rect 125501 338134 339559 338136
rect 125501 338131 125567 338134
rect 339493 338131 339559 338134
rect 160737 337378 160803 337381
rect 166901 337378 166967 337381
rect 160737 337376 166967 337378
rect 160737 337320 160742 337376
rect 160798 337320 166906 337376
rect 166962 337320 166967 337376
rect 160737 337318 166967 337320
rect 160737 337315 160803 337318
rect 166901 337315 166967 337318
rect 135253 337106 135319 337109
rect 160921 337106 160987 337109
rect 135253 337104 160987 337106
rect 135253 337048 135258 337104
rect 135314 337048 160926 337104
rect 160982 337048 160987 337104
rect 135253 337046 160987 337048
rect 135253 337043 135319 337046
rect 160921 337043 160987 337046
rect 66069 336970 66135 336973
rect 159633 336970 159699 336973
rect 66069 336968 159699 336970
rect 66069 336912 66074 336968
rect 66130 336912 159638 336968
rect 159694 336912 159699 336968
rect 66069 336910 159699 336912
rect 66069 336907 66135 336910
rect 159633 336907 159699 336910
rect 91737 336834 91803 336837
rect 185761 336834 185827 336837
rect 91737 336832 185827 336834
rect 91737 336776 91742 336832
rect 91798 336776 185766 336832
rect 185822 336776 185827 336832
rect 91737 336774 185827 336776
rect 91737 336771 91803 336774
rect 185761 336771 185827 336774
rect 114737 335746 114803 335749
rect 159214 335746 159220 335748
rect 114737 335744 159220 335746
rect 114737 335688 114742 335744
rect 114798 335688 159220 335744
rect 114737 335686 159220 335688
rect 114737 335683 114803 335686
rect 159214 335684 159220 335686
rect 159284 335684 159290 335748
rect 74625 335610 74691 335613
rect 181621 335610 181687 335613
rect 74625 335608 181687 335610
rect 74625 335552 74630 335608
rect 74686 335552 181626 335608
rect 181682 335552 181687 335608
rect 74625 335550 181687 335552
rect 74625 335547 74691 335550
rect 181621 335547 181687 335550
rect 89805 335474 89871 335477
rect 304993 335474 305059 335477
rect 89805 335472 305059 335474
rect 89805 335416 89810 335472
rect 89866 335416 304998 335472
rect 305054 335416 305059 335472
rect 89805 335414 305059 335416
rect 89805 335411 89871 335414
rect 304993 335411 305059 335414
rect 112161 334386 112227 334389
rect 212574 334386 212580 334388
rect 112161 334384 212580 334386
rect 112161 334328 112166 334384
rect 112222 334328 212580 334384
rect 112161 334326 212580 334328
rect 112161 334323 112227 334326
rect 212574 334324 212580 334326
rect 212644 334324 212650 334388
rect 70025 334250 70091 334253
rect 195329 334250 195395 334253
rect 70025 334248 195395 334250
rect 70025 334192 70030 334248
rect 70086 334192 195334 334248
rect 195390 334192 195395 334248
rect 70025 334190 195395 334192
rect 70025 334187 70091 334190
rect 195329 334187 195395 334190
rect 88609 334114 88675 334117
rect 295926 334114 295932 334116
rect 88609 334112 295932 334114
rect 88609 334056 88614 334112
rect 88670 334056 295932 334112
rect 88609 334054 295932 334056
rect 88609 334051 88675 334054
rect 295926 334052 295932 334054
rect 295996 334052 296002 334116
rect 95049 333298 95115 333301
rect 115054 333298 115060 333300
rect 95049 333296 115060 333298
rect 95049 333240 95054 333296
rect 95110 333240 115060 333296
rect 95049 333238 115060 333240
rect 95049 333235 95115 333238
rect 115054 333236 115060 333238
rect 115124 333236 115130 333300
rect 64597 332890 64663 332893
rect 155401 332890 155467 332893
rect 64597 332888 155467 332890
rect 64597 332832 64602 332888
rect 64658 332832 155406 332888
rect 155462 332832 155467 332888
rect 64597 332830 155467 332832
rect 64597 332827 64663 332830
rect 155401 332827 155467 332830
rect 117129 332754 117195 332757
rect 233969 332754 234035 332757
rect 117129 332752 234035 332754
rect 117129 332696 117134 332752
rect 117190 332696 233974 332752
rect 234030 332696 234035 332752
rect 117129 332694 234035 332696
rect 117129 332691 117195 332694
rect 233969 332691 234035 332694
rect 105997 332618 106063 332621
rect 222929 332618 222995 332621
rect 105997 332616 222995 332618
rect 105997 332560 106002 332616
rect 106058 332560 222934 332616
rect 222990 332560 222995 332616
rect 105997 332558 222995 332560
rect 105997 332555 106063 332558
rect 222929 332555 222995 332558
rect 92381 332482 92447 332485
rect 93894 332482 93900 332484
rect 92381 332480 93900 332482
rect -960 332196 480 332436
rect 92381 332424 92386 332480
rect 92442 332424 93900 332480
rect 92381 332422 93900 332424
rect 92381 332419 92447 332422
rect 93894 332420 93900 332422
rect 93964 332420 93970 332484
rect 143349 331530 143415 331533
rect 163589 331530 163655 331533
rect 143349 331528 163655 331530
rect 143349 331472 143354 331528
rect 143410 331472 163594 331528
rect 163650 331472 163655 331528
rect 143349 331470 163655 331472
rect 143349 331467 143415 331470
rect 163589 331467 163655 331470
rect 102685 331394 102751 331397
rect 160737 331394 160803 331397
rect 102685 331392 160803 331394
rect 102685 331336 102690 331392
rect 102746 331336 160742 331392
rect 160798 331336 160803 331392
rect 102685 331334 160803 331336
rect 102685 331331 102751 331334
rect 160737 331331 160803 331334
rect 69289 331258 69355 331261
rect 207657 331258 207723 331261
rect 69289 331256 207723 331258
rect 69289 331200 69294 331256
rect 69350 331200 207662 331256
rect 207718 331200 207723 331256
rect 69289 331198 207723 331200
rect 69289 331195 69355 331198
rect 207657 331195 207723 331198
rect 100017 330442 100083 330445
rect 119337 330442 119403 330445
rect 100017 330440 119403 330442
rect 100017 330384 100022 330440
rect 100078 330384 119342 330440
rect 119398 330384 119403 330440
rect 100017 330382 119403 330384
rect 100017 330379 100083 330382
rect 119337 330379 119403 330382
rect 132033 330442 132099 330445
rect 143349 330442 143415 330445
rect 132033 330440 143415 330442
rect 132033 330384 132038 330440
rect 132094 330384 143354 330440
rect 143410 330384 143415 330440
rect 132033 330382 143415 330384
rect 132033 330379 132099 330382
rect 143349 330379 143415 330382
rect 84101 330306 84167 330309
rect 84694 330306 84700 330308
rect 84101 330304 84700 330306
rect 84101 330248 84106 330304
rect 84162 330248 84700 330304
rect 84101 330246 84700 330248
rect 84101 330243 84167 330246
rect 84694 330244 84700 330246
rect 84764 330244 84770 330308
rect 109953 330306 110019 330309
rect 145414 330306 145420 330308
rect 109953 330304 145420 330306
rect 109953 330248 109958 330304
rect 110014 330248 145420 330304
rect 109953 330246 145420 330248
rect 109953 330243 110019 330246
rect 145414 330244 145420 330246
rect 145484 330244 145490 330308
rect 67541 330170 67607 330173
rect 142797 330170 142863 330173
rect 67541 330168 142863 330170
rect 67541 330112 67546 330168
rect 67602 330112 142802 330168
rect 142858 330112 142863 330168
rect 67541 330110 142863 330112
rect 67541 330107 67607 330110
rect 142797 330107 142863 330110
rect 144177 330170 144243 330173
rect 241237 330170 241303 330173
rect 144177 330168 241303 330170
rect 144177 330112 144182 330168
rect 144238 330112 241242 330168
rect 241298 330112 241303 330168
rect 144177 330110 241303 330112
rect 144177 330107 144243 330110
rect 241237 330107 241303 330110
rect 142889 330034 142955 330037
rect 174537 330034 174603 330037
rect 142889 330032 174603 330034
rect 142889 329976 142894 330032
rect 142950 329976 174542 330032
rect 174598 329976 174603 330032
rect 142889 329974 174603 329976
rect 142889 329971 142955 329974
rect 174537 329971 174603 329974
rect 142797 329082 142863 329085
rect 166349 329082 166415 329085
rect 142797 329080 166415 329082
rect 142797 329024 142802 329080
rect 142858 329024 166354 329080
rect 166410 329024 166415 329080
rect 142797 329022 166415 329024
rect 142797 329019 142863 329022
rect 166349 329019 166415 329022
rect 141969 328810 142035 328813
rect 153377 328810 153443 328813
rect 141969 328808 153443 328810
rect 141969 328752 141974 328808
rect 142030 328752 153382 328808
rect 153438 328752 153443 328808
rect 141969 328750 153443 328752
rect 141969 328747 142035 328750
rect 153377 328747 153443 328750
rect 32397 328674 32463 328677
rect 122925 328674 122991 328677
rect 32397 328672 122991 328674
rect 32397 328616 32402 328672
rect 32458 328616 122930 328672
rect 122986 328616 122991 328672
rect 32397 328614 122991 328616
rect 32397 328611 32463 328614
rect 122925 328611 122991 328614
rect 135069 328674 135135 328677
rect 137134 328674 137140 328676
rect 135069 328672 137140 328674
rect 135069 328616 135074 328672
rect 135130 328616 137140 328672
rect 135069 328614 137140 328616
rect 135069 328611 135135 328614
rect 137134 328612 137140 328614
rect 137204 328612 137210 328676
rect 7557 328538 7623 328541
rect 124949 328538 125015 328541
rect 7557 328536 125015 328538
rect 7557 328480 7562 328536
rect 7618 328480 124954 328536
rect 125010 328480 125015 328536
rect 7557 328478 125015 328480
rect 7557 328475 7623 328478
rect 124949 328475 125015 328478
rect 133873 328538 133939 328541
rect 244089 328538 244155 328541
rect 133873 328536 244155 328538
rect 133873 328480 133878 328536
rect 133934 328480 244094 328536
rect 244150 328480 244155 328536
rect 133873 328478 244155 328480
rect 133873 328475 133939 328478
rect 244089 328475 244155 328478
rect 67173 328402 67239 328405
rect 67398 328402 67404 328404
rect 67173 328400 67404 328402
rect 67173 328344 67178 328400
rect 67234 328344 67404 328400
rect 67173 328342 67404 328344
rect 67173 328339 67239 328342
rect 67398 328340 67404 328342
rect 67468 328340 67474 328404
rect 91231 327722 91297 327725
rect 92381 327722 92447 327725
rect 146201 327722 146267 327725
rect 154246 327722 154252 327724
rect 91231 327720 93870 327722
rect 91231 327664 91236 327720
rect 91292 327664 92386 327720
rect 92442 327664 93870 327720
rect 91231 327662 93870 327664
rect 91231 327659 91297 327662
rect 92381 327659 92447 327662
rect 83641 327586 83707 327589
rect 84694 327586 84700 327588
rect 83641 327584 84700 327586
rect 83641 327528 83646 327584
rect 83702 327528 84700 327584
rect 83641 327526 84700 327528
rect 83641 327523 83707 327526
rect 84694 327524 84700 327526
rect 84764 327524 84770 327588
rect 86493 327586 86559 327589
rect 86718 327586 86724 327588
rect 86493 327584 86724 327586
rect 86493 327528 86498 327584
rect 86554 327528 86724 327584
rect 86493 327526 86724 327528
rect 86493 327523 86559 327526
rect 86718 327524 86724 327526
rect 86788 327524 86794 327588
rect 93810 327586 93870 327662
rect 146201 327720 154252 327722
rect 146201 327664 146206 327720
rect 146262 327664 154252 327720
rect 146201 327662 154252 327664
rect 146201 327659 146267 327662
rect 154246 327660 154252 327662
rect 154316 327660 154322 327724
rect 155217 327722 155283 327725
rect 207974 327722 207980 327724
rect 155217 327720 207980 327722
rect 155217 327664 155222 327720
rect 155278 327664 207980 327720
rect 155217 327662 207980 327664
rect 155217 327659 155283 327662
rect 207974 327660 207980 327662
rect 208044 327660 208050 327724
rect 180241 327586 180307 327589
rect 93810 327584 180307 327586
rect 93810 327528 180246 327584
rect 180302 327528 180307 327584
rect 93810 327526 180307 327528
rect 180241 327523 180307 327526
rect 33777 327450 33843 327453
rect 114461 327450 114527 327453
rect 33777 327448 114527 327450
rect 33777 327392 33782 327448
rect 33838 327392 114466 327448
rect 114522 327392 114527 327448
rect 33777 327390 114527 327392
rect 33777 327387 33843 327390
rect 114461 327387 114527 327390
rect 123569 327450 123635 327453
rect 149881 327450 149947 327453
rect 154982 327450 154988 327452
rect 123569 327448 128370 327450
rect 123569 327392 123574 327448
rect 123630 327392 128370 327448
rect 123569 327390 128370 327392
rect 123569 327387 123635 327390
rect 40677 327314 40743 327317
rect 122833 327314 122899 327317
rect 123661 327314 123727 327317
rect 40677 327312 123727 327314
rect 40677 327256 40682 327312
rect 40738 327256 122838 327312
rect 122894 327256 123666 327312
rect 123722 327256 123727 327312
rect 40677 327254 123727 327256
rect 128310 327314 128370 327390
rect 149881 327448 154988 327450
rect 149881 327392 149886 327448
rect 149942 327392 154988 327448
rect 149881 327390 154988 327392
rect 149881 327387 149947 327390
rect 154982 327388 154988 327390
rect 155052 327388 155058 327452
rect 169109 327314 169175 327317
rect 128310 327312 169175 327314
rect 128310 327256 169114 327312
rect 169170 327256 169175 327312
rect 128310 327254 169175 327256
rect 40677 327251 40743 327254
rect 122833 327251 122899 327254
rect 123661 327251 123727 327254
rect 169109 327251 169175 327254
rect 83917 327180 83983 327181
rect 83917 327176 83964 327180
rect 84028 327178 84034 327180
rect 83917 327120 83922 327176
rect 83917 327116 83964 327120
rect 84028 327118 84074 327178
rect 84028 327116 84034 327118
rect 150382 327116 150388 327180
rect 150452 327178 150458 327180
rect 150709 327178 150775 327181
rect 150452 327176 150775 327178
rect 150452 327120 150714 327176
rect 150770 327120 150775 327176
rect 150452 327118 150775 327120
rect 150452 327116 150458 327118
rect 83917 327115 83983 327116
rect 150709 327115 150775 327118
rect 152825 327178 152891 327181
rect 154430 327178 154436 327180
rect 152825 327176 154436 327178
rect 152825 327120 152830 327176
rect 152886 327120 154436 327176
rect 152825 327118 154436 327120
rect 152825 327115 152891 327118
rect 154430 327116 154436 327118
rect 154500 327116 154506 327180
rect 69289 327042 69355 327045
rect 69933 327042 69999 327045
rect 68510 327040 69355 327042
rect 68510 326984 69294 327040
rect 69350 326984 69355 327040
rect 68510 326982 69355 326984
rect 68510 326634 68570 326982
rect 69289 326979 69355 326982
rect 69430 327040 69999 327042
rect 69430 326984 69938 327040
rect 69994 326984 69999 327040
rect 69430 326982 69999 326984
rect 69430 326740 69490 326982
rect 69933 326979 69999 326982
rect 153377 327042 153443 327045
rect 193949 327042 194015 327045
rect 153377 327040 194015 327042
rect 153377 326984 153382 327040
rect 153438 326984 193954 327040
rect 194010 326984 194015 327040
rect 153377 326982 194015 326984
rect 153377 326979 153443 326982
rect 193949 326979 194015 326982
rect 154849 326906 154915 326909
rect 156965 326906 157031 326909
rect 154849 326904 157031 326906
rect 154849 326848 154854 326904
rect 154910 326848 156970 326904
rect 157026 326848 157031 326904
rect 154849 326846 157031 326848
rect 154849 326843 154915 326846
rect 156965 326843 157031 326846
rect 68510 326574 68938 326634
rect 68878 325924 68938 326574
rect 156045 326498 156111 326501
rect 154652 326496 156111 326498
rect 154652 326440 156050 326496
rect 156106 326440 156111 326496
rect 154652 326438 156111 326440
rect 156045 326435 156111 326438
rect 192845 326362 192911 326365
rect 230473 326362 230539 326365
rect 192845 326360 230539 326362
rect 192845 326304 192850 326360
rect 192906 326304 230478 326360
rect 230534 326304 230539 326360
rect 192845 326302 230539 326304
rect 192845 326299 192911 326302
rect 230473 326299 230539 326302
rect 156137 325410 156203 325413
rect 154652 325408 156203 325410
rect 154652 325352 156142 325408
rect 156198 325352 156203 325408
rect 154652 325350 156203 325352
rect 156137 325347 156203 325350
rect 582833 325274 582899 325277
rect 583520 325274 584960 325364
rect 582833 325272 584960 325274
rect 582833 325216 582838 325272
rect 582894 325216 584960 325272
rect 582833 325214 584960 325216
rect 582833 325211 582899 325214
rect 583520 325124 584960 325214
rect 66805 324866 66871 324869
rect 66805 324864 68908 324866
rect 66805 324808 66810 324864
rect 66866 324808 68908 324864
rect 66805 324806 68908 324808
rect 66805 324803 66871 324806
rect 155166 324396 155172 324460
rect 155236 324458 155242 324460
rect 181437 324458 181503 324461
rect 155236 324456 181503 324458
rect 155236 324400 181442 324456
rect 181498 324400 181503 324456
rect 155236 324398 181503 324400
rect 155236 324396 155242 324398
rect 181437 324395 181503 324398
rect 156045 324322 156111 324325
rect 154652 324320 156111 324322
rect 154652 324264 156050 324320
rect 156106 324264 156111 324320
rect 154652 324262 156111 324264
rect 156045 324259 156111 324262
rect 66805 323778 66871 323781
rect 66805 323776 68908 323778
rect 66805 323720 66810 323776
rect 66866 323720 68908 323776
rect 66805 323718 68908 323720
rect 66805 323715 66871 323718
rect 154246 323580 154252 323644
rect 154316 323642 154322 323644
rect 185669 323642 185735 323645
rect 154316 323640 185735 323642
rect 154316 323584 185674 323640
rect 185730 323584 185735 323640
rect 154316 323582 185735 323584
rect 154316 323580 154322 323582
rect 185669 323579 185735 323582
rect 155166 323506 155172 323508
rect 154622 323446 155172 323506
rect 154622 323204 154682 323446
rect 155166 323444 155172 323446
rect 155236 323444 155242 323508
rect 67265 322690 67331 322693
rect 67265 322688 68908 322690
rect 67265 322632 67270 322688
rect 67326 322632 68908 322688
rect 67265 322630 68908 322632
rect 67265 322627 67331 322630
rect 154982 322220 154988 322284
rect 155052 322282 155058 322284
rect 155052 322222 161490 322282
rect 155052 322220 155058 322222
rect 156045 322146 156111 322149
rect 154652 322144 156111 322146
rect 154652 322088 156050 322144
rect 156106 322088 156111 322144
rect 154652 322086 156111 322088
rect 161430 322146 161490 322222
rect 323577 322146 323643 322149
rect 161430 322144 323643 322146
rect 161430 322088 323582 322144
rect 323638 322088 323643 322144
rect 161430 322086 323643 322088
rect 156045 322083 156111 322086
rect 323577 322083 323643 322086
rect 67817 321602 67883 321605
rect 67817 321600 68908 321602
rect 67817 321544 67822 321600
rect 67878 321544 68908 321600
rect 67817 321542 68908 321544
rect 67817 321539 67883 321542
rect 65977 320244 66043 320245
rect 65926 320180 65932 320244
rect 65996 320242 66043 320244
rect 68878 320242 68938 320484
rect 154622 320378 154682 321028
rect 159214 320724 159220 320788
rect 159284 320786 159290 320788
rect 189717 320786 189783 320789
rect 159284 320784 189783 320786
rect 159284 320728 189722 320784
rect 189778 320728 189783 320784
rect 159284 320726 189783 320728
rect 159284 320724 159290 320726
rect 189717 320723 189783 320726
rect 154622 320318 161490 320378
rect 65996 320240 68938 320242
rect 66038 320184 68938 320240
rect 65996 320182 68938 320184
rect 161430 320242 161490 320318
rect 218697 320242 218763 320245
rect 161430 320240 218763 320242
rect 161430 320184 218702 320240
rect 218758 320184 218763 320240
rect 161430 320182 218763 320184
rect 65996 320180 66043 320182
rect 65977 320179 66043 320180
rect 218697 320179 218763 320182
rect 157241 319970 157307 319973
rect 154652 319968 157307 319970
rect 154652 319912 157246 319968
rect 157302 319912 157307 319968
rect 154652 319910 157307 319912
rect 157241 319907 157307 319910
rect 66253 319426 66319 319429
rect 163681 319426 163747 319429
rect 223021 319426 223087 319429
rect 66253 319424 68908 319426
rect -960 319290 480 319380
rect 66253 319368 66258 319424
rect 66314 319368 68908 319424
rect 66253 319366 68908 319368
rect 163681 319424 223087 319426
rect 163681 319368 163686 319424
rect 163742 319368 223026 319424
rect 223082 319368 223087 319424
rect 163681 319366 223087 319368
rect 66253 319363 66319 319366
rect 163681 319363 163747 319366
rect 223021 319363 223087 319366
rect 4061 319290 4127 319293
rect -960 319288 4127 319290
rect -960 319232 4066 319288
rect 4122 319232 4127 319288
rect -960 319230 4127 319232
rect -960 319140 480 319230
rect 4061 319227 4127 319230
rect 157241 318882 157307 318885
rect 154652 318880 157307 318882
rect 154652 318824 157246 318880
rect 157302 318824 157307 318880
rect 154652 318822 157307 318824
rect 157241 318819 157307 318822
rect 66345 318338 66411 318341
rect 154665 318338 154731 318341
rect 238518 318338 238524 318340
rect 66345 318336 68908 318338
rect 66345 318280 66350 318336
rect 66406 318280 68908 318336
rect 66345 318278 68908 318280
rect 154665 318336 238524 318338
rect 154665 318280 154670 318336
rect 154726 318280 238524 318336
rect 154665 318278 238524 318280
rect 66345 318275 66411 318278
rect 154665 318275 154731 318278
rect 238518 318276 238524 318278
rect 238588 318276 238594 318340
rect 155953 318066 156019 318069
rect 156597 318066 156663 318069
rect 154652 318064 156663 318066
rect 154652 318008 155958 318064
rect 156014 318008 156602 318064
rect 156658 318008 156663 318064
rect 154652 318006 156663 318008
rect 155953 318003 156019 318006
rect 156597 318003 156663 318006
rect 66253 317522 66319 317525
rect 66253 317520 68908 317522
rect 66253 317464 66258 317520
rect 66314 317464 68908 317520
rect 66253 317462 68908 317464
rect 66253 317459 66319 317462
rect 157241 316978 157307 316981
rect 154652 316976 157307 316978
rect 154652 316920 157246 316976
rect 157302 316920 157307 316976
rect 154652 316918 157307 316920
rect 157241 316915 157307 316918
rect 66662 316372 66668 316436
rect 66732 316434 66738 316436
rect 66732 316374 68908 316434
rect 66732 316372 66738 316374
rect 69422 315828 69428 315892
rect 69492 315828 69498 315892
rect 157149 315890 157215 315893
rect 154652 315888 157215 315890
rect 154652 315832 157154 315888
rect 157210 315832 157215 315888
rect 154652 315830 157215 315832
rect 66437 315346 66503 315349
rect 69430 315346 69490 315828
rect 157149 315827 157215 315830
rect 66437 315344 69490 315346
rect 66437 315288 66442 315344
rect 66498 315316 69490 315344
rect 169201 315346 169267 315349
rect 240777 315346 240843 315349
rect 169201 315344 240843 315346
rect 66498 315288 69460 315316
rect 66437 315286 69460 315288
rect 169201 315288 169206 315344
rect 169262 315288 240782 315344
rect 240838 315288 240843 315344
rect 169201 315286 240843 315288
rect 66437 315283 66503 315286
rect 169201 315283 169267 315286
rect 240777 315283 240843 315286
rect 157241 314802 157307 314805
rect 154652 314800 157307 314802
rect 154652 314744 157246 314800
rect 157302 314744 157307 314800
rect 154652 314742 157307 314744
rect 157241 314739 157307 314742
rect 66110 314196 66116 314260
rect 66180 314258 66186 314260
rect 66253 314258 66319 314261
rect 66180 314256 68908 314258
rect 66180 314200 66258 314256
rect 66314 314200 68908 314256
rect 66180 314198 68908 314200
rect 66180 314196 66186 314198
rect 66253 314195 66319 314198
rect 154430 313924 154436 313988
rect 154500 313986 154506 313988
rect 333973 313986 334039 313989
rect 154500 313984 334039 313986
rect 154500 313928 333978 313984
rect 334034 313928 334039 313984
rect 154500 313926 334039 313928
rect 154500 313924 154506 313926
rect 333973 313923 334039 313926
rect 154622 313306 154682 313684
rect 195094 313306 195100 313308
rect 154622 313246 195100 313306
rect 195094 313244 195100 313246
rect 195164 313244 195170 313308
rect 61101 313170 61167 313173
rect 61377 313170 61443 313173
rect 61101 313168 68908 313170
rect 61101 313112 61106 313168
rect 61162 313112 61382 313168
rect 61438 313112 68908 313168
rect 61101 313110 68908 313112
rect 61101 313107 61167 313110
rect 61377 313107 61443 313110
rect 157241 312626 157307 312629
rect 154652 312624 157307 312626
rect 154652 312568 157246 312624
rect 157302 312568 157307 312624
rect 154652 312566 157307 312568
rect 157241 312563 157307 312566
rect 66253 312082 66319 312085
rect 583017 312082 583083 312085
rect 583520 312082 584960 312172
rect 66253 312080 68908 312082
rect 66253 312024 66258 312080
rect 66314 312024 68908 312080
rect 66253 312022 68908 312024
rect 583017 312080 584960 312082
rect 583017 312024 583022 312080
rect 583078 312024 584960 312080
rect 583017 312022 584960 312024
rect 66253 312019 66319 312022
rect 583017 312019 583083 312022
rect 583520 311932 584960 312022
rect 157241 311538 157307 311541
rect 154652 311536 157307 311538
rect 154652 311480 157246 311536
rect 157302 311480 157307 311536
rect 154652 311478 157307 311480
rect 157241 311475 157307 311478
rect 162117 311130 162183 311133
rect 191097 311130 191163 311133
rect 162117 311128 191163 311130
rect 162117 311072 162122 311128
rect 162178 311072 191102 311128
rect 191158 311072 191163 311128
rect 162117 311070 191163 311072
rect 162117 311067 162183 311070
rect 191097 311067 191163 311070
rect 66805 310994 66871 310997
rect 66805 310992 68908 310994
rect 66805 310936 66810 310992
rect 66866 310936 68908 310992
rect 66805 310934 68908 310936
rect 66805 310931 66871 310934
rect 208485 310586 208551 310589
rect 209129 310586 209195 310589
rect 266997 310586 267063 310589
rect 208485 310584 267063 310586
rect 208485 310528 208490 310584
rect 208546 310528 209134 310584
rect 209190 310528 267002 310584
rect 267058 310528 267063 310584
rect 208485 310526 267063 310528
rect 208485 310523 208551 310526
rect 209129 310523 209195 310526
rect 266997 310523 267063 310526
rect 157241 310450 157307 310453
rect 154652 310448 157307 310450
rect 154652 310392 157246 310448
rect 157302 310392 157307 310448
rect 154652 310390 157307 310392
rect 157241 310387 157307 310390
rect 66621 309906 66687 309909
rect 66621 309904 68908 309906
rect 66621 309848 66626 309904
rect 66682 309848 68908 309904
rect 66621 309846 68908 309848
rect 66621 309843 66687 309846
rect 157149 309634 157215 309637
rect 154652 309632 157215 309634
rect 154652 309576 157154 309632
rect 157210 309576 157215 309632
rect 154652 309574 157215 309576
rect 157149 309571 157215 309574
rect 157241 309226 157307 309229
rect 302734 309226 302740 309228
rect 157241 309224 302740 309226
rect 157241 309168 157246 309224
rect 157302 309168 302740 309224
rect 157241 309166 302740 309168
rect 157241 309163 157307 309166
rect 302734 309164 302740 309166
rect 302804 309164 302810 309228
rect 67081 309090 67147 309093
rect 67081 309088 68908 309090
rect 67081 309032 67086 309088
rect 67142 309032 68908 309088
rect 67081 309030 68908 309032
rect 67081 309027 67147 309030
rect 157241 308546 157307 308549
rect 154652 308544 157307 308546
rect 154652 308488 157246 308544
rect 157302 308488 157307 308544
rect 154652 308486 157307 308488
rect 157241 308483 157307 308486
rect 159449 308410 159515 308413
rect 338113 308410 338179 308413
rect 159449 308408 338179 308410
rect 159449 308352 159454 308408
rect 159510 308352 338118 308408
rect 338174 308352 338179 308408
rect 159449 308350 338179 308352
rect 159449 308347 159515 308350
rect 338113 308347 338179 308350
rect 67173 308002 67239 308005
rect 67398 308002 67404 308004
rect 67173 308000 67404 308002
rect 67173 307944 67178 308000
rect 67234 307944 67404 308000
rect 67173 307942 67404 307944
rect 67173 307939 67239 307942
rect 67398 307940 67404 307942
rect 67468 308002 67474 308004
rect 67468 307942 68908 308002
rect 67468 307940 67474 307942
rect 67725 306914 67791 306917
rect 67725 306912 68908 306914
rect 67725 306856 67730 306912
rect 67786 306856 68908 306912
rect 67725 306854 68908 306856
rect 67725 306851 67791 306854
rect 154622 306778 154682 307428
rect 154622 306718 161490 306778
rect 161430 306506 161490 306718
rect 318057 306506 318123 306509
rect 161430 306504 318123 306506
rect 161430 306448 318062 306504
rect 318118 306448 318123 306504
rect 161430 306446 318123 306448
rect 318057 306443 318123 306446
rect 157241 306370 157307 306373
rect 154652 306368 157307 306370
rect -960 306234 480 306324
rect 154652 306312 157246 306368
rect 157302 306312 157307 306368
rect 154652 306310 157307 306312
rect 157241 306307 157307 306310
rect 3417 306234 3483 306237
rect -960 306232 3483 306234
rect -960 306176 3422 306232
rect 3478 306176 3483 306232
rect -960 306174 3483 306176
rect -960 306084 480 306174
rect 3417 306171 3483 306174
rect 67357 305826 67423 305829
rect 67357 305824 68908 305826
rect 67357 305768 67362 305824
rect 67418 305768 68908 305824
rect 67357 305766 68908 305768
rect 67357 305763 67423 305766
rect 155401 305690 155467 305693
rect 195973 305690 196039 305693
rect 155401 305688 196039 305690
rect 155401 305632 155406 305688
rect 155462 305632 195978 305688
rect 196034 305632 196039 305688
rect 155401 305630 196039 305632
rect 155401 305627 155467 305630
rect 195973 305627 196039 305630
rect 157241 305282 157307 305285
rect 154652 305280 157307 305282
rect 154652 305224 157246 305280
rect 157302 305224 157307 305280
rect 154652 305222 157307 305224
rect 157241 305219 157307 305222
rect 195973 305010 196039 305013
rect 197261 305010 197327 305013
rect 272517 305010 272583 305013
rect 195973 305008 272583 305010
rect 195973 304952 195978 305008
rect 196034 304952 197266 305008
rect 197322 304952 272522 305008
rect 272578 304952 272583 305008
rect 195973 304950 272583 304952
rect 195973 304947 196039 304950
rect 197261 304947 197327 304950
rect 272517 304947 272583 304950
rect 65517 304738 65583 304741
rect 65517 304736 68908 304738
rect 65517 304680 65522 304736
rect 65578 304680 68908 304736
rect 65517 304678 68908 304680
rect 65517 304675 65583 304678
rect 156045 304194 156111 304197
rect 154652 304192 156111 304194
rect 154652 304136 156050 304192
rect 156106 304136 156111 304192
rect 154652 304134 156111 304136
rect 156045 304131 156111 304134
rect 166441 304194 166507 304197
rect 246246 304194 246252 304196
rect 166441 304192 246252 304194
rect 166441 304136 166446 304192
rect 166502 304136 246252 304192
rect 166441 304134 246252 304136
rect 166441 304131 166507 304134
rect 246246 304132 246252 304134
rect 246316 304132 246322 304196
rect 57830 303724 57836 303788
rect 57900 303786 57906 303788
rect 57900 303726 68938 303786
rect 57900 303724 57906 303726
rect 68878 303620 68938 303726
rect 157241 303106 157307 303109
rect 154652 303104 157307 303106
rect 154652 303048 157246 303104
rect 157302 303048 157307 303104
rect 154652 303046 157307 303048
rect 157241 303043 157307 303046
rect 159357 302834 159423 302837
rect 233969 302834 234035 302837
rect 159357 302832 234035 302834
rect 159357 302776 159362 302832
rect 159418 302776 233974 302832
rect 234030 302776 234035 302832
rect 159357 302774 234035 302776
rect 159357 302771 159423 302774
rect 233969 302771 234035 302774
rect 66069 302562 66135 302565
rect 66069 302560 68908 302562
rect 66069 302504 66074 302560
rect 66130 302504 68908 302560
rect 66069 302502 68908 302504
rect 66069 302499 66135 302502
rect 176101 302290 176167 302293
rect 176561 302290 176627 302293
rect 298737 302290 298803 302293
rect 176101 302288 298803 302290
rect 176101 302232 176106 302288
rect 176162 302232 176566 302288
rect 176622 302232 298742 302288
rect 298798 302232 298803 302288
rect 176101 302230 298803 302232
rect 176101 302227 176167 302230
rect 176561 302227 176627 302230
rect 298737 302227 298803 302230
rect 66805 301474 66871 301477
rect 154622 301474 154682 301988
rect 66805 301472 68908 301474
rect 66805 301416 66810 301472
rect 66866 301416 68908 301472
rect 66805 301414 68908 301416
rect 154622 301414 161490 301474
rect 66805 301411 66871 301414
rect 154622 300930 154682 301172
rect 161430 301066 161490 301414
rect 188286 301066 188292 301068
rect 161430 301006 188292 301066
rect 188286 301004 188292 301006
rect 188356 301004 188362 301068
rect 316677 300930 316743 300933
rect 154622 300928 316743 300930
rect 154622 300872 316682 300928
rect 316738 300872 316743 300928
rect 154622 300870 316743 300872
rect 316677 300867 316743 300870
rect 66437 300658 66503 300661
rect 66437 300656 68908 300658
rect 66437 300600 66442 300656
rect 66498 300600 68908 300656
rect 66437 300598 68908 300600
rect 66437 300595 66503 300598
rect 154622 299706 154682 300084
rect 244038 299706 244044 299708
rect 154622 299646 244044 299706
rect 244038 299644 244044 299646
rect 244108 299644 244114 299708
rect 66805 299570 66871 299573
rect 240777 299570 240843 299573
rect 583109 299570 583175 299573
rect 66805 299568 68908 299570
rect 66805 299512 66810 299568
rect 66866 299512 68908 299568
rect 66805 299510 68908 299512
rect 240777 299568 583175 299570
rect 240777 299512 240782 299568
rect 240838 299512 583114 299568
rect 583170 299512 583175 299568
rect 240777 299510 583175 299512
rect 66805 299507 66871 299510
rect 240777 299507 240843 299510
rect 583109 299507 583175 299510
rect 164141 299434 164207 299437
rect 171225 299434 171291 299437
rect 172421 299434 172487 299437
rect 164141 299432 172487 299434
rect 164141 299376 164146 299432
rect 164202 299376 171230 299432
rect 171286 299376 172426 299432
rect 172482 299376 172487 299432
rect 164141 299374 172487 299376
rect 164141 299371 164207 299374
rect 171225 299371 171291 299374
rect 172421 299371 172487 299374
rect 157241 299026 157307 299029
rect 154652 299024 157307 299026
rect 154652 298968 157246 299024
rect 157302 298968 157307 299024
rect 154652 298966 157307 298968
rect 157241 298963 157307 298966
rect 172421 298754 172487 298757
rect 213637 298754 213703 298757
rect 172421 298752 213703 298754
rect 172421 298696 172426 298752
rect 172482 298696 213642 298752
rect 213698 298696 213703 298752
rect 172421 298694 213703 298696
rect 172421 298691 172487 298694
rect 213637 298691 213703 298694
rect 225597 298754 225663 298757
rect 235533 298754 235599 298757
rect 225597 298752 235599 298754
rect 225597 298696 225602 298752
rect 225658 298696 235538 298752
rect 235594 298696 235599 298752
rect 225597 298694 235599 298696
rect 225597 298691 225663 298694
rect 235533 298691 235599 298694
rect 583385 298754 583451 298757
rect 583520 298754 584960 298844
rect 583385 298752 584960 298754
rect 583385 298696 583390 298752
rect 583446 298696 584960 298752
rect 583385 298694 584960 298696
rect 583385 298691 583451 298694
rect 583520 298604 584960 298694
rect 67541 298482 67607 298485
rect 67541 298480 68908 298482
rect 67541 298424 67546 298480
rect 67602 298424 68908 298480
rect 67541 298422 68908 298424
rect 67541 298419 67607 298422
rect 206277 298210 206343 298213
rect 582925 298210 582991 298213
rect 206277 298208 582991 298210
rect 206277 298152 206282 298208
rect 206338 298152 582930 298208
rect 582986 298152 582991 298208
rect 206277 298150 582991 298152
rect 206277 298147 206343 298150
rect 582925 298147 582991 298150
rect 235257 298074 235323 298077
rect 236177 298074 236243 298077
rect 235257 298072 236243 298074
rect 235257 298016 235262 298072
rect 235318 298016 236182 298072
rect 236238 298016 236243 298072
rect 235257 298014 236243 298016
rect 235257 298011 235323 298014
rect 236177 298011 236243 298014
rect 156413 297938 156479 297941
rect 154652 297936 156479 297938
rect 154652 297880 156418 297936
rect 156474 297880 156479 297936
rect 154652 297878 156479 297880
rect 156413 297875 156479 297878
rect 177573 297530 177639 297533
rect 214046 297530 214052 297532
rect 177573 297528 214052 297530
rect 177573 297472 177578 297528
rect 177634 297472 214052 297528
rect 177573 297470 214052 297472
rect 177573 297467 177639 297470
rect 214046 297468 214052 297470
rect 214116 297468 214122 297532
rect 66621 297394 66687 297397
rect 165705 297394 165771 297397
rect 256785 297394 256851 297397
rect 66621 297392 68908 297394
rect 66621 297336 66626 297392
rect 66682 297336 68908 297392
rect 66621 297334 68908 297336
rect 165705 297392 256851 297394
rect 165705 297336 165710 297392
rect 165766 297336 256790 297392
rect 256846 297336 256851 297392
rect 165705 297334 256851 297336
rect 66621 297331 66687 297334
rect 165705 297331 165771 297334
rect 256785 297331 256851 297334
rect 156689 296850 156755 296853
rect 154652 296848 156755 296850
rect 154652 296792 156694 296848
rect 156750 296792 156755 296848
rect 154652 296790 156755 296792
rect 156689 296787 156755 296790
rect 236177 296850 236243 296853
rect 574737 296850 574803 296853
rect 236177 296848 574803 296850
rect 236177 296792 236182 296848
rect 236238 296792 574742 296848
rect 574798 296792 574803 296848
rect 236177 296790 574803 296792
rect 236177 296787 236243 296790
rect 574737 296787 574803 296790
rect 66437 296306 66503 296309
rect 66437 296304 68908 296306
rect 66437 296248 66442 296304
rect 66498 296248 68908 296304
rect 66437 296246 68908 296248
rect 66437 296243 66503 296246
rect 69422 295428 69428 295492
rect 69492 295428 69498 295492
rect 67541 295218 67607 295221
rect 69430 295218 69490 295428
rect 154622 295354 154682 295732
rect 220169 295490 220235 295493
rect 220721 295490 220787 295493
rect 268377 295490 268443 295493
rect 220169 295488 268443 295490
rect 220169 295432 220174 295488
rect 220230 295432 220726 295488
rect 220782 295432 268382 295488
rect 268438 295432 268443 295488
rect 220169 295430 268443 295432
rect 220169 295427 220235 295430
rect 220721 295427 220787 295430
rect 268377 295427 268443 295430
rect 160134 295354 160140 295356
rect 154622 295294 160140 295354
rect 160134 295292 160140 295294
rect 160204 295354 160210 295356
rect 160829 295354 160895 295357
rect 160204 295352 160895 295354
rect 160204 295296 160834 295352
rect 160890 295296 160895 295352
rect 160204 295294 160895 295296
rect 160204 295292 160210 295294
rect 160829 295291 160895 295294
rect 184381 295354 184447 295357
rect 224309 295354 224375 295357
rect 184381 295352 224375 295354
rect 184381 295296 184386 295352
rect 184442 295296 224314 295352
rect 224370 295296 224375 295352
rect 184381 295294 224375 295296
rect 184381 295291 184447 295294
rect 224309 295291 224375 295294
rect 233693 295354 233759 295357
rect 233969 295354 234035 295357
rect 583661 295354 583727 295357
rect 233693 295352 583727 295354
rect 233693 295296 233698 295352
rect 233754 295296 233974 295352
rect 234030 295296 583666 295352
rect 583722 295296 583727 295352
rect 233693 295294 583727 295296
rect 233693 295291 233759 295294
rect 233969 295291 234035 295294
rect 583661 295291 583727 295294
rect 67541 295216 69490 295218
rect 67541 295160 67546 295216
rect 67602 295188 69490 295216
rect 67602 295160 69460 295188
rect 67541 295158 69460 295160
rect 67541 295155 67607 295158
rect 156321 294674 156387 294677
rect 154652 294672 156387 294674
rect 154652 294616 156326 294672
rect 156382 294616 156387 294672
rect 154652 294614 156387 294616
rect 156321 294611 156387 294614
rect 242249 294674 242315 294677
rect 248689 294674 248755 294677
rect 242249 294672 248755 294674
rect 242249 294616 242254 294672
rect 242310 294616 248694 294672
rect 248750 294616 248755 294672
rect 242249 294614 248755 294616
rect 242249 294611 242315 294614
rect 248689 294611 248755 294614
rect 240225 294538 240291 294541
rect 583753 294538 583819 294541
rect 240225 294536 583819 294538
rect 240225 294480 240230 294536
rect 240286 294480 583758 294536
rect 583814 294480 583819 294536
rect 240225 294478 583819 294480
rect 240225 294475 240291 294478
rect 583753 294475 583819 294478
rect 66805 294130 66871 294133
rect 215293 294130 215359 294133
rect 229737 294130 229803 294133
rect 66805 294128 68908 294130
rect 66805 294072 66810 294128
rect 66866 294072 68908 294128
rect 66805 294070 68908 294072
rect 215293 294128 229803 294130
rect 215293 294072 215298 294128
rect 215354 294072 229742 294128
rect 229798 294072 229803 294128
rect 215293 294070 229803 294072
rect 66805 294067 66871 294070
rect 215293 294067 215359 294070
rect 229737 294067 229803 294070
rect 239029 294130 239095 294133
rect 240225 294130 240291 294133
rect 239029 294128 240291 294130
rect 239029 294072 239034 294128
rect 239090 294072 240230 294128
rect 240286 294072 240291 294128
rect 239029 294070 240291 294072
rect 239029 294067 239095 294070
rect 240225 294067 240291 294070
rect 177481 293994 177547 293997
rect 251449 293994 251515 293997
rect 177481 293992 251515 293994
rect 177481 293936 177486 293992
rect 177542 293936 251454 293992
rect 251510 293936 251515 293992
rect 177481 293934 251515 293936
rect 177481 293931 177547 293934
rect 251449 293931 251515 293934
rect 156505 293586 156571 293589
rect 154652 293584 156571 293586
rect 154652 293528 156510 293584
rect 156566 293528 156571 293584
rect 154652 293526 156571 293528
rect 156505 293523 156571 293526
rect -960 293178 480 293268
rect 2773 293178 2839 293181
rect -960 293176 2839 293178
rect -960 293120 2778 293176
rect 2834 293120 2839 293176
rect -960 293118 2839 293120
rect -960 293028 480 293118
rect 2773 293115 2839 293118
rect 159357 293178 159423 293181
rect 215293 293178 215359 293181
rect 159357 293176 215359 293178
rect 159357 293120 159362 293176
rect 159418 293120 215298 293176
rect 215354 293120 215359 293176
rect 159357 293118 215359 293120
rect 159357 293115 159423 293118
rect 215293 293115 215359 293118
rect 66989 293042 67055 293045
rect 66989 293040 68908 293042
rect 66989 292984 66994 293040
rect 67050 292984 68908 293040
rect 66989 292982 68908 292984
rect 66989 292979 67055 292982
rect 210509 292906 210575 292909
rect 216949 292906 217015 292909
rect 210509 292904 217015 292906
rect 210509 292848 210514 292904
rect 210570 292848 216954 292904
rect 217010 292848 217015 292904
rect 210509 292846 217015 292848
rect 210509 292843 210575 292846
rect 216949 292843 217015 292846
rect 157241 292770 157307 292773
rect 252553 292770 252619 292773
rect 154652 292768 157307 292770
rect 154652 292712 157246 292768
rect 157302 292712 157307 292768
rect 154652 292710 157307 292712
rect 157241 292707 157307 292710
rect 197126 292710 200130 292770
rect 191189 292634 191255 292637
rect 191741 292634 191807 292637
rect 197126 292634 197186 292710
rect 191189 292632 197186 292634
rect 191189 292576 191194 292632
rect 191250 292576 191746 292632
rect 191802 292576 197186 292632
rect 191189 292574 197186 292576
rect 197261 292634 197327 292637
rect 197854 292634 197860 292636
rect 197261 292632 197860 292634
rect 197261 292576 197266 292632
rect 197322 292576 197860 292632
rect 197261 292574 197860 292576
rect 191189 292571 191255 292574
rect 191741 292571 191807 292574
rect 197261 292571 197327 292574
rect 197854 292572 197860 292574
rect 197924 292572 197930 292636
rect 200070 292634 200130 292710
rect 216814 292768 252619 292770
rect 216814 292712 252558 292768
rect 252614 292712 252619 292768
rect 216814 292710 252619 292712
rect 209957 292634 210023 292637
rect 200070 292632 210023 292634
rect 200070 292576 209962 292632
rect 210018 292576 210023 292632
rect 200070 292574 210023 292576
rect 209957 292571 210023 292574
rect 215293 292634 215359 292637
rect 215937 292634 216003 292637
rect 216814 292634 216874 292710
rect 252553 292707 252619 292710
rect 215293 292632 216874 292634
rect 215293 292576 215298 292632
rect 215354 292576 215942 292632
rect 215998 292576 216874 292632
rect 215293 292574 216874 292576
rect 216949 292634 217015 292637
rect 251541 292634 251607 292637
rect 216949 292632 251607 292634
rect 216949 292576 216954 292632
rect 217010 292576 251546 292632
rect 251602 292576 251607 292632
rect 216949 292574 251607 292576
rect 215293 292571 215359 292574
rect 215937 292571 216003 292574
rect 216949 292571 217015 292574
rect 251541 292571 251607 292574
rect 66897 292226 66963 292229
rect 66897 292224 68908 292226
rect 66897 292168 66902 292224
rect 66958 292168 68908 292224
rect 66897 292166 68908 292168
rect 66897 292163 66963 292166
rect 213821 291818 213887 291821
rect 582465 291818 582531 291821
rect 213821 291816 582531 291818
rect 213821 291760 213826 291816
rect 213882 291760 582470 291816
rect 582526 291760 582531 291816
rect 213821 291758 582531 291760
rect 213821 291755 213887 291758
rect 582465 291755 582531 291758
rect 156045 291682 156111 291685
rect 154652 291680 156111 291682
rect 154652 291624 156050 291680
rect 156106 291624 156111 291680
rect 154652 291622 156111 291624
rect 156045 291619 156111 291622
rect 199326 291484 199332 291548
rect 199396 291546 199402 291548
rect 232773 291546 232839 291549
rect 199396 291544 232839 291546
rect 199396 291488 232778 291544
rect 232834 291488 232839 291544
rect 199396 291486 232839 291488
rect 199396 291484 199402 291486
rect 232773 291483 232839 291486
rect 174629 291410 174695 291413
rect 213453 291410 213519 291413
rect 213821 291410 213887 291413
rect 174629 291408 213887 291410
rect 174629 291352 174634 291408
rect 174690 291352 213458 291408
rect 213514 291352 213826 291408
rect 213882 291352 213887 291408
rect 174629 291350 213887 291352
rect 174629 291347 174695 291350
rect 213453 291347 213519 291350
rect 213821 291347 213887 291350
rect 164877 291274 164943 291277
rect 249977 291274 250043 291277
rect 164877 291272 250043 291274
rect 164877 291216 164882 291272
rect 164938 291216 249982 291272
rect 250038 291216 250043 291272
rect 164877 291214 250043 291216
rect 164877 291211 164943 291214
rect 249977 291211 250043 291214
rect 66805 291138 66871 291141
rect 66805 291136 68908 291138
rect 66805 291080 66810 291136
rect 66866 291080 68908 291136
rect 66805 291078 68908 291080
rect 66805 291075 66871 291078
rect 156454 291076 156460 291140
rect 156524 291138 156530 291140
rect 156781 291138 156847 291141
rect 156524 291136 156847 291138
rect 156524 291080 156786 291136
rect 156842 291080 156847 291136
rect 156524 291078 156847 291080
rect 156524 291076 156530 291078
rect 156781 291075 156847 291078
rect 193949 291138 194015 291141
rect 194501 291138 194567 291141
rect 193949 291136 194567 291138
rect 193949 291080 193954 291136
rect 194010 291080 194506 291136
rect 194562 291080 194567 291136
rect 193949 291078 194567 291080
rect 193949 291075 194015 291078
rect 194501 291075 194567 291078
rect 200757 291138 200823 291141
rect 582557 291138 582623 291141
rect 200757 291136 582623 291138
rect 200757 291080 200762 291136
rect 200818 291080 582562 291136
rect 582618 291080 582623 291136
rect 200757 291078 582623 291080
rect 200757 291075 200823 291078
rect 582557 291075 582623 291078
rect 157241 290594 157307 290597
rect 154652 290592 157307 290594
rect 154652 290536 157246 290592
rect 157302 290536 157307 290592
rect 154652 290534 157307 290536
rect 157241 290531 157307 290534
rect 213637 290458 213703 290461
rect 227897 290458 227963 290461
rect 213637 290456 227963 290458
rect 213637 290400 213642 290456
rect 213698 290400 227902 290456
rect 227958 290400 227963 290456
rect 213637 290398 227963 290400
rect 213637 290395 213703 290398
rect 227897 290395 227963 290398
rect 156781 290186 156847 290189
rect 247217 290186 247283 290189
rect 156781 290184 247283 290186
rect 156781 290128 156786 290184
rect 156842 290128 247222 290184
rect 247278 290128 247283 290184
rect 156781 290126 247283 290128
rect 156781 290123 156847 290126
rect 247217 290123 247283 290126
rect 66805 290050 66871 290053
rect 194501 290050 194567 290053
rect 203149 290050 203215 290053
rect 66805 290048 68908 290050
rect 66805 289992 66810 290048
rect 66866 289992 68908 290048
rect 66805 289990 68908 289992
rect 194501 290048 203215 290050
rect 194501 289992 194506 290048
rect 194562 289992 203154 290048
rect 203210 289992 203215 290048
rect 194501 289990 203215 289992
rect 66805 289987 66871 289990
rect 194501 289987 194567 289990
rect 203149 289987 203215 289990
rect 157241 289506 157307 289509
rect 154652 289504 157307 289506
rect 154652 289448 157246 289504
rect 157302 289448 157307 289504
rect 154652 289446 157307 289448
rect 157241 289443 157307 289446
rect 66713 288962 66779 288965
rect 66713 288960 68908 288962
rect 66713 288904 66718 288960
rect 66774 288904 68908 288960
rect 66713 288902 68908 288904
rect 66713 288899 66779 288902
rect 197077 288826 197143 288829
rect 230749 288826 230815 288829
rect 197077 288824 230815 288826
rect 197077 288768 197082 288824
rect 197138 288768 230754 288824
rect 230810 288768 230815 288824
rect 197077 288766 230815 288768
rect 197077 288763 197143 288766
rect 230749 288763 230815 288766
rect 181529 288690 181595 288693
rect 217317 288690 217383 288693
rect 181529 288688 217383 288690
rect 181529 288632 181534 288688
rect 181590 288632 217322 288688
rect 217378 288632 217383 288688
rect 181529 288630 217383 288632
rect 181529 288627 181595 288630
rect 217317 288627 217383 288630
rect 226977 288690 227043 288693
rect 249742 288690 249748 288692
rect 226977 288688 249748 288690
rect 226977 288632 226982 288688
rect 227038 288632 249748 288688
rect 226977 288630 249748 288632
rect 226977 288627 227043 288630
rect 249742 288628 249748 288630
rect 249812 288628 249818 288692
rect 202229 288554 202295 288557
rect 285622 288554 285628 288556
rect 202229 288552 285628 288554
rect 202229 288496 202234 288552
rect 202290 288496 285628 288552
rect 202229 288494 285628 288496
rect 202229 288491 202295 288494
rect 285622 288492 285628 288494
rect 285692 288492 285698 288556
rect 157241 288418 157307 288421
rect 154652 288416 157307 288418
rect 154652 288360 157246 288416
rect 157302 288360 157307 288416
rect 154652 288358 157307 288360
rect 157241 288355 157307 288358
rect 66621 287874 66687 287877
rect 66621 287872 68908 287874
rect 66621 287816 66626 287872
rect 66682 287816 68908 287872
rect 66621 287814 68908 287816
rect 66621 287811 66687 287814
rect 211981 287602 212047 287605
rect 284334 287602 284340 287604
rect 200070 287600 284340 287602
rect 200070 287544 211986 287600
rect 212042 287544 284340 287600
rect 200070 287542 284340 287544
rect 198181 287466 198247 287469
rect 200070 287466 200130 287542
rect 211981 287539 212047 287542
rect 284334 287540 284340 287542
rect 284404 287540 284410 287604
rect 238109 287466 238175 287469
rect 260097 287466 260163 287469
rect 198181 287464 200130 287466
rect 198181 287408 198186 287464
rect 198242 287408 200130 287464
rect 198181 287406 200130 287408
rect 219390 287464 260163 287466
rect 219390 287408 238114 287464
rect 238170 287408 260102 287464
rect 260158 287408 260163 287464
rect 219390 287406 260163 287408
rect 198181 287403 198247 287406
rect 174721 287330 174787 287333
rect 219390 287330 219450 287406
rect 238109 287403 238175 287406
rect 260097 287403 260163 287406
rect 239949 287330 240015 287333
rect 288433 287330 288499 287333
rect 174721 287328 219450 287330
rect 154622 287194 154682 287300
rect 174721 287272 174726 287328
rect 174782 287272 219450 287328
rect 174721 287270 219450 287272
rect 238710 287328 288499 287330
rect 238710 287272 239954 287328
rect 240010 287272 288438 287328
rect 288494 287272 288499 287328
rect 238710 287270 288499 287272
rect 174721 287267 174787 287270
rect 173014 287194 173020 287196
rect 154622 287134 173020 287194
rect 173014 287132 173020 287134
rect 173084 287132 173090 287196
rect 229737 287058 229803 287061
rect 238710 287058 238770 287270
rect 239949 287267 240015 287270
rect 288433 287267 288499 287270
rect 229737 287056 238770 287058
rect 229737 287000 229742 287056
rect 229798 287000 238770 287056
rect 229737 286998 238770 287000
rect 229737 286995 229803 286998
rect 66805 286786 66871 286789
rect 66805 286784 68908 286786
rect 66805 286728 66810 286784
rect 66866 286728 68908 286784
rect 66805 286726 68908 286728
rect 66805 286723 66871 286726
rect 215201 286650 215267 286653
rect 221549 286650 221615 286653
rect 215201 286648 221615 286650
rect 215201 286592 215206 286648
rect 215262 286592 221554 286648
rect 221610 286592 221615 286648
rect 215201 286590 221615 286592
rect 215201 286587 215267 286590
rect 221549 286587 221615 286590
rect 228357 286650 228423 286653
rect 230381 286650 230447 286653
rect 228357 286648 230447 286650
rect 228357 286592 228362 286648
rect 228418 286592 230386 286648
rect 230442 286592 230447 286648
rect 228357 286590 230447 286592
rect 228357 286587 228423 286590
rect 230381 286587 230447 286590
rect 159214 286316 159220 286380
rect 159284 286378 159290 286380
rect 164877 286378 164943 286381
rect 159284 286376 164943 286378
rect 159284 286320 164882 286376
rect 164938 286320 164943 286376
rect 159284 286318 164943 286320
rect 159284 286316 159290 286318
rect 164877 286315 164943 286318
rect 188429 286378 188495 286381
rect 195462 286378 195468 286380
rect 188429 286376 195468 286378
rect 188429 286320 188434 286376
rect 188490 286320 195468 286376
rect 188429 286318 195468 286320
rect 188429 286315 188495 286318
rect 195462 286316 195468 286318
rect 195532 286316 195538 286380
rect 236729 286378 236795 286381
rect 236729 286376 238770 286378
rect 236729 286320 236734 286376
rect 236790 286320 238770 286376
rect 236729 286318 238770 286320
rect 236729 286315 236795 286318
rect 157057 286242 157123 286245
rect 154652 286240 157123 286242
rect 154652 286184 157062 286240
rect 157118 286184 157123 286240
rect 154652 286182 157123 286184
rect 157057 286179 157123 286182
rect 190361 286106 190427 286109
rect 219157 286106 219223 286109
rect 190361 286104 219223 286106
rect 190361 286048 190366 286104
rect 190422 286048 219162 286104
rect 219218 286048 219223 286104
rect 190361 286046 219223 286048
rect 190361 286043 190427 286046
rect 219157 286043 219223 286046
rect 178861 285834 178927 285837
rect 203701 285834 203767 285837
rect 178861 285832 203767 285834
rect 178861 285776 178866 285832
rect 178922 285776 203706 285832
rect 203762 285776 203767 285832
rect 178861 285774 203767 285776
rect 178861 285771 178927 285774
rect 203701 285771 203767 285774
rect 210734 285772 210740 285836
rect 210804 285834 210810 285836
rect 220077 285834 220143 285837
rect 210804 285832 220143 285834
rect 210804 285776 220082 285832
rect 220138 285776 220143 285832
rect 210804 285774 220143 285776
rect 210804 285772 210810 285774
rect 220077 285771 220143 285774
rect 223481 285834 223547 285837
rect 226517 285834 226583 285837
rect 223481 285832 226583 285834
rect 223481 285776 223486 285832
rect 223542 285776 226522 285832
rect 226578 285776 226583 285832
rect 223481 285774 226583 285776
rect 238710 285834 238770 286318
rect 239581 285834 239647 285837
rect 262857 285834 262923 285837
rect 238710 285832 262923 285834
rect 238710 285776 239586 285832
rect 239642 285776 262862 285832
rect 262918 285776 262923 285832
rect 238710 285774 262923 285776
rect 223481 285771 223547 285774
rect 226517 285771 226583 285774
rect 239581 285771 239647 285774
rect 262857 285771 262923 285774
rect 66989 285698 67055 285701
rect 195329 285698 195395 285701
rect 200757 285698 200823 285701
rect 66989 285696 68908 285698
rect 66989 285640 66994 285696
rect 67050 285640 68908 285696
rect 66989 285638 68908 285640
rect 195329 285696 200823 285698
rect 195329 285640 195334 285696
rect 195390 285640 200762 285696
rect 200818 285640 200823 285696
rect 195329 285638 200823 285640
rect 66989 285635 67055 285638
rect 195329 285635 195395 285638
rect 200757 285635 200823 285638
rect 201401 285698 201467 285701
rect 206093 285698 206159 285701
rect 201401 285696 206159 285698
rect 201401 285640 201406 285696
rect 201462 285640 206098 285696
rect 206154 285640 206159 285696
rect 201401 285638 206159 285640
rect 201401 285635 201467 285638
rect 206093 285635 206159 285638
rect 223614 285636 223620 285700
rect 223684 285698 223690 285700
rect 223941 285698 224007 285701
rect 223684 285696 224007 285698
rect 223684 285640 223946 285696
rect 224002 285640 224007 285696
rect 223684 285638 224007 285640
rect 223684 285636 223690 285638
rect 223941 285635 224007 285638
rect 224309 285698 224375 285701
rect 225413 285698 225479 285701
rect 224309 285696 225479 285698
rect 224309 285640 224314 285696
rect 224370 285640 225418 285696
rect 225474 285640 225479 285696
rect 224309 285638 225479 285640
rect 224309 285635 224375 285638
rect 225413 285635 225479 285638
rect 232497 285698 232563 285701
rect 234613 285698 234679 285701
rect 232497 285696 234679 285698
rect 232497 285640 232502 285696
rect 232558 285640 234618 285696
rect 234674 285640 234679 285696
rect 232497 285638 234679 285640
rect 232497 285635 232563 285638
rect 234613 285635 234679 285638
rect 235993 285698 236059 285701
rect 236494 285698 236500 285700
rect 235993 285696 236500 285698
rect 235993 285640 235998 285696
rect 236054 285640 236500 285696
rect 235993 285638 236500 285640
rect 235993 285635 236059 285638
rect 236494 285636 236500 285638
rect 236564 285636 236570 285700
rect 240777 285698 240843 285701
rect 243813 285698 243879 285701
rect 310513 285698 310579 285701
rect 240777 285696 243879 285698
rect 240777 285640 240782 285696
rect 240838 285640 243818 285696
rect 243874 285640 243879 285696
rect 240777 285638 243879 285640
rect 240777 285635 240843 285638
rect 243813 285635 243879 285638
rect 244046 285696 310579 285698
rect 244046 285640 310518 285696
rect 310574 285640 310579 285696
rect 244046 285638 310579 285640
rect 157149 285562 157215 285565
rect 167637 285562 167703 285565
rect 157149 285560 167703 285562
rect 157149 285504 157154 285560
rect 157210 285504 167642 285560
rect 167698 285504 167703 285560
rect 157149 285502 167703 285504
rect 157149 285499 157215 285502
rect 167637 285499 167703 285502
rect 242157 285562 242223 285565
rect 242617 285562 242683 285565
rect 244046 285562 244106 285638
rect 310513 285635 310579 285638
rect 242157 285560 244106 285562
rect 242157 285504 242162 285560
rect 242218 285504 242622 285560
rect 242678 285504 244106 285560
rect 242157 285502 244106 285504
rect 242157 285499 242223 285502
rect 242617 285499 242683 285502
rect 583520 285276 584960 285516
rect 156413 285154 156479 285157
rect 154652 285152 156479 285154
rect 154652 285096 156418 285152
rect 156474 285096 156479 285152
rect 154652 285094 156479 285096
rect 156413 285091 156479 285094
rect 185761 284882 185827 284885
rect 204989 284882 205055 284885
rect 185761 284880 205055 284882
rect 185761 284824 185766 284880
rect 185822 284824 204994 284880
rect 205050 284824 205055 284880
rect 185761 284822 205055 284824
rect 185761 284819 185827 284822
rect 204989 284819 205055 284822
rect 67081 284610 67147 284613
rect 67081 284608 68908 284610
rect 67081 284552 67086 284608
rect 67142 284552 68908 284608
rect 67081 284550 68908 284552
rect 67081 284547 67147 284550
rect 198774 284548 198780 284612
rect 198844 284610 198850 284612
rect 200021 284610 200087 284613
rect 198844 284608 200087 284610
rect 198844 284552 200026 284608
rect 200082 284552 200087 284608
rect 198844 284550 200087 284552
rect 198844 284548 198850 284550
rect 200021 284547 200087 284550
rect 200614 284548 200620 284612
rect 200684 284610 200690 284612
rect 200757 284610 200823 284613
rect 200684 284608 200823 284610
rect 200684 284552 200762 284608
rect 200818 284552 200823 284608
rect 200684 284550 200823 284552
rect 200684 284548 200690 284550
rect 200757 284547 200823 284550
rect 216765 284610 216831 284613
rect 237414 284610 237420 284612
rect 216765 284608 237420 284610
rect 216765 284552 216770 284608
rect 216826 284552 237420 284608
rect 216765 284550 237420 284552
rect 216765 284547 216831 284550
rect 237414 284548 237420 284550
rect 237484 284548 237490 284612
rect 169201 284474 169267 284477
rect 204253 284474 204319 284477
rect 169201 284472 204319 284474
rect 169201 284416 169206 284472
rect 169262 284416 204258 284472
rect 204314 284416 204319 284472
rect 169201 284414 204319 284416
rect 169201 284411 169267 284414
rect 204253 284411 204319 284414
rect 212349 284474 212415 284477
rect 264237 284474 264303 284477
rect 212349 284472 264303 284474
rect 212349 284416 212354 284472
rect 212410 284416 264242 284472
rect 264298 284416 264303 284472
rect 212349 284414 264303 284416
rect 212349 284411 212415 284414
rect 264237 284411 264303 284414
rect 157149 284338 157215 284341
rect 154652 284336 157215 284338
rect 154652 284280 157154 284336
rect 157210 284280 157215 284336
rect 154652 284278 157215 284280
rect 157149 284275 157215 284278
rect 198733 284338 198799 284341
rect 210877 284338 210943 284341
rect 198733 284336 210943 284338
rect 198733 284280 198738 284336
rect 198794 284280 210882 284336
rect 210938 284280 210943 284336
rect 198733 284278 210943 284280
rect 198733 284275 198799 284278
rect 210877 284275 210943 284278
rect 214741 284338 214807 284341
rect 304257 284338 304323 284341
rect 214741 284336 304323 284338
rect 214741 284280 214746 284336
rect 214802 284280 304262 284336
rect 304318 284280 304323 284336
rect 214741 284278 304323 284280
rect 214741 284275 214807 284278
rect 304257 284275 304323 284278
rect 201953 284066 202019 284069
rect 180750 284064 202019 284066
rect 180750 284008 201958 284064
rect 202014 284008 202019 284064
rect 180750 284006 202019 284008
rect 66110 283732 66116 283796
rect 66180 283794 66186 283796
rect 66180 283734 68908 283794
rect 66180 283732 66186 283734
rect 154246 283460 154252 283524
rect 154316 283522 154322 283524
rect 180750 283522 180810 284006
rect 201953 284003 202019 284006
rect 220721 284066 220787 284069
rect 222694 284066 222700 284068
rect 220721 284064 222700 284066
rect 220721 284008 220726 284064
rect 220782 284008 222700 284064
rect 220721 284006 222700 284008
rect 220721 284003 220787 284006
rect 222694 284004 222700 284006
rect 222764 284004 222770 284068
rect 223757 284066 223823 284069
rect 226926 284066 226932 284068
rect 223757 284064 226932 284066
rect 223757 284008 223762 284064
rect 223818 284008 226932 284064
rect 223757 284006 226932 284008
rect 223757 284003 223823 284006
rect 226926 284004 226932 284006
rect 226996 284004 227002 284068
rect 243629 284066 243695 284069
rect 244089 284066 244155 284069
rect 243629 284064 244155 284066
rect 243629 284008 243634 284064
rect 243690 284008 244094 284064
rect 244150 284008 244155 284064
rect 243629 284006 244155 284008
rect 243629 284003 243695 284006
rect 244089 284003 244155 284006
rect 205357 283932 205423 283933
rect 205357 283930 205404 283932
rect 205312 283928 205404 283930
rect 205312 283872 205362 283928
rect 205312 283870 205404 283872
rect 205357 283868 205404 283870
rect 205468 283868 205474 283932
rect 211613 283930 211679 283933
rect 214465 283932 214531 283933
rect 215937 283932 216003 283933
rect 212390 283930 212396 283932
rect 211613 283928 212396 283930
rect 211613 283872 211618 283928
rect 211674 283872 212396 283928
rect 211613 283870 212396 283872
rect 205357 283867 205423 283868
rect 211613 283867 211679 283870
rect 212390 283868 212396 283870
rect 212460 283868 212466 283932
rect 214414 283930 214420 283932
rect 214374 283870 214420 283930
rect 214484 283928 214531 283932
rect 215886 283930 215892 283932
rect 214526 283872 214531 283928
rect 214414 283868 214420 283870
rect 214484 283868 214531 283872
rect 215846 283870 215892 283930
rect 215956 283928 216003 283932
rect 215998 283872 216003 283928
rect 215886 283868 215892 283870
rect 215956 283868 216003 283872
rect 216622 283868 216628 283932
rect 216692 283930 216698 283932
rect 217409 283930 217475 283933
rect 221273 283932 221339 283933
rect 216692 283928 217475 283930
rect 216692 283872 217414 283928
rect 217470 283872 217475 283928
rect 216692 283870 217475 283872
rect 216692 283868 216698 283870
rect 214465 283867 214531 283868
rect 215937 283867 216003 283868
rect 217409 283867 217475 283870
rect 221222 283868 221228 283932
rect 221292 283930 221339 283932
rect 224677 283932 224743 283933
rect 224677 283930 224724 283932
rect 221292 283928 221384 283930
rect 221334 283872 221384 283928
rect 221292 283870 221384 283872
rect 224632 283928 224724 283930
rect 224632 283872 224682 283928
rect 224632 283870 224724 283872
rect 221292 283868 221339 283870
rect 221273 283867 221339 283868
rect 224677 283868 224724 283870
rect 224788 283868 224794 283932
rect 225229 283930 225295 283933
rect 226190 283930 226196 283932
rect 225229 283928 226196 283930
rect 225229 283872 225234 283928
rect 225290 283872 226196 283928
rect 225229 283870 226196 283872
rect 224677 283867 224743 283868
rect 225229 283867 225295 283870
rect 226190 283868 226196 283870
rect 226260 283868 226266 283932
rect 230105 283930 230171 283933
rect 230238 283930 230244 283932
rect 230105 283928 230244 283930
rect 230105 283872 230110 283928
rect 230166 283872 230244 283928
rect 230105 283870 230244 283872
rect 230105 283867 230171 283870
rect 230238 283868 230244 283870
rect 230308 283868 230314 283932
rect 231577 283930 231643 283933
rect 231710 283930 231716 283932
rect 231577 283928 231716 283930
rect 231577 283872 231582 283928
rect 231638 283872 231716 283928
rect 231577 283870 231716 283872
rect 231577 283867 231643 283870
rect 231710 283868 231716 283870
rect 231780 283868 231786 283932
rect 236494 283868 236500 283932
rect 236564 283930 236570 283932
rect 236729 283930 236795 283933
rect 236564 283928 236795 283930
rect 236564 283872 236734 283928
rect 236790 283872 236795 283928
rect 236564 283870 236795 283872
rect 236564 283868 236570 283870
rect 236729 283867 236795 283870
rect 238661 283930 238727 283933
rect 240358 283930 240364 283932
rect 238661 283928 240364 283930
rect 238661 283872 238666 283928
rect 238722 283872 240364 283928
rect 238661 283870 240364 283872
rect 238661 283867 238727 283870
rect 240358 283868 240364 283870
rect 240428 283868 240434 283932
rect 154316 283462 180810 283522
rect 154316 283460 154322 283462
rect 157241 283250 157307 283253
rect 154652 283248 157307 283250
rect 154652 283192 157246 283248
rect 157302 283192 157307 283248
rect 154652 283190 157307 283192
rect 157241 283187 157307 283190
rect 180241 283250 180307 283253
rect 200254 283250 200314 283764
rect 244046 283522 244106 283764
rect 251265 283522 251331 283525
rect 244046 283520 251331 283522
rect 244046 283464 251270 283520
rect 251326 283464 251331 283520
rect 244046 283462 251331 283464
rect 251265 283459 251331 283462
rect 246297 283250 246363 283253
rect 180241 283248 200314 283250
rect 180241 283192 180246 283248
rect 180302 283192 200314 283248
rect 180241 283190 200314 283192
rect 244076 283248 246363 283250
rect 244076 283192 246302 283248
rect 246358 283192 246363 283248
rect 244076 283190 246363 283192
rect 180241 283187 180307 283190
rect 246297 283187 246363 283190
rect 200021 282978 200087 282981
rect 244089 282978 244155 282981
rect 314653 282978 314719 282981
rect 200021 282976 200284 282978
rect 200021 282920 200026 282976
rect 200082 282920 200284 282976
rect 200021 282918 200284 282920
rect 244089 282976 314719 282978
rect 244089 282920 244094 282976
rect 244150 282920 314658 282976
rect 314714 282920 314719 282976
rect 244089 282918 314719 282920
rect 200021 282915 200087 282918
rect 244089 282915 244155 282918
rect 314653 282915 314719 282918
rect 199469 282842 199535 282845
rect 154622 282840 199535 282842
rect 154622 282784 199474 282840
rect 199530 282784 199535 282840
rect 154622 282782 199535 282784
rect 67541 282706 67607 282709
rect 67541 282704 68908 282706
rect 67541 282648 67546 282704
rect 67602 282648 68908 282704
rect 67541 282646 68908 282648
rect 67541 282643 67607 282646
rect 154622 282132 154682 282782
rect 199469 282779 199535 282782
rect 197353 282434 197419 282437
rect 244406 282434 244412 282436
rect 197353 282432 200284 282434
rect 197353 282376 197358 282432
rect 197414 282376 200284 282432
rect 197353 282374 200284 282376
rect 244076 282374 244412 282434
rect 197353 282371 197419 282374
rect 244406 282372 244412 282374
rect 244476 282372 244482 282436
rect 66805 281618 66871 281621
rect 197997 281618 198063 281621
rect 245929 281618 245995 281621
rect 66805 281616 68908 281618
rect 66805 281560 66810 281616
rect 66866 281560 68908 281616
rect 66805 281558 68908 281560
rect 197997 281616 200284 281618
rect 197997 281560 198002 281616
rect 198058 281560 200284 281616
rect 197997 281558 200284 281560
rect 244076 281616 245995 281618
rect 244076 281560 245934 281616
rect 245990 281560 245995 281616
rect 244076 281558 245995 281560
rect 66805 281555 66871 281558
rect 197997 281555 198063 281558
rect 245929 281555 245995 281558
rect 157241 281074 157307 281077
rect 245929 281074 245995 281077
rect 154652 281072 157307 281074
rect 154652 281016 157246 281072
rect 157302 281016 157307 281072
rect 154652 281014 157307 281016
rect 244076 281072 245995 281074
rect 244076 281016 245934 281072
rect 245990 281016 245995 281072
rect 244076 281014 245995 281016
rect 157241 281011 157307 281014
rect 245929 281011 245995 281014
rect 184054 280740 184060 280804
rect 184124 280802 184130 280804
rect 196566 280802 196572 280804
rect 184124 280742 196572 280802
rect 184124 280740 184130 280742
rect 196566 280740 196572 280742
rect 196636 280740 196642 280804
rect 197353 280802 197419 280805
rect 197353 280800 200284 280802
rect 197353 280744 197358 280800
rect 197414 280744 200284 280800
rect 197353 280742 200284 280744
rect 197353 280739 197419 280742
rect 66805 280530 66871 280533
rect 66805 280528 68908 280530
rect 66805 280472 66810 280528
rect 66866 280472 68908 280528
rect 66805 280470 68908 280472
rect 66805 280467 66871 280470
rect 197353 280258 197419 280261
rect 244549 280258 244615 280261
rect 245469 280258 245535 280261
rect 197353 280256 200284 280258
rect -960 279972 480 280212
rect 197353 280200 197358 280256
rect 197414 280200 200284 280256
rect 197353 280198 200284 280200
rect 244076 280256 245535 280258
rect 244076 280200 244554 280256
rect 244610 280200 245474 280256
rect 245530 280200 245535 280256
rect 244076 280198 245535 280200
rect 197353 280195 197419 280198
rect 244549 280195 244615 280198
rect 245469 280195 245535 280198
rect 157241 279986 157307 279989
rect 154652 279984 157307 279986
rect 154652 279928 157246 279984
rect 157302 279928 157307 279984
rect 154652 279926 157307 279928
rect 157241 279923 157307 279926
rect 67173 279442 67239 279445
rect 67950 279442 67956 279444
rect 67173 279440 67956 279442
rect 67173 279384 67178 279440
rect 67234 279384 67956 279440
rect 67173 279382 67956 279384
rect 67173 279379 67239 279382
rect 67950 279380 67956 279382
rect 68020 279442 68026 279444
rect 188429 279442 188495 279445
rect 199326 279442 199332 279444
rect 68020 279382 68908 279442
rect 188429 279440 199332 279442
rect 188429 279384 188434 279440
rect 188490 279384 199332 279440
rect 188429 279382 199332 279384
rect 68020 279380 68026 279382
rect 188429 279379 188495 279382
rect 199326 279380 199332 279382
rect 199396 279380 199402 279444
rect 245929 279442 245995 279445
rect 244076 279440 245995 279442
rect 155309 279306 155375 279309
rect 196893 279306 196959 279309
rect 155309 279304 196959 279306
rect 155309 279248 155314 279304
rect 155370 279248 196898 279304
rect 196954 279248 196959 279304
rect 155309 279246 196959 279248
rect 155309 279243 155375 279246
rect 196893 279243 196959 279246
rect 157241 278898 157307 278901
rect 154652 278896 157307 278898
rect 154652 278840 157246 278896
rect 157302 278840 157307 278896
rect 154652 278838 157307 278840
rect 157241 278835 157307 278838
rect 188981 278898 189047 278901
rect 200254 278898 200314 279412
rect 244076 279384 245934 279440
rect 245990 279384 245995 279440
rect 244076 279382 245995 279384
rect 245929 279379 245995 279382
rect 245653 278898 245719 278901
rect 251265 278900 251331 278901
rect 251214 278898 251220 278900
rect 188981 278896 200314 278898
rect 188981 278840 188986 278896
rect 189042 278840 200314 278896
rect 188981 278838 200314 278840
rect 244076 278896 245719 278898
rect 244076 278840 245658 278896
rect 245714 278840 245719 278896
rect 244076 278838 245719 278840
rect 251174 278838 251220 278898
rect 251284 278896 251331 278900
rect 251326 278840 251331 278896
rect 188981 278835 189047 278838
rect 245653 278835 245719 278838
rect 251214 278836 251220 278838
rect 251284 278836 251331 278840
rect 251265 278835 251331 278836
rect 198089 278762 198155 278765
rect 198641 278762 198707 278765
rect 198089 278760 200130 278762
rect 198089 278704 198094 278760
rect 198150 278704 198646 278760
rect 198702 278704 200130 278760
rect 198089 278702 200130 278704
rect 198089 278699 198155 278702
rect 198641 278699 198707 278702
rect 200070 278626 200130 278702
rect 200070 278566 200284 278626
rect 66437 278354 66503 278357
rect 66437 278352 68908 278354
rect 66437 278296 66442 278352
rect 66498 278296 68908 278352
rect 66437 278294 68908 278296
rect 66437 278291 66503 278294
rect 197353 278082 197419 278085
rect 245929 278082 245995 278085
rect 197353 278080 200284 278082
rect 197353 278024 197358 278080
rect 197414 278024 200284 278080
rect 197353 278022 200284 278024
rect 244076 278080 245995 278082
rect 244076 278024 245934 278080
rect 245990 278024 245995 278080
rect 244076 278022 245995 278024
rect 197353 278019 197419 278022
rect 245929 278019 245995 278022
rect 157241 277810 157307 277813
rect 154652 277808 157307 277810
rect 154652 277752 157246 277808
rect 157302 277752 157307 277808
rect 154652 277750 157307 277752
rect 157241 277747 157307 277750
rect 246021 277538 246087 277541
rect 244076 277536 246087 277538
rect 244076 277480 246026 277536
rect 246082 277480 246087 277536
rect 244076 277478 246087 277480
rect 246021 277475 246087 277478
rect 66805 277266 66871 277269
rect 66805 277264 68908 277266
rect 66805 277208 66810 277264
rect 66866 277208 68908 277264
rect 66805 277206 68908 277208
rect 66805 277203 66871 277206
rect 197854 277204 197860 277268
rect 197924 277266 197930 277268
rect 197924 277206 200284 277266
rect 197924 277204 197930 277206
rect 155309 276722 155375 276725
rect 154652 276720 155375 276722
rect 154652 276664 155314 276720
rect 155370 276664 155375 276720
rect 154652 276662 155375 276664
rect 155309 276659 155375 276662
rect 197353 276722 197419 276725
rect 245745 276722 245811 276725
rect 197353 276720 200284 276722
rect 197353 276664 197358 276720
rect 197414 276664 200284 276720
rect 197353 276662 200284 276664
rect 244076 276720 245811 276722
rect 244076 276664 245750 276720
rect 245806 276664 245811 276720
rect 244076 276662 245811 276664
rect 197353 276659 197419 276662
rect 245745 276659 245811 276662
rect 66161 276178 66227 276181
rect 67950 276178 67956 276180
rect 66161 276176 67956 276178
rect 66161 276120 66166 276176
rect 66222 276120 67956 276176
rect 66161 276118 67956 276120
rect 66161 276115 66227 276118
rect 67950 276116 67956 276118
rect 68020 276178 68026 276180
rect 68020 276118 68908 276178
rect 68020 276116 68026 276118
rect 156873 275906 156939 275909
rect 245929 275906 245995 275909
rect 154652 275904 156939 275906
rect 154652 275848 156878 275904
rect 156934 275848 156939 275904
rect 244076 275904 245995 275906
rect 154652 275846 156939 275848
rect 156873 275843 156939 275846
rect 66805 275362 66871 275365
rect 164877 275362 164943 275365
rect 200254 275362 200314 275876
rect 244076 275848 245934 275904
rect 245990 275848 245995 275904
rect 244076 275846 245995 275848
rect 245929 275843 245995 275846
rect 244222 275634 244228 275636
rect 66805 275360 68908 275362
rect 66805 275304 66810 275360
rect 66866 275304 68908 275360
rect 66805 275302 68908 275304
rect 164877 275360 200314 275362
rect 164877 275304 164882 275360
rect 164938 275304 200314 275360
rect 244046 275574 244228 275634
rect 244046 275332 244106 275574
rect 244222 275572 244228 275574
rect 244292 275572 244298 275636
rect 164877 275302 200314 275304
rect 66805 275299 66871 275302
rect 164877 275299 164943 275302
rect 197353 275090 197419 275093
rect 197353 275088 200284 275090
rect 197353 275032 197358 275088
rect 197414 275032 200284 275088
rect 197353 275030 200284 275032
rect 197353 275027 197419 275030
rect 157241 274818 157307 274821
rect 154652 274816 157307 274818
rect 154652 274760 157246 274816
rect 157302 274760 157307 274816
rect 154652 274758 157307 274760
rect 157241 274755 157307 274758
rect 200021 274546 200087 274549
rect 244273 274546 244339 274549
rect 246481 274546 246547 274549
rect 200021 274544 200284 274546
rect 200021 274488 200026 274544
rect 200082 274488 200284 274544
rect 200021 274486 200284 274488
rect 244076 274544 246547 274546
rect 244076 274488 244278 274544
rect 244334 274488 246486 274544
rect 246542 274488 246547 274544
rect 244076 274486 246547 274488
rect 200021 274483 200087 274486
rect 244273 274483 244339 274486
rect 246481 274483 246547 274486
rect 66805 274274 66871 274277
rect 66805 274272 68908 274274
rect 66805 274216 66810 274272
rect 66866 274216 68908 274272
rect 66805 274214 68908 274216
rect 66805 274211 66871 274214
rect 156505 273730 156571 273733
rect 245653 273730 245719 273733
rect 154652 273728 156571 273730
rect 154652 273672 156510 273728
rect 156566 273672 156571 273728
rect 244076 273728 245719 273730
rect 154652 273670 156571 273672
rect 156505 273667 156571 273670
rect 186313 273458 186379 273461
rect 200254 273458 200314 273700
rect 244076 273672 245658 273728
rect 245714 273672 245719 273728
rect 244076 273670 245719 273672
rect 245653 273667 245719 273670
rect 186313 273456 200314 273458
rect 186313 273400 186318 273456
rect 186374 273400 200314 273456
rect 186313 273398 200314 273400
rect 186313 273395 186379 273398
rect 246246 273322 246252 273324
rect 246070 273262 246252 273322
rect 66805 273186 66871 273189
rect 245837 273186 245903 273189
rect 66805 273184 68908 273186
rect 66805 273128 66810 273184
rect 66866 273128 68908 273184
rect 66805 273126 68908 273128
rect 244076 273184 245903 273186
rect 244076 273128 245842 273184
rect 245898 273128 245903 273184
rect 244076 273126 245903 273128
rect 66805 273123 66871 273126
rect 245837 273123 245903 273126
rect 197353 272914 197419 272917
rect 246070 272914 246130 273262
rect 246246 273260 246252 273262
rect 246316 273322 246322 273324
rect 307753 273322 307819 273325
rect 246316 273320 307819 273322
rect 246316 273264 307758 273320
rect 307814 273264 307819 273320
rect 246316 273262 307819 273264
rect 246316 273260 246322 273262
rect 307753 273259 307819 273262
rect 197353 272912 200284 272914
rect 197353 272856 197358 272912
rect 197414 272856 200284 272912
rect 197353 272854 200284 272856
rect 244046 272854 246130 272914
rect 197353 272851 197419 272854
rect 156965 272642 157031 272645
rect 154652 272640 157031 272642
rect 154652 272584 156970 272640
rect 157026 272584 157031 272640
rect 154652 272582 157031 272584
rect 156965 272579 157031 272582
rect 197445 272370 197511 272373
rect 197445 272368 200284 272370
rect 197445 272312 197450 272368
rect 197506 272312 200284 272368
rect 244046 272340 244106 272854
rect 197445 272310 200284 272312
rect 197445 272307 197511 272310
rect 246113 272234 246179 272237
rect 246389 272234 246455 272237
rect 274582 272234 274588 272236
rect 246113 272232 274588 272234
rect 246113 272176 246118 272232
rect 246174 272176 246394 272232
rect 246450 272176 274588 272232
rect 246113 272174 274588 272176
rect 246113 272171 246179 272174
rect 246389 272171 246455 272174
rect 274582 272172 274588 272174
rect 274652 272172 274658 272236
rect 580349 272234 580415 272237
rect 583520 272234 584960 272324
rect 580349 272232 584960 272234
rect 580349 272176 580354 272232
rect 580410 272176 584960 272232
rect 580349 272174 584960 272176
rect 580349 272171 580415 272174
rect 65885 272098 65951 272101
rect 65885 272096 68908 272098
rect 65885 272040 65890 272096
rect 65946 272040 68908 272096
rect 583520 272084 584960 272174
rect 65885 272038 68908 272040
rect 65885 272035 65951 272038
rect 197445 271554 197511 271557
rect 245837 271554 245903 271557
rect 197445 271552 200284 271554
rect 66805 271010 66871 271013
rect 66805 271008 68908 271010
rect 66805 270952 66810 271008
rect 66866 270952 68908 271008
rect 66805 270950 68908 270952
rect 66805 270947 66871 270950
rect 154622 270874 154682 271524
rect 197445 271496 197450 271552
rect 197506 271496 200284 271552
rect 197445 271494 200284 271496
rect 244076 271552 245903 271554
rect 244076 271496 245842 271552
rect 245898 271496 245903 271552
rect 244076 271494 245903 271496
rect 197445 271491 197511 271494
rect 245837 271491 245903 271494
rect 198549 271010 198615 271013
rect 246113 271010 246179 271013
rect 198549 271008 200284 271010
rect 198549 270952 198554 271008
rect 198610 270952 200284 271008
rect 198549 270950 200284 270952
rect 244076 271008 246179 271010
rect 244076 270952 246118 271008
rect 246174 270952 246179 271008
rect 244076 270950 246179 270952
rect 198549 270947 198615 270950
rect 246113 270947 246179 270950
rect 154622 270814 161490 270874
rect 161430 270602 161490 270814
rect 175917 270602 175983 270605
rect 161430 270600 175983 270602
rect 161430 270544 175922 270600
rect 175978 270544 175983 270600
rect 161430 270542 175983 270544
rect 175917 270539 175983 270542
rect 244222 270540 244228 270604
rect 244292 270602 244298 270604
rect 309225 270602 309291 270605
rect 244292 270600 309291 270602
rect 244292 270544 309230 270600
rect 309286 270544 309291 270600
rect 244292 270542 309291 270544
rect 244292 270540 244298 270542
rect 309225 270539 309291 270542
rect 157241 270466 157307 270469
rect 154652 270464 157307 270466
rect 154652 270408 157246 270464
rect 157302 270408 157307 270464
rect 154652 270406 157307 270408
rect 157241 270403 157307 270406
rect 199377 270194 199443 270197
rect 246297 270194 246363 270197
rect 199377 270192 200284 270194
rect 199377 270136 199382 270192
rect 199438 270136 200284 270192
rect 199377 270134 200284 270136
rect 244076 270192 246363 270194
rect 244076 270136 246302 270192
rect 246358 270136 246363 270192
rect 244076 270134 246363 270136
rect 199377 270131 199443 270134
rect 246297 270131 246363 270134
rect 66805 269922 66871 269925
rect 66805 269920 68908 269922
rect 66805 269864 66810 269920
rect 66866 269864 68908 269920
rect 66805 269862 68908 269864
rect 66805 269859 66871 269862
rect 245929 269650 245995 269653
rect 244076 269648 245995 269650
rect 244076 269592 245934 269648
rect 245990 269592 245995 269648
rect 244076 269590 245995 269592
rect 245929 269587 245995 269590
rect 161974 269378 161980 269380
rect 154652 269318 161980 269378
rect 161974 269316 161980 269318
rect 162044 269316 162050 269380
rect 197353 269378 197419 269381
rect 197353 269376 200284 269378
rect 197353 269320 197358 269376
rect 197414 269320 200284 269376
rect 197353 269318 200284 269320
rect 197353 269315 197419 269318
rect 244038 269044 244044 269108
rect 244108 269044 244114 269108
rect 67633 268834 67699 268837
rect 197353 268834 197419 268837
rect 67633 268832 68908 268834
rect 67633 268776 67638 268832
rect 67694 268776 68908 268832
rect 67633 268774 68908 268776
rect 197353 268832 200284 268834
rect 197353 268776 197358 268832
rect 197414 268776 200284 268832
rect 244046 268804 244106 269044
rect 197353 268774 200284 268776
rect 67633 268771 67699 268774
rect 197353 268771 197419 268774
rect 156413 268290 156479 268293
rect 154652 268288 156479 268290
rect 154652 268232 156418 268288
rect 156474 268232 156479 268288
rect 154652 268230 156479 268232
rect 156413 268227 156479 268230
rect 197353 268018 197419 268021
rect 245745 268018 245811 268021
rect 197353 268016 200284 268018
rect 197353 267960 197358 268016
rect 197414 267960 200284 268016
rect 197353 267958 200284 267960
rect 244076 268016 245811 268018
rect 244076 267960 245750 268016
rect 245806 267960 245811 268016
rect 244076 267958 245811 267960
rect 197353 267955 197419 267958
rect 245745 267955 245811 267958
rect 66621 267746 66687 267749
rect 66621 267744 68908 267746
rect 66621 267688 66626 267744
rect 66682 267688 68908 267744
rect 66621 267686 68908 267688
rect 66621 267683 66687 267686
rect 156321 267474 156387 267477
rect 245929 267474 245995 267477
rect 154652 267472 156387 267474
rect 154652 267416 156326 267472
rect 156382 267416 156387 267472
rect 154652 267414 156387 267416
rect 244076 267472 245995 267474
rect 244076 267416 245934 267472
rect 245990 267416 245995 267472
rect 244076 267414 245995 267416
rect 156321 267411 156387 267414
rect 245929 267411 245995 267414
rect -960 267202 480 267292
rect 3417 267202 3483 267205
rect -960 267200 3483 267202
rect -960 267144 3422 267200
rect 3478 267144 3483 267200
rect -960 267142 3483 267144
rect -960 267052 480 267142
rect 3417 267139 3483 267142
rect 197353 267202 197419 267205
rect 197353 267200 200284 267202
rect 197353 267144 197358 267200
rect 197414 267144 200284 267200
rect 197353 267142 200284 267144
rect 197353 267139 197419 267142
rect 159449 267066 159515 267069
rect 198181 267066 198247 267069
rect 159449 267064 198247 267066
rect 159449 267008 159454 267064
rect 159510 267008 198186 267064
rect 198242 267008 198247 267064
rect 159449 267006 198247 267008
rect 159449 267003 159515 267006
rect 198181 267003 198247 267006
rect 67398 266868 67404 266932
rect 67468 266930 67474 266932
rect 67468 266870 68908 266930
rect 67468 266868 67474 266870
rect 197445 266658 197511 266661
rect 197445 266656 200284 266658
rect 197445 266600 197450 266656
rect 197506 266600 200284 266656
rect 197445 266598 200284 266600
rect 244076 266598 248430 266658
rect 197445 266595 197511 266598
rect 248370 266522 248430 266598
rect 263685 266522 263751 266525
rect 248370 266520 263751 266522
rect 248370 266464 263690 266520
rect 263746 266464 263751 266520
rect 248370 266462 263751 266464
rect 263685 266459 263751 266462
rect 157241 266386 157307 266389
rect 154652 266384 157307 266386
rect 154652 266328 157246 266384
rect 157302 266328 157307 266384
rect 154652 266326 157307 266328
rect 157241 266323 157307 266326
rect 66805 265842 66871 265845
rect 196617 265842 196683 265845
rect 245929 265842 245995 265845
rect 66805 265840 68908 265842
rect 66805 265784 66810 265840
rect 66866 265784 68908 265840
rect 66805 265782 68908 265784
rect 196617 265840 200284 265842
rect 196617 265784 196622 265840
rect 196678 265784 200284 265840
rect 196617 265782 200284 265784
rect 244076 265840 245995 265842
rect 244076 265784 245934 265840
rect 245990 265784 245995 265840
rect 244076 265782 245995 265784
rect 66805 265779 66871 265782
rect 196617 265779 196683 265782
rect 245929 265779 245995 265782
rect 166206 265508 166212 265572
rect 166276 265570 166282 265572
rect 198774 265570 198780 265572
rect 166276 265510 198780 265570
rect 166276 265508 166282 265510
rect 198774 265508 198780 265510
rect 198844 265508 198850 265572
rect 157241 265298 157307 265301
rect 154652 265296 157307 265298
rect 154652 265240 157246 265296
rect 157302 265240 157307 265296
rect 154652 265238 157307 265240
rect 157241 265235 157307 265238
rect 197353 265298 197419 265301
rect 245745 265298 245811 265301
rect 197353 265296 200284 265298
rect 197353 265240 197358 265296
rect 197414 265240 200284 265296
rect 197353 265238 200284 265240
rect 244076 265296 245811 265298
rect 244076 265240 245750 265296
rect 245806 265240 245811 265296
rect 244076 265238 245811 265240
rect 197353 265235 197419 265238
rect 245745 265235 245811 265238
rect 66713 264754 66779 264757
rect 66713 264752 68908 264754
rect 66713 264696 66718 264752
rect 66774 264696 68908 264752
rect 66713 264694 68908 264696
rect 66713 264691 66779 264694
rect 197445 264482 197511 264485
rect 244549 264482 244615 264485
rect 197445 264480 200284 264482
rect 197445 264424 197450 264480
rect 197506 264424 200284 264480
rect 197445 264422 200284 264424
rect 244076 264480 244615 264482
rect 244076 264424 244554 264480
rect 244610 264424 244615 264480
rect 244076 264422 244615 264424
rect 197445 264419 197511 264422
rect 244549 264419 244615 264422
rect 155217 264210 155283 264213
rect 154652 264208 155283 264210
rect 154652 264152 155222 264208
rect 155278 264152 155283 264208
rect 154652 264150 155283 264152
rect 155217 264147 155283 264150
rect 155350 264148 155356 264212
rect 155420 264210 155426 264212
rect 174629 264210 174695 264213
rect 155420 264208 174695 264210
rect 155420 264152 174634 264208
rect 174690 264152 174695 264208
rect 155420 264150 174695 264152
rect 155420 264148 155426 264150
rect 174629 264147 174695 264150
rect 245837 263938 245903 263941
rect 244076 263936 245903 263938
rect 244076 263880 245842 263936
rect 245898 263880 245903 263936
rect 244076 263878 245903 263880
rect 245837 263875 245903 263878
rect 66805 263666 66871 263669
rect 197353 263666 197419 263669
rect 66805 263664 68908 263666
rect 66805 263608 66810 263664
rect 66866 263608 68908 263664
rect 66805 263606 68908 263608
rect 197353 263664 200284 263666
rect 197353 263608 197358 263664
rect 197414 263608 200284 263664
rect 197353 263606 200284 263608
rect 66805 263603 66871 263606
rect 197353 263603 197419 263606
rect 156413 263122 156479 263125
rect 245653 263122 245719 263125
rect 154652 263120 156479 263122
rect 154652 263064 156418 263120
rect 156474 263064 156479 263120
rect 244076 263120 245719 263122
rect 154652 263062 156479 263064
rect 156413 263059 156479 263062
rect 66805 262578 66871 262581
rect 174629 262578 174695 262581
rect 200254 262578 200314 263092
rect 244076 263064 245658 263120
rect 245714 263064 245719 263120
rect 244076 263062 245719 263064
rect 245653 263059 245719 263062
rect 66805 262576 68908 262578
rect 66805 262520 66810 262576
rect 66866 262520 68908 262576
rect 66805 262518 68908 262520
rect 174629 262576 200314 262578
rect 174629 262520 174634 262576
rect 174690 262520 200314 262576
rect 174629 262518 200314 262520
rect 66805 262515 66871 262518
rect 174629 262515 174695 262518
rect 196617 262306 196683 262309
rect 247125 262306 247191 262309
rect 196617 262304 200284 262306
rect 196617 262248 196622 262304
rect 196678 262248 200284 262304
rect 196617 262246 200284 262248
rect 244076 262304 247191 262306
rect 244076 262248 247130 262304
rect 247186 262248 247191 262304
rect 244076 262246 247191 262248
rect 196617 262243 196683 262246
rect 247125 262243 247191 262246
rect 156965 262034 157031 262037
rect 154652 262032 157031 262034
rect 154652 261976 156970 262032
rect 157026 261976 157031 262032
rect 154652 261974 157031 261976
rect 156965 261971 157031 261974
rect 66805 261490 66871 261493
rect 197353 261490 197419 261493
rect 66805 261488 68908 261490
rect 66805 261432 66810 261488
rect 66866 261432 68908 261488
rect 66805 261430 68908 261432
rect 197353 261488 200284 261490
rect 197353 261432 197358 261488
rect 197414 261432 200284 261488
rect 197353 261430 200284 261432
rect 66805 261427 66871 261430
rect 197353 261427 197419 261430
rect 244046 261218 244106 261732
rect 256785 261218 256851 261221
rect 244046 261216 256851 261218
rect 244046 261160 256790 261216
rect 256846 261160 256851 261216
rect 244046 261158 256851 261160
rect 256785 261155 256851 261158
rect 157241 260946 157307 260949
rect 154652 260944 157307 260946
rect 154652 260888 157246 260944
rect 157302 260888 157307 260944
rect 154652 260886 157307 260888
rect 157241 260883 157307 260886
rect 197997 260946 198063 260949
rect 246389 260946 246455 260949
rect 197997 260944 200284 260946
rect 197997 260888 198002 260944
rect 198058 260888 200284 260944
rect 197997 260886 200284 260888
rect 244076 260944 246455 260946
rect 244076 260888 246394 260944
rect 246450 260888 246455 260944
rect 244076 260886 246455 260888
rect 197997 260883 198063 260886
rect 246389 260883 246455 260886
rect 67817 260402 67883 260405
rect 67817 260400 68908 260402
rect 67817 260344 67822 260400
rect 67878 260344 68908 260400
rect 67817 260342 68908 260344
rect 67817 260339 67883 260342
rect 197353 260130 197419 260133
rect 245745 260130 245811 260133
rect 197353 260128 200284 260130
rect 197353 260072 197358 260128
rect 197414 260072 200284 260128
rect 197353 260070 200284 260072
rect 244076 260128 245811 260130
rect 244076 260072 245750 260128
rect 245806 260072 245811 260128
rect 244076 260070 245811 260072
rect 197353 260067 197419 260070
rect 245745 260067 245811 260070
rect 156689 259858 156755 259861
rect 154652 259856 156755 259858
rect 154652 259800 156694 259856
rect 156750 259800 156755 259856
rect 154652 259798 156755 259800
rect 156689 259795 156755 259798
rect 244457 259586 244523 259589
rect 244076 259584 244523 259586
rect 244076 259528 244462 259584
rect 244518 259528 244523 259584
rect 244076 259526 244523 259528
rect 244457 259523 244523 259526
rect 198549 259450 198615 259453
rect 198774 259450 198780 259452
rect 198549 259448 198780 259450
rect 198549 259392 198554 259448
rect 198610 259392 198780 259448
rect 198549 259390 198780 259392
rect 198549 259387 198615 259390
rect 198774 259388 198780 259390
rect 198844 259388 198850 259452
rect 197353 259314 197419 259317
rect 243997 259314 244063 259317
rect 197353 259312 200284 259314
rect 69430 258772 69490 259284
rect 197353 259256 197358 259312
rect 197414 259256 200284 259312
rect 197353 259254 200284 259256
rect 243997 259312 244106 259314
rect 243997 259256 244002 259312
rect 244058 259256 244106 259312
rect 197353 259251 197419 259254
rect 243997 259251 244106 259256
rect 69422 258708 69428 258772
rect 69492 258708 69498 258772
rect 66253 258090 66319 258093
rect 66253 258088 66362 258090
rect 66253 258032 66258 258088
rect 66314 258032 66362 258088
rect 66253 258027 66362 258032
rect 66302 257954 66362 258027
rect 68878 257954 68938 258468
rect 154622 258362 154682 259012
rect 197445 258770 197511 258773
rect 244046 258770 244106 259251
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 245837 258770 245903 258773
rect 197445 258768 200284 258770
rect 197445 258712 197450 258768
rect 197506 258712 200284 258768
rect 244046 258768 245903 258770
rect 244046 258740 245842 258768
rect 197445 258710 200284 258712
rect 244076 258712 245842 258740
rect 245898 258712 245903 258768
rect 583520 258756 584960 258846
rect 244076 258710 245903 258712
rect 197445 258707 197511 258710
rect 245837 258707 245903 258710
rect 154622 258302 164250 258362
rect 156873 257954 156939 257957
rect 66302 257894 68938 257954
rect 154652 257952 156939 257954
rect 154652 257896 156878 257952
rect 156934 257896 156939 257952
rect 154652 257894 156939 257896
rect 164190 257954 164250 258302
rect 245929 258226 245995 258229
rect 244076 258224 245995 258226
rect 244076 258168 245934 258224
rect 245990 258168 245995 258224
rect 244076 258166 245995 258168
rect 245929 258163 245995 258166
rect 168966 258028 168972 258092
rect 169036 258028 169042 258092
rect 168974 257954 169034 258028
rect 164190 257894 169034 257954
rect 197445 257954 197511 257957
rect 197445 257952 200284 257954
rect 197445 257896 197450 257952
rect 197506 257896 200284 257952
rect 197445 257894 200284 257896
rect 156873 257891 156939 257894
rect 197445 257891 197511 257894
rect 65977 257410 66043 257413
rect 245653 257410 245719 257413
rect 65977 257408 68908 257410
rect 65977 257352 65982 257408
rect 66038 257352 68908 257408
rect 65977 257350 68908 257352
rect 200070 257350 200284 257410
rect 244076 257408 245719 257410
rect 244076 257352 245658 257408
rect 245714 257352 245719 257408
rect 244076 257350 245719 257352
rect 65977 257347 66043 257350
rect 161013 257274 161079 257277
rect 180057 257274 180123 257277
rect 161013 257272 180123 257274
rect 161013 257216 161018 257272
rect 161074 257216 180062 257272
rect 180118 257216 180123 257272
rect 161013 257214 180123 257216
rect 161013 257211 161079 257214
rect 180057 257211 180123 257214
rect 183461 257274 183527 257277
rect 200070 257274 200130 257350
rect 245653 257347 245719 257350
rect 183461 257272 200130 257274
rect 183461 257216 183466 257272
rect 183522 257216 200130 257272
rect 183461 257214 200130 257216
rect 183461 257211 183527 257214
rect 157241 256866 157307 256869
rect 154652 256864 157307 256866
rect 154652 256808 157246 256864
rect 157302 256808 157307 256864
rect 154652 256806 157307 256808
rect 157241 256803 157307 256806
rect 182173 256730 182239 256733
rect 183461 256730 183527 256733
rect 182173 256728 183527 256730
rect 182173 256672 182178 256728
rect 182234 256672 183466 256728
rect 183522 256672 183527 256728
rect 182173 256670 183527 256672
rect 182173 256667 182239 256670
rect 183461 256667 183527 256670
rect 199561 256594 199627 256597
rect 245929 256594 245995 256597
rect 199561 256592 200284 256594
rect 199561 256536 199566 256592
rect 199622 256536 200284 256592
rect 199561 256534 200284 256536
rect 244076 256592 245995 256594
rect 244076 256536 245934 256592
rect 245990 256536 245995 256592
rect 244076 256534 245995 256536
rect 199561 256531 199627 256534
rect 245929 256531 245995 256534
rect 66805 256322 66871 256325
rect 66805 256320 68908 256322
rect 66805 256264 66810 256320
rect 66866 256264 68908 256320
rect 66805 256262 68908 256264
rect 66805 256259 66871 256262
rect 247217 256050 247283 256053
rect 244076 256048 247283 256050
rect 244076 255992 247222 256048
rect 247278 255992 247283 256048
rect 244076 255990 247283 255992
rect 247217 255987 247283 255990
rect 160829 255914 160895 255917
rect 189901 255914 189967 255917
rect 160829 255912 189967 255914
rect 160829 255856 160834 255912
rect 160890 255856 189906 255912
rect 189962 255856 189967 255912
rect 160829 255854 189967 255856
rect 160829 255851 160895 255854
rect 189901 255851 189967 255854
rect 156505 255778 156571 255781
rect 154652 255776 156571 255778
rect 154652 255720 156510 255776
rect 156566 255720 156571 255776
rect 154652 255718 156571 255720
rect 156505 255715 156571 255718
rect 197353 255778 197419 255781
rect 197353 255776 200284 255778
rect 197353 255720 197358 255776
rect 197414 255720 200284 255776
rect 197353 255718 200284 255720
rect 197353 255715 197419 255718
rect 67449 255234 67515 255237
rect 197353 255234 197419 255237
rect 245929 255234 245995 255237
rect 67449 255232 68908 255234
rect 67449 255176 67454 255232
rect 67510 255176 68908 255232
rect 67449 255174 68908 255176
rect 197353 255232 200284 255234
rect 197353 255176 197358 255232
rect 197414 255176 200284 255232
rect 197353 255174 200284 255176
rect 244076 255232 245995 255234
rect 244076 255176 245934 255232
rect 245990 255176 245995 255232
rect 244076 255174 245995 255176
rect 67449 255171 67515 255174
rect 197353 255171 197419 255174
rect 245929 255171 245995 255174
rect 157241 254690 157307 254693
rect 154652 254688 157307 254690
rect 154652 254632 157246 254688
rect 157302 254632 157307 254688
rect 154652 254630 157307 254632
rect 157241 254627 157307 254630
rect 162669 254554 162735 254557
rect 178677 254554 178743 254557
rect 162669 254552 178743 254554
rect 162669 254496 162674 254552
rect 162730 254496 178682 254552
rect 178738 254496 178743 254552
rect 162669 254494 178743 254496
rect 162669 254491 162735 254494
rect 178677 254491 178743 254494
rect 193806 254356 193812 254420
rect 193876 254418 193882 254420
rect 245837 254418 245903 254421
rect 193876 254358 200284 254418
rect 244076 254416 245903 254418
rect 244076 254360 245842 254416
rect 245898 254360 245903 254416
rect 244076 254358 245903 254360
rect 193876 254356 193882 254358
rect 245837 254355 245903 254358
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 66805 254146 66871 254149
rect 66805 254144 68908 254146
rect 66805 254088 66810 254144
rect 66866 254088 68908 254144
rect 66805 254086 68908 254088
rect 66805 254083 66871 254086
rect 245929 253874 245995 253877
rect 244076 253872 245995 253874
rect 244076 253816 245934 253872
rect 245990 253816 245995 253872
rect 244076 253814 245995 253816
rect 245929 253811 245995 253814
rect 157241 253602 157307 253605
rect 154652 253600 157307 253602
rect 154652 253544 157246 253600
rect 157302 253544 157307 253600
rect 154652 253542 157307 253544
rect 157241 253539 157307 253542
rect 197445 253602 197511 253605
rect 197445 253600 200284 253602
rect 197445 253544 197450 253600
rect 197506 253544 200284 253600
rect 197445 253542 200284 253544
rect 197445 253539 197511 253542
rect 167637 253194 167703 253197
rect 191189 253194 191255 253197
rect 167637 253192 191255 253194
rect 167637 253136 167642 253192
rect 167698 253136 191194 253192
rect 191250 253136 191255 253192
rect 167637 253134 191255 253136
rect 167637 253131 167703 253134
rect 191189 253131 191255 253134
rect 66805 253058 66871 253061
rect 197353 253058 197419 253061
rect 244365 253058 244431 253061
rect 245653 253058 245719 253061
rect 66805 253056 68908 253058
rect 66805 253000 66810 253056
rect 66866 253000 68908 253056
rect 66805 252998 68908 253000
rect 197353 253056 200284 253058
rect 197353 253000 197358 253056
rect 197414 253000 200284 253056
rect 197353 252998 200284 253000
rect 244076 253056 245719 253058
rect 244076 253000 244370 253056
rect 244426 253000 245658 253056
rect 245714 253000 245719 253056
rect 244076 252998 245719 253000
rect 66805 252995 66871 252998
rect 197353 252995 197419 252998
rect 244365 252995 244431 252998
rect 245653 252995 245719 252998
rect 157149 252514 157215 252517
rect 154652 252512 157215 252514
rect 154652 252456 157154 252512
rect 157210 252456 157215 252512
rect 154652 252454 157215 252456
rect 157149 252451 157215 252454
rect 197997 252242 198063 252245
rect 245929 252242 245995 252245
rect 197997 252240 200284 252242
rect 197997 252184 198002 252240
rect 198058 252184 200284 252240
rect 197997 252182 200284 252184
rect 244076 252240 245995 252242
rect 244076 252184 245934 252240
rect 245990 252184 245995 252240
rect 244076 252182 245995 252184
rect 197997 252179 198063 252182
rect 245929 252179 245995 252182
rect 66662 251908 66668 251972
rect 66732 251970 66738 251972
rect 66732 251910 68908 251970
rect 66732 251908 66738 251910
rect 197353 251698 197419 251701
rect 245837 251698 245903 251701
rect 197353 251696 200284 251698
rect 197353 251640 197358 251696
rect 197414 251640 200284 251696
rect 197353 251638 200284 251640
rect 244076 251696 245903 251698
rect 244076 251640 245842 251696
rect 245898 251640 245903 251696
rect 244076 251638 245903 251640
rect 197353 251635 197419 251638
rect 245837 251635 245903 251638
rect 157241 251426 157307 251429
rect 154652 251424 157307 251426
rect 154652 251368 157246 251424
rect 157302 251368 157307 251424
rect 154652 251366 157307 251368
rect 157241 251363 157307 251366
rect 67725 250882 67791 250885
rect 197353 250882 197419 250885
rect 67725 250880 68908 250882
rect 67725 250824 67730 250880
rect 67786 250824 68908 250880
rect 67725 250822 68908 250824
rect 197353 250880 200284 250882
rect 197353 250824 197358 250880
rect 197414 250824 200284 250880
rect 197353 250822 200284 250824
rect 67725 250819 67791 250822
rect 197353 250819 197419 250822
rect 157241 250610 157307 250613
rect 244046 250612 244106 250852
rect 154652 250608 157307 250610
rect 154652 250552 157246 250608
rect 157302 250552 157307 250608
rect 154652 250550 157307 250552
rect 157241 250547 157307 250550
rect 244038 250548 244044 250612
rect 244108 250548 244114 250612
rect 245101 250338 245167 250341
rect 244076 250336 245167 250338
rect 244076 250280 245106 250336
rect 245162 250280 245167 250336
rect 244076 250278 245167 250280
rect 245101 250275 245167 250278
rect 66437 250066 66503 250069
rect 66437 250064 68908 250066
rect 66437 250008 66442 250064
rect 66498 250008 68908 250064
rect 66437 250006 68908 250008
rect 200070 250006 200284 250066
rect 66437 250003 66503 250006
rect 178953 249930 179019 249933
rect 200070 249930 200130 250006
rect 178953 249928 200130 249930
rect 178953 249872 178958 249928
rect 179014 249872 200130 249928
rect 178953 249870 200130 249872
rect 178953 249867 179019 249870
rect 156505 249522 156571 249525
rect 154652 249520 156571 249522
rect 154652 249464 156510 249520
rect 156566 249464 156571 249520
rect 154652 249462 156571 249464
rect 156505 249459 156571 249462
rect 197353 249522 197419 249525
rect 245929 249522 245995 249525
rect 197353 249520 200284 249522
rect 197353 249464 197358 249520
rect 197414 249464 200284 249520
rect 197353 249462 200284 249464
rect 244076 249520 245995 249522
rect 244076 249464 245934 249520
rect 245990 249464 245995 249520
rect 244076 249462 245995 249464
rect 197353 249459 197419 249462
rect 245929 249459 245995 249462
rect 67766 248916 67772 248980
rect 67836 248978 67842 248980
rect 67836 248918 68908 248978
rect 67836 248916 67842 248918
rect 197353 248706 197419 248709
rect 197353 248704 200284 248706
rect 197353 248648 197358 248704
rect 197414 248648 200284 248704
rect 197353 248646 200284 248648
rect 197353 248643 197419 248646
rect 244046 248437 244106 248676
rect 156965 248434 157031 248437
rect 154652 248432 157031 248434
rect 154652 248376 156970 248432
rect 157026 248376 157031 248432
rect 154652 248374 157031 248376
rect 156965 248371 157031 248374
rect 243997 248432 244106 248437
rect 243997 248376 244002 248432
rect 244058 248376 244106 248432
rect 243997 248374 244106 248376
rect 243997 248371 244063 248374
rect 245929 248162 245995 248165
rect 244076 248160 245995 248162
rect 244076 248104 245934 248160
rect 245990 248104 245995 248160
rect 244076 248102 245995 248104
rect 245929 248099 245995 248102
rect 66805 247890 66871 247893
rect 197353 247890 197419 247893
rect 66805 247888 68908 247890
rect 66805 247832 66810 247888
rect 66866 247832 68908 247888
rect 66805 247830 68908 247832
rect 197353 247888 200284 247890
rect 197353 247832 197358 247888
rect 197414 247832 200284 247888
rect 197353 247830 200284 247832
rect 66805 247827 66871 247830
rect 197353 247827 197419 247830
rect 156781 247346 156847 247349
rect 154652 247344 156847 247346
rect 154652 247288 156786 247344
rect 156842 247288 156847 247344
rect 154652 247286 156847 247288
rect 156781 247283 156847 247286
rect 187049 247346 187115 247349
rect 245694 247346 245700 247348
rect 187049 247344 200284 247346
rect 187049 247288 187054 247344
rect 187110 247288 200284 247344
rect 187049 247286 200284 247288
rect 244076 247286 245700 247346
rect 187049 247283 187115 247286
rect 245694 247284 245700 247286
rect 245764 247284 245770 247348
rect 158713 247210 158779 247213
rect 158713 247208 180810 247210
rect 158713 247152 158718 247208
rect 158774 247152 180810 247208
rect 158713 247150 180810 247152
rect 158713 247147 158779 247150
rect 180750 247074 180810 247150
rect 198774 247074 198780 247076
rect 180750 247014 198780 247074
rect 198774 247012 198780 247014
rect 198844 247074 198850 247076
rect 199878 247074 199884 247076
rect 198844 247014 199884 247074
rect 198844 247012 198850 247014
rect 199878 247012 199884 247014
rect 199948 247012 199954 247076
rect 67265 246802 67331 246805
rect 67265 246800 68908 246802
rect 67265 246744 67270 246800
rect 67326 246744 68908 246800
rect 67265 246742 68908 246744
rect 67265 246739 67331 246742
rect 197353 246530 197419 246533
rect 245837 246530 245903 246533
rect 197353 246528 200284 246530
rect 197353 246472 197358 246528
rect 197414 246472 200284 246528
rect 197353 246470 200284 246472
rect 244076 246528 245903 246530
rect 244076 246472 245842 246528
rect 245898 246472 245903 246528
rect 244076 246470 245903 246472
rect 197353 246467 197419 246470
rect 245837 246467 245903 246470
rect 157241 246258 157307 246261
rect 196617 246258 196683 246261
rect 154652 246256 157307 246258
rect 154652 246200 157246 246256
rect 157302 246200 157307 246256
rect 154652 246198 157307 246200
rect 157241 246195 157307 246198
rect 161430 246256 196683 246258
rect 161430 246200 196622 246256
rect 196678 246200 196683 246256
rect 161430 246198 196683 246200
rect 156781 246122 156847 246125
rect 161430 246122 161490 246198
rect 196617 246195 196683 246198
rect 156781 246120 161490 246122
rect 156781 246064 156786 246120
rect 156842 246064 161490 246120
rect 156781 246062 161490 246064
rect 156781 246059 156847 246062
rect 195462 245924 195468 245988
rect 195532 245986 195538 245988
rect 246389 245986 246455 245989
rect 195532 245926 200284 245986
rect 244076 245984 246455 245986
rect 244076 245928 246394 245984
rect 246450 245928 246455 245984
rect 244076 245926 246455 245928
rect 195532 245924 195538 245926
rect 246389 245923 246455 245926
rect 67633 245714 67699 245717
rect 67633 245712 68908 245714
rect 67633 245656 67638 245712
rect 67694 245656 68908 245712
rect 67633 245654 68908 245656
rect 67633 245651 67699 245654
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 160737 245170 160803 245173
rect 154652 245168 160803 245170
rect 154652 245112 160742 245168
rect 160798 245112 160803 245168
rect 154652 245110 160803 245112
rect 160737 245107 160803 245110
rect 197077 245170 197143 245173
rect 244365 245170 244431 245173
rect 197077 245168 200284 245170
rect 197077 245112 197082 245168
rect 197138 245112 200284 245168
rect 197077 245110 200284 245112
rect 244076 245168 244431 245170
rect 244076 245112 244370 245168
rect 244426 245112 244431 245168
rect 244076 245110 244431 245112
rect 197077 245107 197143 245110
rect 244365 245107 244431 245110
rect 66621 244626 66687 244629
rect 245929 244626 245995 244629
rect 66621 244624 68908 244626
rect 66621 244568 66626 244624
rect 66682 244568 68908 244624
rect 66621 244566 68908 244568
rect 244076 244624 245995 244626
rect 244076 244568 245934 244624
rect 245990 244568 245995 244624
rect 244076 244566 245995 244568
rect 66621 244563 66687 244566
rect 245929 244563 245995 244566
rect 197445 244354 197511 244357
rect 197445 244352 200284 244354
rect 197445 244296 197450 244352
rect 197506 244296 200284 244352
rect 197445 244294 200284 244296
rect 197445 244291 197511 244294
rect 156045 244082 156111 244085
rect 154652 244080 156111 244082
rect 154652 244024 156050 244080
rect 156106 244024 156111 244080
rect 154652 244022 156111 244024
rect 156045 244019 156111 244022
rect 154430 243884 154436 243948
rect 154500 243946 154506 243948
rect 174721 243946 174787 243949
rect 154500 243944 174787 243946
rect 154500 243888 174726 243944
rect 174782 243888 174787 243944
rect 154500 243886 174787 243888
rect 154500 243884 154506 243886
rect 174721 243883 174787 243886
rect 195278 243748 195284 243812
rect 195348 243810 195354 243812
rect 244641 243810 244707 243813
rect 195348 243750 200284 243810
rect 244076 243808 244707 243810
rect 244076 243752 244646 243808
rect 244702 243752 244707 243808
rect 244076 243750 244707 243752
rect 195348 243748 195354 243750
rect 244641 243747 244707 243750
rect 66805 243538 66871 243541
rect 66805 243536 68908 243538
rect 66805 243480 66810 243536
rect 66866 243480 68908 243536
rect 66805 243478 68908 243480
rect 66805 243475 66871 243478
rect 65885 243402 65951 243405
rect 69422 243402 69428 243404
rect 65885 243400 69428 243402
rect 65885 243344 65890 243400
rect 65946 243344 69428 243400
rect 65885 243342 69428 243344
rect 65885 243339 65951 243342
rect 69422 243340 69428 243342
rect 69492 243340 69498 243404
rect 154798 243204 154804 243268
rect 154868 243266 154874 243268
rect 154941 243266 155007 243269
rect 154868 243264 155007 243266
rect 154868 243208 154946 243264
rect 155002 243208 155007 243264
rect 154868 243206 155007 243208
rect 154868 243204 154874 243206
rect 154941 243203 155007 243206
rect 155401 242994 155467 242997
rect 154652 242992 155467 242994
rect 154652 242936 155406 242992
rect 155462 242936 155467 242992
rect 154652 242934 155467 242936
rect 155401 242931 155467 242934
rect 197353 242994 197419 242997
rect 248454 242994 248460 242996
rect 197353 242992 200284 242994
rect 197353 242936 197358 242992
rect 197414 242936 200284 242992
rect 197353 242934 200284 242936
rect 244076 242934 248460 242994
rect 197353 242931 197419 242934
rect 248454 242932 248460 242934
rect 248524 242932 248530 242996
rect 67081 242858 67147 242861
rect 67398 242858 67404 242860
rect 67081 242856 67404 242858
rect 67081 242800 67086 242856
rect 67142 242800 67404 242856
rect 67081 242798 67404 242800
rect 67081 242795 67147 242798
rect 67398 242796 67404 242798
rect 67468 242796 67474 242860
rect 191649 242586 191715 242589
rect 197997 242586 198063 242589
rect 191649 242584 198063 242586
rect 191649 242528 191654 242584
rect 191710 242528 198002 242584
rect 198058 242528 198063 242584
rect 191649 242526 198063 242528
rect 191649 242523 191715 242526
rect 197997 242523 198063 242526
rect 245929 242450 245995 242453
rect 244076 242448 245995 242450
rect 69430 241906 69490 242420
rect 244076 242392 245934 242448
rect 245990 242392 245995 242448
rect 244076 242390 245995 242392
rect 245929 242387 245995 242390
rect 156229 242178 156295 242181
rect 154652 242176 156295 242178
rect 154652 242120 156234 242176
rect 156290 242120 156295 242176
rect 154652 242118 156295 242120
rect 156229 242115 156295 242118
rect 197537 242178 197603 242181
rect 197537 242176 200284 242178
rect 197537 242120 197542 242176
rect 197598 242120 200284 242176
rect 197537 242118 200284 242120
rect 197537 242115 197603 242118
rect 135989 242044 136055 242045
rect 135989 242042 136036 242044
rect 135944 242040 136036 242042
rect 135944 241984 135994 242040
rect 135944 241982 136036 241984
rect 135989 241980 136036 241982
rect 136100 241980 136106 242044
rect 138054 241980 138060 242044
rect 138124 242042 138130 242044
rect 138197 242042 138263 242045
rect 138124 242040 138263 242042
rect 138124 241984 138202 242040
rect 138258 241984 138263 242040
rect 138124 241982 138263 241984
rect 138124 241980 138130 241982
rect 135989 241979 136055 241980
rect 138197 241979 138263 241982
rect 146753 242042 146819 242045
rect 147438 242042 147444 242044
rect 146753 242040 147444 242042
rect 146753 241984 146758 242040
rect 146814 241984 147444 242040
rect 146753 241982 147444 241984
rect 146753 241979 146819 241982
rect 147438 241980 147444 241982
rect 147508 241980 147514 242044
rect 151854 241980 151860 242044
rect 151924 242042 151930 242044
rect 152549 242042 152615 242045
rect 151924 242040 152615 242042
rect 151924 241984 152554 242040
rect 152610 241984 152615 242040
rect 151924 241982 152615 241984
rect 151924 241980 151930 241982
rect 152549 241979 152615 241982
rect 70301 241906 70367 241909
rect 69430 241904 70367 241906
rect 69430 241848 70306 241904
rect 70362 241848 70367 241904
rect 69430 241846 70367 241848
rect 70301 241843 70367 241846
rect 67449 241770 67515 241773
rect 69657 241770 69723 241773
rect 67449 241768 69723 241770
rect 67449 241712 67454 241768
rect 67510 241712 69662 241768
rect 69718 241712 69723 241768
rect 67449 241710 69723 241712
rect 67449 241707 67515 241710
rect 69657 241707 69723 241710
rect 154021 241634 154087 241637
rect 158713 241634 158779 241637
rect 191649 241636 191715 241637
rect 191598 241634 191604 241636
rect 154021 241632 158779 241634
rect 154021 241576 154026 241632
rect 154082 241576 158718 241632
rect 158774 241576 158779 241632
rect 154021 241574 158779 241576
rect 191558 241574 191604 241634
rect 191668 241632 191715 241636
rect 191710 241576 191715 241632
rect 154021 241571 154087 241574
rect 158713 241571 158779 241574
rect 191598 241572 191604 241574
rect 191668 241572 191715 241576
rect 191649 241571 191715 241572
rect 197353 241634 197419 241637
rect 197353 241632 200284 241634
rect 197353 241576 197358 241632
rect 197414 241576 200284 241632
rect 197353 241574 200284 241576
rect 197353 241571 197419 241574
rect 57881 241498 57947 241501
rect 82951 241498 83017 241501
rect 84101 241498 84167 241501
rect 57881 241496 84167 241498
rect 57881 241440 57886 241496
rect 57942 241440 82956 241496
rect 83012 241440 84106 241496
rect 84162 241440 84167 241496
rect 57881 241438 84167 241440
rect 57881 241435 57947 241438
rect 82951 241435 83017 241438
rect 84101 241435 84167 241438
rect 149053 241498 149119 241501
rect 168373 241498 168439 241501
rect 149053 241496 168439 241498
rect 149053 241440 149058 241496
rect 149114 241440 168378 241496
rect 168434 241440 168439 241496
rect 149053 241438 168439 241440
rect 149053 241435 149119 241438
rect 168373 241435 168439 241438
rect 179045 241498 179111 241501
rect 198733 241498 198799 241501
rect 179045 241496 198799 241498
rect 179045 241440 179050 241496
rect 179106 241440 198738 241496
rect 198794 241440 198799 241496
rect 179045 241438 198799 241440
rect 179045 241435 179111 241438
rect 198733 241435 198799 241438
rect 244046 241365 244106 241604
rect 244046 241360 244155 241365
rect 244046 241304 244094 241360
rect 244150 241304 244155 241360
rect 244046 241302 244155 241304
rect 244089 241299 244155 241302
rect -960 241090 480 241180
rect 3417 241090 3483 241093
rect -960 241088 3483 241090
rect -960 241032 3422 241088
rect 3478 241032 3483 241088
rect -960 241030 3483 241032
rect -960 240940 480 241030
rect 3417 241027 3483 241030
rect 75361 240954 75427 240957
rect 126697 240954 126763 240957
rect 75361 240952 126763 240954
rect 75361 240896 75366 240952
rect 75422 240896 126702 240952
rect 126758 240896 126763 240952
rect 75361 240894 126763 240896
rect 75361 240891 75427 240894
rect 126697 240891 126763 240894
rect 69606 240756 69612 240820
rect 69676 240818 69682 240820
rect 122925 240818 122991 240821
rect 69676 240816 122991 240818
rect 69676 240760 122930 240816
rect 122986 240760 122991 240816
rect 69676 240758 122991 240760
rect 69676 240756 69682 240758
rect 122925 240755 122991 240758
rect 126237 240818 126303 240821
rect 149145 240818 149211 240821
rect 126237 240816 149211 240818
rect 126237 240760 126242 240816
rect 126298 240760 149150 240816
rect 149206 240760 149211 240816
rect 126237 240758 149211 240760
rect 126237 240755 126303 240758
rect 149145 240755 149211 240758
rect 197353 240818 197419 240821
rect 197353 240816 200284 240818
rect 197353 240760 197358 240816
rect 197414 240788 200284 240816
rect 197414 240760 200314 240788
rect 197353 240758 200314 240760
rect 197353 240755 197419 240758
rect 145925 240410 145991 240413
rect 154430 240410 154436 240412
rect 145925 240408 154436 240410
rect 145925 240352 145930 240408
rect 145986 240352 154436 240408
rect 145925 240350 154436 240352
rect 145925 240347 145991 240350
rect 154430 240348 154436 240350
rect 154500 240348 154506 240412
rect 200113 240410 200179 240413
rect 200254 240410 200314 240758
rect 243862 240549 243922 240788
rect 243862 240544 243971 240549
rect 243862 240488 243910 240544
rect 243966 240488 243971 240544
rect 243862 240486 243971 240488
rect 243905 240483 243971 240486
rect 200113 240408 200314 240410
rect 200113 240352 200118 240408
rect 200174 240352 200314 240408
rect 200113 240350 200314 240352
rect 200113 240347 200179 240350
rect 124305 240274 124371 240277
rect 178861 240274 178927 240277
rect 124305 240272 178927 240274
rect 124305 240216 124310 240272
rect 124366 240216 178866 240272
rect 178922 240216 178927 240272
rect 124305 240214 178927 240216
rect 124305 240211 124371 240214
rect 178861 240211 178927 240214
rect 198825 240274 198891 240277
rect 245878 240274 245884 240276
rect 198825 240272 199946 240274
rect 198825 240216 198830 240272
rect 198886 240216 199946 240272
rect 198825 240214 199946 240216
rect 244076 240214 245884 240274
rect 198825 240211 198891 240214
rect 43989 240138 44055 240141
rect 77293 240138 77359 240141
rect 77937 240138 78003 240141
rect 43989 240136 78003 240138
rect 43989 240080 43994 240136
rect 44050 240080 77298 240136
rect 77354 240080 77942 240136
rect 77998 240080 78003 240136
rect 43989 240078 78003 240080
rect 199886 240138 199946 240214
rect 245878 240212 245884 240214
rect 245948 240212 245954 240276
rect 200246 240138 200252 240140
rect 199886 240078 200252 240138
rect 43989 240075 44055 240078
rect 77293 240075 77359 240078
rect 77937 240075 78003 240078
rect 200246 240076 200252 240078
rect 200316 240076 200322 240140
rect 200430 240076 200436 240140
rect 200500 240138 200506 240140
rect 200941 240138 201007 240141
rect 200500 240136 201007 240138
rect 200500 240080 200946 240136
rect 201002 240080 201007 240136
rect 200500 240078 201007 240080
rect 200500 240076 200506 240078
rect 200941 240075 201007 240078
rect 218646 240076 218652 240140
rect 218716 240138 218722 240140
rect 219525 240138 219591 240141
rect 218716 240136 219591 240138
rect 218716 240080 219530 240136
rect 219586 240080 219591 240136
rect 218716 240078 219591 240080
rect 218716 240076 218722 240078
rect 219525 240075 219591 240078
rect 228214 240076 228220 240140
rect 228284 240138 228290 240140
rect 230565 240138 230631 240141
rect 228284 240136 230631 240138
rect 228284 240080 230570 240136
rect 230626 240080 230631 240136
rect 228284 240078 230631 240080
rect 228284 240076 228290 240078
rect 230565 240075 230631 240078
rect 233734 240076 233740 240140
rect 233804 240138 233810 240140
rect 236453 240138 236519 240141
rect 233804 240136 236519 240138
rect 233804 240080 236458 240136
rect 236514 240080 236519 240136
rect 233804 240078 236519 240080
rect 233804 240076 233810 240078
rect 236453 240075 236519 240078
rect 237925 240138 237991 240141
rect 238518 240138 238524 240140
rect 237925 240136 238524 240138
rect 237925 240080 237930 240136
rect 237986 240080 238524 240136
rect 237925 240078 238524 240080
rect 237925 240075 237991 240078
rect 238518 240076 238524 240078
rect 238588 240076 238594 240140
rect 258073 240138 258139 240141
rect 580165 240138 580231 240141
rect 258030 240136 580231 240138
rect 258030 240080 258078 240136
rect 258134 240080 580170 240136
rect 580226 240080 580231 240136
rect 258030 240078 580231 240080
rect 258030 240075 258139 240078
rect 580165 240075 580231 240078
rect 50889 240002 50955 240005
rect 74717 240002 74783 240005
rect 75453 240002 75519 240005
rect 50889 240000 75519 240002
rect 50889 239944 50894 240000
rect 50950 239944 74722 240000
rect 74778 239944 75458 240000
rect 75514 239944 75519 240000
rect 50889 239942 75519 239944
rect 50889 239939 50955 239942
rect 74717 239939 74783 239942
rect 75453 239939 75519 239942
rect 112529 240002 112595 240005
rect 222285 240002 222351 240005
rect 112529 240000 222351 240002
rect 112529 239944 112534 240000
rect 112590 239944 222290 240000
rect 222346 239944 222351 240000
rect 112529 239942 222351 239944
rect 112529 239939 112595 239942
rect 222285 239939 222351 239942
rect 239213 240002 239279 240005
rect 258030 240002 258090 240075
rect 239213 240000 258090 240002
rect 239213 239944 239218 240000
rect 239274 239944 258090 240000
rect 239213 239942 258090 239944
rect 239213 239939 239279 239942
rect 84009 239866 84075 239869
rect 84009 239864 200130 239866
rect 84009 239808 84014 239864
rect 84070 239808 200130 239864
rect 84009 239806 200130 239808
rect 84009 239803 84075 239806
rect 200070 239594 200130 239806
rect 200246 239668 200252 239732
rect 200316 239730 200322 239732
rect 200573 239730 200639 239733
rect 204897 239730 204963 239733
rect 200316 239728 204963 239730
rect 200316 239672 200578 239728
rect 200634 239672 204902 239728
rect 204958 239672 204963 239728
rect 200316 239670 204963 239672
rect 200316 239668 200322 239670
rect 200573 239667 200639 239670
rect 204897 239667 204963 239670
rect 222285 239730 222351 239733
rect 228357 239730 228423 239733
rect 222285 239728 228423 239730
rect 222285 239672 222290 239728
rect 222346 239672 228362 239728
rect 228418 239672 228423 239728
rect 222285 239670 228423 239672
rect 222285 239667 222351 239670
rect 228357 239667 228423 239670
rect 207933 239594 207999 239597
rect 200070 239592 207999 239594
rect 200070 239536 207938 239592
rect 207994 239536 207999 239592
rect 200070 239534 207999 239536
rect 207933 239531 207999 239534
rect 207974 239396 207980 239460
rect 208044 239458 208050 239460
rect 219433 239458 219499 239461
rect 208044 239456 219499 239458
rect 208044 239400 219438 239456
rect 219494 239400 219499 239456
rect 208044 239398 219499 239400
rect 208044 239396 208050 239398
rect 219433 239395 219499 239398
rect 219525 238914 219591 238917
rect 243629 238914 243695 238917
rect 219525 238912 243695 238914
rect 219525 238856 219530 238912
rect 219586 238856 243634 238912
rect 243690 238856 243695 238912
rect 219525 238854 243695 238856
rect 219525 238851 219591 238854
rect 243629 238851 243695 238854
rect 238937 238780 239003 238781
rect 238886 238778 238892 238780
rect 238846 238718 238892 238778
rect 238956 238776 239003 238780
rect 238998 238720 239003 238776
rect 238886 238716 238892 238718
rect 238956 238716 239003 238720
rect 238937 238715 239003 238716
rect 202045 238642 202111 238645
rect 203006 238642 203012 238644
rect 202045 238640 203012 238642
rect 202045 238584 202050 238640
rect 202106 238584 203012 238640
rect 202045 238582 203012 238584
rect 202045 238579 202111 238582
rect 203006 238580 203012 238582
rect 203076 238580 203082 238644
rect 212574 238580 212580 238644
rect 212644 238642 212650 238644
rect 213637 238642 213703 238645
rect 212644 238640 213703 238642
rect 212644 238584 213642 238640
rect 213698 238584 213703 238640
rect 212644 238582 213703 238584
rect 212644 238580 212650 238582
rect 213637 238579 213703 238582
rect 214046 238580 214052 238644
rect 214116 238642 214122 238644
rect 215201 238642 215267 238645
rect 214116 238640 215267 238642
rect 214116 238584 215206 238640
rect 215262 238584 215267 238640
rect 214116 238582 215267 238584
rect 214116 238580 214122 238582
rect 215201 238579 215267 238582
rect 232446 238580 232452 238644
rect 232516 238642 232522 238644
rect 235901 238642 235967 238645
rect 232516 238640 235967 238642
rect 232516 238584 235906 238640
rect 235962 238584 235967 238640
rect 232516 238582 235967 238584
rect 232516 238580 232522 238582
rect 235901 238579 235967 238582
rect 241789 238642 241855 238645
rect 258165 238642 258231 238645
rect 241789 238640 258231 238642
rect 241789 238584 241794 238640
rect 241850 238584 258170 238640
rect 258226 238584 258231 238640
rect 241789 238582 258231 238584
rect 241789 238579 241855 238582
rect 258165 238579 258231 238582
rect 96613 238506 96679 238509
rect 214189 238506 214255 238509
rect 96613 238504 214255 238506
rect 96613 238448 96618 238504
rect 96674 238448 214194 238504
rect 214250 238448 214255 238504
rect 96613 238446 214255 238448
rect 96613 238443 96679 238446
rect 214189 238443 214255 238446
rect 120257 238370 120323 238373
rect 226701 238370 226767 238373
rect 120257 238368 226767 238370
rect 120257 238312 120262 238368
rect 120318 238312 226706 238368
rect 226762 238312 226767 238368
rect 120257 238310 226767 238312
rect 120257 238307 120323 238310
rect 226701 238307 226767 238310
rect 73153 238234 73219 238237
rect 202229 238234 202295 238237
rect 73153 238232 202295 238234
rect 73153 238176 73158 238232
rect 73214 238176 202234 238232
rect 202290 238176 202295 238232
rect 73153 238174 202295 238176
rect 73153 238171 73219 238174
rect 202229 238171 202295 238174
rect 58985 237962 59051 237965
rect 75085 237962 75151 237965
rect 58985 237960 75151 237962
rect 58985 237904 58990 237960
rect 59046 237904 75090 237960
rect 75146 237904 75151 237960
rect 58985 237902 75151 237904
rect 58985 237899 59051 237902
rect 75085 237899 75151 237902
rect 234061 237554 234127 237557
rect 241789 237554 241855 237557
rect 242014 237554 242020 237556
rect 234061 237552 238770 237554
rect 234061 237496 234066 237552
rect 234122 237496 238770 237552
rect 234061 237494 238770 237496
rect 234061 237491 234127 237494
rect 220169 237418 220235 237421
rect 221365 237418 221431 237421
rect 220169 237416 221431 237418
rect 220169 237360 220174 237416
rect 220230 237360 221370 237416
rect 221426 237360 221431 237416
rect 220169 237358 221431 237360
rect 220169 237355 220235 237358
rect 221365 237355 221431 237358
rect 235257 237418 235323 237421
rect 237373 237418 237439 237421
rect 235257 237416 237439 237418
rect 235257 237360 235262 237416
rect 235318 237360 237378 237416
rect 237434 237360 237439 237416
rect 235257 237358 237439 237360
rect 238710 237418 238770 237494
rect 241789 237552 242020 237554
rect 241789 237496 241794 237552
rect 241850 237496 242020 237552
rect 241789 237494 242020 237496
rect 241789 237491 241855 237494
rect 242014 237492 242020 237494
rect 242084 237492 242090 237556
rect 307845 237418 307911 237421
rect 238710 237416 307911 237418
rect 238710 237360 307850 237416
rect 307906 237360 307911 237416
rect 238710 237358 307911 237360
rect 235257 237355 235323 237358
rect 237373 237355 237439 237358
rect 307845 237355 307911 237358
rect 137093 237284 137159 237285
rect 137093 237280 137140 237284
rect 137204 237282 137210 237284
rect 149053 237282 149119 237285
rect 155350 237282 155356 237284
rect 137093 237224 137098 237280
rect 137093 237220 137140 237224
rect 137204 237222 137250 237282
rect 149053 237280 155356 237282
rect 149053 237224 149058 237280
rect 149114 237224 155356 237280
rect 149053 237222 155356 237224
rect 137204 237220 137210 237222
rect 137093 237219 137159 237220
rect 149053 237219 149119 237222
rect 155350 237220 155356 237222
rect 155420 237220 155426 237284
rect 208894 237220 208900 237284
rect 208964 237282 208970 237284
rect 214557 237282 214623 237285
rect 208964 237280 214623 237282
rect 208964 237224 214562 237280
rect 214618 237224 214623 237280
rect 208964 237222 214623 237224
rect 208964 237220 208970 237222
rect 214557 237219 214623 237222
rect 216581 237282 216647 237285
rect 583477 237282 583543 237285
rect 216581 237280 583543 237282
rect 216581 237224 216586 237280
rect 216642 237224 583482 237280
rect 583538 237224 583543 237280
rect 216581 237222 583543 237224
rect 216581 237219 216647 237222
rect 583477 237219 583543 237222
rect 60549 237146 60615 237149
rect 226885 237146 226951 237149
rect 60549 237144 226951 237146
rect 60549 237088 60554 237144
rect 60610 237088 226890 237144
rect 226946 237088 226951 237144
rect 60549 237086 226951 237088
rect 60549 237083 60615 237086
rect 226885 237083 226951 237086
rect 162761 237010 162827 237013
rect 240685 237010 240751 237013
rect 162761 237008 240751 237010
rect 162761 236952 162766 237008
rect 162822 236952 240690 237008
rect 240746 236952 240751 237008
rect 162761 236950 240751 236952
rect 162761 236947 162827 236950
rect 240685 236947 240751 236950
rect 137093 236874 137159 236877
rect 178953 236874 179019 236877
rect 137093 236872 179019 236874
rect 137093 236816 137098 236872
rect 137154 236816 178958 236872
rect 179014 236816 179019 236872
rect 137093 236814 179019 236816
rect 137093 236811 137159 236814
rect 178953 236811 179019 236814
rect 67357 236602 67423 236605
rect 133597 236602 133663 236605
rect 67357 236600 133663 236602
rect 67357 236544 67362 236600
rect 67418 236544 133602 236600
rect 133658 236544 133663 236600
rect 67357 236542 133663 236544
rect 67357 236539 67423 236542
rect 133597 236539 133663 236542
rect 216029 236058 216095 236061
rect 216581 236058 216647 236061
rect 216029 236056 216647 236058
rect 216029 236000 216034 236056
rect 216090 236000 216586 236056
rect 216642 236000 216647 236056
rect 216029 235998 216647 236000
rect 216029 235995 216095 235998
rect 216581 235995 216647 235998
rect 66161 235922 66227 235925
rect 245837 235922 245903 235925
rect 66161 235920 245903 235922
rect 66161 235864 66166 235920
rect 66222 235864 245842 235920
rect 245898 235864 245903 235920
rect 66161 235862 245903 235864
rect 66161 235859 66227 235862
rect 245837 235859 245903 235862
rect 252502 235860 252508 235924
rect 252572 235922 252578 235924
rect 252921 235922 252987 235925
rect 252572 235920 252987 235922
rect 252572 235864 252926 235920
rect 252982 235864 252987 235920
rect 252572 235862 252987 235864
rect 252572 235860 252578 235862
rect 252921 235859 252987 235862
rect 48129 235786 48195 235789
rect 119337 235786 119403 235789
rect 48129 235784 119403 235786
rect 48129 235728 48134 235784
rect 48190 235728 119342 235784
rect 119398 235728 119403 235784
rect 48129 235726 119403 235728
rect 48129 235723 48195 235726
rect 119337 235723 119403 235726
rect 142337 235786 142403 235789
rect 159214 235786 159220 235788
rect 142337 235784 159220 235786
rect 142337 235728 142342 235784
rect 142398 235728 159220 235784
rect 142337 235726 159220 235728
rect 142337 235723 142403 235726
rect 159214 235724 159220 235726
rect 159284 235724 159290 235788
rect 178677 235786 178743 235789
rect 242709 235786 242775 235789
rect 178677 235784 242775 235786
rect 178677 235728 178682 235784
rect 178738 235728 242714 235784
rect 242770 235728 242775 235784
rect 178677 235726 242775 235728
rect 178677 235723 178743 235726
rect 242709 235723 242775 235726
rect 72366 235588 72372 235652
rect 72436 235650 72442 235652
rect 102133 235650 102199 235653
rect 72436 235648 102199 235650
rect 72436 235592 102138 235648
rect 102194 235592 102199 235648
rect 72436 235590 102199 235592
rect 72436 235588 72442 235590
rect 102133 235587 102199 235590
rect 136633 235650 136699 235653
rect 195278 235650 195284 235652
rect 136633 235648 195284 235650
rect 136633 235592 136638 235648
rect 136694 235592 195284 235648
rect 136633 235590 195284 235592
rect 136633 235587 136699 235590
rect 195278 235588 195284 235590
rect 195348 235588 195354 235652
rect 196566 235588 196572 235652
rect 196636 235650 196642 235652
rect 211061 235650 211127 235653
rect 232589 235650 232655 235653
rect 196636 235590 200130 235650
rect 196636 235588 196642 235590
rect 200070 235514 200130 235590
rect 211061 235648 232655 235650
rect 211061 235592 211066 235648
rect 211122 235592 232594 235648
rect 232650 235592 232655 235648
rect 211061 235590 232655 235592
rect 211061 235587 211127 235590
rect 232589 235587 232655 235590
rect 210325 235514 210391 235517
rect 200070 235512 210391 235514
rect 200070 235456 210330 235512
rect 210386 235456 210391 235512
rect 200070 235454 210391 235456
rect 210325 235451 210391 235454
rect 102133 234698 102199 234701
rect 102777 234698 102843 234701
rect 102133 234696 102843 234698
rect 102133 234640 102138 234696
rect 102194 234640 102782 234696
rect 102838 234640 102843 234696
rect 102133 234638 102843 234640
rect 102133 234635 102199 234638
rect 102777 234635 102843 234638
rect 136633 234698 136699 234701
rect 137369 234698 137435 234701
rect 136633 234696 137435 234698
rect 136633 234640 136638 234696
rect 136694 234640 137374 234696
rect 137430 234640 137435 234696
rect 136633 234638 137435 234640
rect 136633 234635 136699 234638
rect 137369 234635 137435 234638
rect 75085 234562 75151 234565
rect 169201 234562 169267 234565
rect 75085 234560 169267 234562
rect 75085 234504 75090 234560
rect 75146 234504 169206 234560
rect 169262 234504 169267 234560
rect 75085 234502 169267 234504
rect 75085 234499 75151 234502
rect 169201 234499 169267 234502
rect 181437 234562 181503 234565
rect 228173 234562 228239 234565
rect 229093 234562 229159 234565
rect 181437 234560 228239 234562
rect 181437 234504 181442 234560
rect 181498 234504 228178 234560
rect 228234 234504 228239 234560
rect 181437 234502 228239 234504
rect 181437 234499 181503 234502
rect 228173 234499 228239 234502
rect 229050 234560 229159 234562
rect 229050 234504 229098 234560
rect 229154 234504 229159 234560
rect 229050 234499 229159 234504
rect 150433 234426 150499 234429
rect 163589 234426 163655 234429
rect 150433 234424 163655 234426
rect 150433 234368 150438 234424
rect 150494 234368 163594 234424
rect 163650 234368 163655 234424
rect 150433 234366 163655 234368
rect 150433 234363 150499 234366
rect 163589 234363 163655 234366
rect 195513 234426 195579 234429
rect 203517 234426 203583 234429
rect 204069 234426 204135 234429
rect 195513 234424 204135 234426
rect 195513 234368 195518 234424
rect 195574 234368 203522 234424
rect 203578 234368 204074 234424
rect 204130 234368 204135 234424
rect 195513 234366 204135 234368
rect 195513 234363 195579 234366
rect 203517 234363 203583 234366
rect 204069 234363 204135 234366
rect 69790 234228 69796 234292
rect 69860 234290 69866 234292
rect 153837 234290 153903 234293
rect 69860 234288 153903 234290
rect 69860 234232 153842 234288
rect 153898 234232 153903 234288
rect 69860 234230 153903 234232
rect 69860 234228 69866 234230
rect 153837 234227 153903 234230
rect 164969 233882 165035 233885
rect 195145 233882 195211 233885
rect 164969 233880 195211 233882
rect 164969 233824 164974 233880
rect 165030 233824 195150 233880
rect 195206 233824 195211 233880
rect 164969 233822 195211 233824
rect 164969 233819 165035 233822
rect 195145 233819 195211 233822
rect 201585 233882 201651 233885
rect 224217 233882 224283 233885
rect 201585 233880 224283 233882
rect 201585 233824 201590 233880
rect 201646 233824 224222 233880
rect 224278 233824 224283 233880
rect 201585 233822 224283 233824
rect 201585 233819 201651 233822
rect 224217 233819 224283 233822
rect 227713 233882 227779 233885
rect 229050 233882 229110 234499
rect 231117 234018 231183 234021
rect 240358 234018 240364 234020
rect 231117 234016 240364 234018
rect 231117 233960 231122 234016
rect 231178 233960 240364 234016
rect 231117 233958 240364 233960
rect 231117 233955 231183 233958
rect 240358 233956 240364 233958
rect 240428 233956 240434 234020
rect 287237 233882 287303 233885
rect 227713 233880 287303 233882
rect 227713 233824 227718 233880
rect 227774 233824 287242 233880
rect 287298 233824 287303 233880
rect 227713 233822 287303 233824
rect 227713 233819 227779 233822
rect 287237 233819 287303 233822
rect 61837 233202 61903 233205
rect 234981 233202 235047 233205
rect 61837 233200 235047 233202
rect 61837 233144 61842 233200
rect 61898 233144 234986 233200
rect 235042 233144 235047 233200
rect 61837 233142 235047 233144
rect 61837 233139 61903 233142
rect 234981 233139 235047 233142
rect 130377 233066 130443 233069
rect 132534 233066 132540 233068
rect 130377 233064 132540 233066
rect 130377 233008 130382 233064
rect 130438 233008 132540 233064
rect 130377 233006 132540 233008
rect 130377 233003 130443 233006
rect 132534 233004 132540 233006
rect 132604 233004 132610 233068
rect 151813 233066 151879 233069
rect 173801 233066 173867 233069
rect 238845 233066 238911 233069
rect 151813 233064 161490 233066
rect 151813 233008 151818 233064
rect 151874 233008 161490 233064
rect 151813 233006 161490 233008
rect 151813 233003 151879 233006
rect 74717 232930 74783 232933
rect 157333 232930 157399 232933
rect 74717 232928 157399 232930
rect 74717 232872 74722 232928
rect 74778 232872 157338 232928
rect 157394 232872 157399 232928
rect 74717 232870 157399 232872
rect 74717 232867 74783 232870
rect 157333 232867 157399 232870
rect 161430 232794 161490 233006
rect 173801 233064 238911 233066
rect 173801 233008 173806 233064
rect 173862 233008 238850 233064
rect 238906 233008 238911 233064
rect 173801 233006 238911 233008
rect 173801 233003 173867 233006
rect 238845 233003 238911 233006
rect 171869 232930 171935 232933
rect 194685 232930 194751 232933
rect 171869 232928 194751 232930
rect 171869 232872 171874 232928
rect 171930 232872 194690 232928
rect 194746 232872 194751 232928
rect 171869 232870 194751 232872
rect 171869 232867 171935 232870
rect 194685 232867 194751 232870
rect 195145 232930 195211 232933
rect 230197 232930 230263 232933
rect 195145 232928 230263 232930
rect 195145 232872 195150 232928
rect 195206 232872 230202 232928
rect 230258 232872 230263 232928
rect 195145 232870 230263 232872
rect 195145 232867 195211 232870
rect 230197 232867 230263 232870
rect 173157 232794 173223 232797
rect 161430 232792 173223 232794
rect 161430 232736 173162 232792
rect 173218 232736 173223 232792
rect 161430 232734 173223 232736
rect 173157 232731 173223 232734
rect 582649 232386 582715 232389
rect 583520 232386 584960 232476
rect 582649 232384 584960 232386
rect 582649 232328 582654 232384
rect 582710 232328 584960 232384
rect 582649 232326 584960 232328
rect 582649 232323 582715 232326
rect 583520 232236 584960 232326
rect 49601 231842 49667 231845
rect 231485 231842 231551 231845
rect 49601 231840 231551 231842
rect 49601 231784 49606 231840
rect 49662 231784 231490 231840
rect 231546 231784 231551 231840
rect 49601 231782 231551 231784
rect 49601 231779 49667 231782
rect 231485 231779 231551 231782
rect 128169 231706 128235 231709
rect 227713 231706 227779 231709
rect 128169 231704 227779 231706
rect 128169 231648 128174 231704
rect 128230 231648 227718 231704
rect 227774 231648 227779 231704
rect 128169 231646 227779 231648
rect 128169 231643 128235 231646
rect 227713 231643 227779 231646
rect 189809 231570 189875 231573
rect 247217 231570 247283 231573
rect 189809 231568 247283 231570
rect 189809 231512 189814 231568
rect 189870 231512 247222 231568
rect 247278 231512 247283 231568
rect 189809 231510 247283 231512
rect 189809 231507 189875 231510
rect 247217 231507 247283 231510
rect 114369 231162 114435 231165
rect 143441 231162 143507 231165
rect 143574 231162 143580 231164
rect 114369 231160 143580 231162
rect 114369 231104 114374 231160
rect 114430 231104 143446 231160
rect 143502 231104 143580 231160
rect 114369 231102 143580 231104
rect 114369 231099 114435 231102
rect 143441 231099 143507 231102
rect 143574 231100 143580 231102
rect 143644 231100 143650 231164
rect 66069 230482 66135 230485
rect 185761 230482 185827 230485
rect 66069 230480 185827 230482
rect 66069 230424 66074 230480
rect 66130 230424 185766 230480
rect 185822 230424 185827 230480
rect 66069 230422 185827 230424
rect 66069 230419 66135 230422
rect 185761 230419 185827 230422
rect 187693 230482 187759 230485
rect 216622 230482 216628 230484
rect 187693 230480 216628 230482
rect 187693 230424 187698 230480
rect 187754 230424 216628 230480
rect 187693 230422 216628 230424
rect 187693 230419 187759 230422
rect 216622 230420 216628 230422
rect 216692 230420 216698 230484
rect 72969 230346 73035 230349
rect 154062 230346 154068 230348
rect 72969 230344 154068 230346
rect 72969 230288 72974 230344
rect 73030 230288 154068 230344
rect 72969 230286 154068 230288
rect 72969 230283 73035 230286
rect 154062 230284 154068 230286
rect 154132 230284 154138 230348
rect 163497 230346 163563 230349
rect 245694 230346 245700 230348
rect 161430 230344 245700 230346
rect 161430 230288 163502 230344
rect 163558 230288 245700 230344
rect 161430 230286 245700 230288
rect 129549 230210 129615 230213
rect 161430 230210 161490 230286
rect 163497 230283 163563 230286
rect 245694 230284 245700 230286
rect 245764 230284 245770 230348
rect 129549 230208 161490 230210
rect 129549 230152 129554 230208
rect 129610 230152 161490 230208
rect 129549 230150 161490 230152
rect 129549 230147 129615 230150
rect 200297 229802 200363 229805
rect 303705 229802 303771 229805
rect 200297 229800 303771 229802
rect 200297 229744 200302 229800
rect 200358 229744 303710 229800
rect 303766 229744 303771 229800
rect 200297 229742 303771 229744
rect 200297 229739 200363 229742
rect 303705 229739 303771 229742
rect 67950 228924 67956 228988
rect 68020 228986 68026 228988
rect 233509 228986 233575 228989
rect 68020 228984 233575 228986
rect 68020 228928 233514 228984
rect 233570 228928 233575 228984
rect 68020 228926 233575 228928
rect 68020 228924 68026 228926
rect 233509 228923 233575 228926
rect 102777 228850 102843 228853
rect 232957 228850 233023 228853
rect 102777 228848 233023 228850
rect 102777 228792 102782 228848
rect 102838 228792 232962 228848
rect 233018 228792 233023 228848
rect 102777 228790 233023 228792
rect 102777 228787 102843 228790
rect 232957 228787 233023 228790
rect 79317 228714 79383 228717
rect 201493 228714 201559 228717
rect 79317 228712 201559 228714
rect 79317 228656 79322 228712
rect 79378 228656 201498 228712
rect 201554 228656 201559 228712
rect 79317 228654 201559 228656
rect 79317 228651 79383 228654
rect 201493 228651 201559 228654
rect 233877 228306 233943 228309
rect 243261 228306 243327 228309
rect 233877 228304 243327 228306
rect 233877 228248 233882 228304
rect 233938 228248 243266 228304
rect 243322 228248 243327 228304
rect 233877 228246 243327 228248
rect 233877 228243 233943 228246
rect 243261 228243 243327 228246
rect -960 227884 480 228124
rect 84694 227564 84700 227628
rect 84764 227626 84770 227628
rect 245878 227626 245884 227628
rect 84764 227566 245884 227626
rect 84764 227564 84770 227566
rect 245878 227564 245884 227566
rect 245948 227564 245954 227628
rect 86718 227428 86724 227492
rect 86788 227490 86794 227492
rect 216029 227490 216095 227493
rect 86788 227488 216095 227490
rect 86788 227432 216034 227488
rect 216090 227432 216095 227488
rect 86788 227430 216095 227432
rect 86788 227428 86794 227430
rect 216029 227427 216095 227430
rect 128997 227354 129063 227357
rect 159449 227354 159515 227357
rect 128997 227352 159515 227354
rect 128997 227296 129002 227352
rect 129058 227296 159454 227352
rect 159510 227296 159515 227352
rect 128997 227294 159515 227296
rect 128997 227291 129063 227294
rect 159449 227291 159515 227294
rect 191741 226946 191807 226949
rect 282269 226946 282335 226949
rect 191741 226944 282335 226946
rect 191741 226888 191746 226944
rect 191802 226888 282274 226944
rect 282330 226888 282335 226944
rect 191741 226886 282335 226888
rect 191741 226883 191807 226886
rect 282269 226883 282335 226886
rect 215937 226404 216003 226405
rect 215886 226402 215892 226404
rect 215846 226342 215892 226402
rect 215956 226400 216003 226404
rect 215998 226344 216003 226400
rect 215886 226340 215892 226342
rect 215956 226340 216003 226344
rect 215937 226339 216003 226340
rect 52269 226266 52335 226269
rect 227621 226266 227687 226269
rect 52269 226264 227687 226266
rect 52269 226208 52274 226264
rect 52330 226208 227626 226264
rect 227682 226208 227687 226264
rect 52269 226206 227687 226208
rect 52269 226203 52335 226206
rect 227621 226203 227687 226206
rect 146753 226130 146819 226133
rect 165521 226130 165587 226133
rect 204989 226130 205055 226133
rect 146753 226128 205055 226130
rect 146753 226072 146758 226128
rect 146814 226072 165526 226128
rect 165582 226072 204994 226128
rect 205050 226072 205055 226128
rect 146753 226070 205055 226072
rect 146753 226067 146819 226070
rect 165521 226067 165587 226070
rect 204989 226067 205055 226070
rect 191281 225994 191347 225997
rect 223614 225994 223620 225996
rect 191281 225992 223620 225994
rect 191281 225936 191286 225992
rect 191342 225936 223620 225992
rect 191281 225934 223620 225936
rect 191281 225931 191347 225934
rect 223614 225932 223620 225934
rect 223684 225994 223690 225996
rect 224861 225994 224927 225997
rect 223684 225992 224927 225994
rect 223684 225936 224866 225992
rect 224922 225936 224927 225992
rect 223684 225934 224927 225936
rect 223684 225932 223690 225934
rect 224861 225931 224927 225934
rect 137461 225586 137527 225589
rect 155493 225586 155559 225589
rect 137461 225584 155559 225586
rect 137461 225528 137466 225584
rect 137522 225528 155498 225584
rect 155554 225528 155559 225584
rect 137461 225526 155559 225528
rect 137461 225523 137527 225526
rect 155493 225523 155559 225526
rect 230238 225116 230244 225180
rect 230308 225178 230314 225180
rect 234613 225178 234679 225181
rect 230308 225176 234679 225178
rect 230308 225120 234618 225176
rect 234674 225120 234679 225176
rect 230308 225118 234679 225120
rect 230308 225116 230314 225118
rect 234613 225115 234679 225118
rect 119429 225042 119495 225045
rect 135161 225042 135227 225045
rect 119429 225040 135227 225042
rect 119429 224984 119434 225040
rect 119490 224984 135166 225040
rect 135222 224984 135227 225040
rect 119429 224982 135227 224984
rect 119429 224979 119495 224982
rect 135161 224979 135227 224982
rect 212165 225042 212231 225045
rect 215385 225042 215451 225045
rect 582649 225042 582715 225045
rect 212165 225040 582715 225042
rect 212165 224984 212170 225040
rect 212226 224984 215390 225040
rect 215446 224984 582654 225040
rect 582710 224984 582715 225040
rect 212165 224982 582715 224984
rect 212165 224979 212231 224982
rect 215385 224979 215451 224982
rect 582649 224979 582715 224982
rect 64597 224906 64663 224909
rect 263593 224906 263659 224909
rect 64597 224904 263659 224906
rect 64597 224848 64602 224904
rect 64658 224848 263598 224904
rect 263654 224848 263659 224904
rect 64597 224846 263659 224848
rect 64597 224843 64663 224846
rect 263593 224843 263659 224846
rect 84101 224770 84167 224773
rect 239765 224770 239831 224773
rect 244273 224772 244339 224773
rect 84101 224768 239831 224770
rect 84101 224712 84106 224768
rect 84162 224712 239770 224768
rect 239826 224712 239831 224768
rect 84101 224710 239831 224712
rect 84101 224707 84167 224710
rect 239765 224707 239831 224710
rect 244222 224708 244228 224772
rect 244292 224770 244339 224772
rect 244292 224768 244384 224770
rect 244334 224712 244384 224768
rect 244292 224710 244384 224712
rect 244292 224708 244339 224710
rect 244273 224707 244339 224708
rect 156597 224634 156663 224637
rect 226977 224634 227043 224637
rect 156597 224632 227043 224634
rect 156597 224576 156602 224632
rect 156658 224576 226982 224632
rect 227038 224576 227043 224632
rect 156597 224574 227043 224576
rect 156597 224571 156663 224574
rect 226977 224571 227043 224574
rect 263593 224498 263659 224501
rect 264237 224498 264303 224501
rect 263593 224496 264303 224498
rect 263593 224440 263598 224496
rect 263654 224440 264242 224496
rect 264298 224440 264303 224496
rect 263593 224438 264303 224440
rect 263593 224435 263659 224438
rect 264237 224435 264303 224438
rect 51717 224226 51783 224229
rect 150382 224226 150388 224228
rect 51717 224224 150388 224226
rect 51717 224168 51722 224224
rect 51778 224168 150388 224224
rect 51717 224166 150388 224168
rect 51717 224163 51783 224166
rect 150382 224164 150388 224166
rect 150452 224164 150458 224228
rect 60457 223546 60523 223549
rect 163681 223546 163747 223549
rect 60457 223544 163747 223546
rect 60457 223488 60462 223544
rect 60518 223488 163686 223544
rect 163742 223488 163747 223544
rect 60457 223486 163747 223488
rect 60457 223483 60523 223486
rect 163681 223483 163747 223486
rect 158069 223138 158135 223141
rect 158713 223138 158779 223141
rect 251214 223138 251220 223140
rect 158069 223136 251220 223138
rect 158069 223080 158074 223136
rect 158130 223080 158718 223136
rect 158774 223080 251220 223136
rect 158069 223078 251220 223080
rect 158069 223075 158135 223078
rect 158713 223075 158779 223078
rect 251214 223076 251220 223078
rect 251284 223076 251290 223140
rect 36537 223002 36603 223005
rect 156597 223002 156663 223005
rect 36537 223000 156663 223002
rect 36537 222944 36542 223000
rect 36598 222944 156602 223000
rect 156658 222944 156663 223000
rect 36537 222942 156663 222944
rect 36537 222939 36603 222942
rect 156597 222939 156663 222942
rect 195421 223002 195487 223005
rect 200205 223002 200271 223005
rect 302417 223002 302483 223005
rect 195421 223000 302483 223002
rect 195421 222944 195426 223000
rect 195482 222944 200210 223000
rect 200266 222944 302422 223000
rect 302478 222944 302483 223000
rect 195421 222942 302483 222944
rect 195421 222939 195487 222942
rect 200205 222939 200271 222942
rect 302417 222939 302483 222942
rect 77201 222866 77267 222869
rect 202781 222866 202847 222869
rect 203057 222866 203123 222869
rect 77201 222864 203123 222866
rect 77201 222808 77206 222864
rect 77262 222808 202786 222864
rect 202842 222808 203062 222864
rect 203118 222808 203123 222864
rect 77201 222806 203123 222808
rect 77201 222803 77267 222806
rect 202781 222803 202847 222806
rect 203057 222803 203123 222806
rect 216622 222804 216628 222868
rect 216692 222866 216698 222868
rect 227713 222866 227779 222869
rect 216692 222864 227779 222866
rect 216692 222808 227718 222864
rect 227774 222808 227779 222864
rect 216692 222806 227779 222808
rect 216692 222804 216698 222806
rect 227713 222803 227779 222806
rect 125409 222186 125475 222189
rect 214097 222186 214163 222189
rect 125409 222184 214163 222186
rect 125409 222128 125414 222184
rect 125470 222128 214102 222184
rect 214158 222128 214163 222184
rect 125409 222126 214163 222128
rect 125409 222123 125475 222126
rect 214097 222123 214163 222126
rect 137277 222050 137343 222053
rect 171133 222050 171199 222053
rect 187693 222050 187759 222053
rect 137277 222048 187759 222050
rect 137277 221992 137282 222048
rect 137338 221992 171138 222048
rect 171194 221992 187698 222048
rect 187754 221992 187759 222048
rect 137277 221990 187759 221992
rect 137277 221987 137343 221990
rect 171133 221987 171199 221990
rect 187693 221987 187759 221990
rect 191097 221642 191163 221645
rect 245745 221642 245811 221645
rect 191097 221640 245811 221642
rect 191097 221584 191102 221640
rect 191158 221584 245750 221640
rect 245806 221584 245811 221640
rect 191097 221582 245811 221584
rect 191097 221579 191163 221582
rect 245745 221579 245811 221582
rect 101949 221506 102015 221509
rect 196617 221506 196683 221509
rect 101949 221504 196683 221506
rect 101949 221448 101954 221504
rect 102010 221448 196622 221504
rect 196678 221448 196683 221504
rect 101949 221446 196683 221448
rect 101949 221443 102015 221446
rect 196617 221443 196683 221446
rect 59077 220826 59143 220829
rect 193806 220826 193812 220828
rect 59077 220824 193812 220826
rect 59077 220768 59082 220824
rect 59138 220768 193812 220824
rect 59077 220766 193812 220768
rect 59077 220763 59143 220766
rect 193806 220764 193812 220766
rect 193876 220764 193882 220828
rect 204805 220826 204871 220829
rect 205357 220826 205423 220829
rect 204805 220824 205423 220826
rect 204805 220768 204810 220824
rect 204866 220768 205362 220824
rect 205418 220768 205423 220824
rect 204805 220766 205423 220768
rect 204805 220763 204871 220766
rect 205357 220763 205423 220766
rect 73797 220690 73863 220693
rect 159357 220690 159423 220693
rect 73797 220688 159423 220690
rect 73797 220632 73802 220688
rect 73858 220632 159362 220688
rect 159418 220632 159423 220688
rect 73797 220630 159423 220632
rect 73797 220627 73863 220630
rect 159357 220627 159423 220630
rect 192477 220282 192543 220285
rect 207749 220282 207815 220285
rect 192477 220280 207815 220282
rect 192477 220224 192482 220280
rect 192538 220224 207754 220280
rect 207810 220224 207815 220280
rect 192477 220222 207815 220224
rect 192477 220219 192543 220222
rect 207749 220219 207815 220222
rect 90909 220146 90975 220149
rect 298093 220146 298159 220149
rect 90909 220144 298159 220146
rect 90909 220088 90914 220144
rect 90970 220088 298098 220144
rect 298154 220088 298159 220144
rect 90909 220086 298159 220088
rect 90909 220083 90975 220086
rect 298093 220083 298159 220086
rect 204805 219466 204871 219469
rect 280286 219466 280292 219468
rect 204805 219464 280292 219466
rect 204805 219408 204810 219464
rect 204866 219408 280292 219464
rect 204805 219406 280292 219408
rect 204805 219403 204871 219406
rect 280286 219404 280292 219406
rect 280356 219404 280362 219468
rect 128261 219330 128327 219333
rect 152457 219330 152523 219333
rect 128261 219328 152523 219330
rect 128261 219272 128266 219328
rect 128322 219272 152462 219328
rect 152518 219272 152523 219328
rect 128261 219270 152523 219272
rect 128261 219267 128327 219270
rect 152457 219267 152523 219270
rect 199469 219330 199535 219333
rect 223389 219330 223455 219333
rect 199469 219328 223455 219330
rect 199469 219272 199474 219328
rect 199530 219272 223394 219328
rect 223450 219272 223455 219328
rect 199469 219270 223455 219272
rect 199469 219267 199535 219270
rect 223389 219267 223455 219270
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect 82721 218786 82787 218789
rect 162301 218786 162367 218789
rect 82721 218784 162367 218786
rect 82721 218728 82726 218784
rect 82782 218728 162306 218784
rect 162362 218728 162367 218784
rect 82721 218726 162367 218728
rect 82721 218723 82787 218726
rect 162301 218723 162367 218726
rect 163037 218786 163103 218789
rect 204805 218786 204871 218789
rect 163037 218784 204871 218786
rect 163037 218728 163042 218784
rect 163098 218728 204810 218784
rect 204866 218728 204871 218784
rect 163037 218726 204871 218728
rect 163037 218723 163103 218726
rect 204805 218723 204871 218726
rect 111609 218650 111675 218653
rect 306465 218650 306531 218653
rect 111609 218648 306531 218650
rect 111609 218592 111614 218648
rect 111670 218592 306470 218648
rect 306526 218592 306531 218648
rect 111609 218590 306531 218592
rect 111609 218587 111675 218590
rect 306465 218587 306531 218590
rect 222929 218242 222995 218245
rect 223389 218242 223455 218245
rect 222929 218240 223455 218242
rect 222929 218184 222934 218240
rect 222990 218184 223394 218240
rect 223450 218184 223455 218240
rect 222929 218182 223455 218184
rect 222929 218179 222995 218182
rect 223389 218179 223455 218182
rect 207381 218106 207447 218109
rect 283005 218106 283071 218109
rect 207381 218104 283071 218106
rect 207381 218048 207386 218104
rect 207442 218048 283010 218104
rect 283066 218048 283071 218104
rect 207381 218046 283071 218048
rect 207381 218043 207447 218046
rect 283005 218043 283071 218046
rect 122649 217970 122715 217973
rect 225597 217970 225663 217973
rect 122649 217968 225663 217970
rect 122649 217912 122654 217968
rect 122710 217912 225602 217968
rect 225658 217912 225663 217968
rect 122649 217910 225663 217912
rect 122649 217907 122715 217910
rect 225597 217907 225663 217910
rect 93853 217834 93919 217837
rect 158253 217834 158319 217837
rect 93853 217832 158319 217834
rect 93853 217776 93858 217832
rect 93914 217776 158258 217832
rect 158314 217776 158319 217832
rect 93853 217774 158319 217776
rect 93853 217771 93919 217774
rect 158253 217771 158319 217774
rect 64689 217290 64755 217293
rect 342253 217290 342319 217293
rect 64689 217288 342319 217290
rect 64689 217232 64694 217288
rect 64750 217232 342258 217288
rect 342314 217232 342319 217288
rect 64689 217230 342319 217232
rect 64689 217227 64755 217230
rect 342253 217227 342319 217230
rect 231853 216748 231919 216749
rect 231853 216746 231900 216748
rect 231808 216744 231900 216746
rect 231808 216688 231858 216744
rect 231808 216686 231900 216688
rect 231853 216684 231900 216686
rect 231964 216684 231970 216748
rect 231853 216683 231919 216684
rect 108297 216610 108363 216613
rect 195421 216610 195487 216613
rect 108297 216608 195487 216610
rect 108297 216552 108302 216608
rect 108358 216552 195426 216608
rect 195482 216552 195487 216608
rect 108297 216550 195487 216552
rect 108297 216547 108363 216550
rect 195421 216547 195487 216550
rect 204989 216202 205055 216205
rect 242249 216202 242315 216205
rect 204989 216200 242315 216202
rect 204989 216144 204994 216200
rect 205050 216144 242254 216200
rect 242310 216144 242315 216200
rect 204989 216142 242315 216144
rect 204989 216139 205055 216142
rect 242249 216139 242315 216142
rect 197169 216066 197235 216069
rect 276749 216066 276815 216069
rect 197169 216064 276815 216066
rect 197169 216008 197174 216064
rect 197230 216008 276754 216064
rect 276810 216008 276815 216064
rect 197169 216006 276815 216008
rect 197169 216003 197235 216006
rect 276749 216003 276815 216006
rect 67265 215930 67331 215933
rect 356053 215930 356119 215933
rect 67265 215928 356119 215930
rect 67265 215872 67270 215928
rect 67326 215872 356058 215928
rect 356114 215872 356119 215928
rect 67265 215870 356119 215872
rect 67265 215867 67331 215870
rect 356053 215867 356119 215870
rect 69749 215250 69815 215253
rect 226333 215250 226399 215253
rect 69749 215248 226399 215250
rect 69749 215192 69754 215248
rect 69810 215192 226338 215248
rect 226394 215192 226399 215248
rect 69749 215190 226399 215192
rect 69749 215187 69815 215190
rect 226333 215187 226399 215190
rect -960 214978 480 215068
rect 3325 214978 3391 214981
rect -960 214976 3391 214978
rect -960 214920 3330 214976
rect 3386 214920 3391 214976
rect -960 214918 3391 214920
rect -960 214828 480 214918
rect 3325 214915 3391 214918
rect 226333 214842 226399 214845
rect 226977 214842 227043 214845
rect 226333 214840 227043 214842
rect 226333 214784 226338 214840
rect 226394 214784 226982 214840
rect 227038 214784 227043 214840
rect 226333 214782 227043 214784
rect 226333 214779 226399 214782
rect 226977 214779 227043 214782
rect 111701 214706 111767 214709
rect 191189 214706 191255 214709
rect 111701 214704 191255 214706
rect 111701 214648 111706 214704
rect 111762 214648 191194 214704
rect 191250 214648 191255 214704
rect 111701 214646 191255 214648
rect 111701 214643 111767 214646
rect 191189 214643 191255 214646
rect 93761 214570 93827 214573
rect 299606 214570 299612 214572
rect 93761 214568 299612 214570
rect 93761 214512 93766 214568
rect 93822 214512 299612 214568
rect 93761 214510 299612 214512
rect 93761 214507 93827 214510
rect 299606 214508 299612 214510
rect 299676 214508 299682 214572
rect 53465 213890 53531 213893
rect 156597 213890 156663 213893
rect 156781 213890 156847 213893
rect 53465 213888 156847 213890
rect 53465 213832 53470 213888
rect 53526 213832 156602 213888
rect 156658 213832 156786 213888
rect 156842 213832 156847 213888
rect 53465 213830 156847 213832
rect 53465 213827 53531 213830
rect 156597 213827 156663 213830
rect 156781 213827 156847 213830
rect 217409 213890 217475 213893
rect 221917 213890 221983 213893
rect 217409 213888 221983 213890
rect 217409 213832 217414 213888
rect 217470 213832 221922 213888
rect 221978 213832 221983 213888
rect 217409 213830 221983 213832
rect 217409 213827 217475 213830
rect 221917 213827 221983 213830
rect 122741 213346 122807 213349
rect 180057 213346 180123 213349
rect 122741 213344 180123 213346
rect 122741 213288 122746 213344
rect 122802 213288 180062 213344
rect 180118 213288 180123 213344
rect 122741 213286 180123 213288
rect 122741 213283 122807 213286
rect 180057 213283 180123 213286
rect 92381 213210 92447 213213
rect 340873 213210 340939 213213
rect 92381 213208 340939 213210
rect 92381 213152 92386 213208
rect 92442 213152 340878 213208
rect 340934 213152 340939 213208
rect 92381 213150 340939 213152
rect 92381 213147 92447 213150
rect 340873 213147 340939 213150
rect 197997 212666 198063 212669
rect 213085 212666 213151 212669
rect 213729 212666 213795 212669
rect 197997 212664 213795 212666
rect 197997 212608 198002 212664
rect 198058 212608 213090 212664
rect 213146 212608 213734 212664
rect 213790 212608 213795 212664
rect 197997 212606 213795 212608
rect 197997 212603 198063 212606
rect 213085 212603 213151 212606
rect 213729 212603 213795 212606
rect 104249 212530 104315 212533
rect 203333 212530 203399 212533
rect 104249 212528 203399 212530
rect 104249 212472 104254 212528
rect 104310 212472 203338 212528
rect 203394 212472 203399 212528
rect 104249 212470 203399 212472
rect 104249 212467 104315 212470
rect 203333 212467 203399 212470
rect 81249 211986 81315 211989
rect 304257 211986 304323 211989
rect 81249 211984 304323 211986
rect 81249 211928 81254 211984
rect 81310 211928 304262 211984
rect 304318 211928 304323 211984
rect 81249 211926 304323 211928
rect 81249 211923 81315 211926
rect 304257 211923 304323 211926
rect 95141 211850 95207 211853
rect 351913 211850 351979 211853
rect 95141 211848 351979 211850
rect 95141 211792 95146 211848
rect 95202 211792 351918 211848
rect 351974 211792 351979 211848
rect 95141 211790 351979 211792
rect 95141 211787 95207 211790
rect 351913 211787 351979 211790
rect 191598 211108 191604 211172
rect 191668 211170 191674 211172
rect 198273 211170 198339 211173
rect 214465 211172 214531 211173
rect 214414 211170 214420 211172
rect 191668 211168 198339 211170
rect 191668 211112 198278 211168
rect 198334 211112 198339 211168
rect 191668 211110 198339 211112
rect 214374 211110 214420 211170
rect 214484 211168 214531 211172
rect 214526 211112 214531 211168
rect 191668 211108 191674 211110
rect 198273 211107 198339 211110
rect 214414 211108 214420 211110
rect 214484 211108 214531 211112
rect 214465 211107 214531 211108
rect 143349 211034 143415 211037
rect 163037 211034 163103 211037
rect 143349 211032 163103 211034
rect 143349 210976 143354 211032
rect 143410 210976 163042 211032
rect 163098 210976 163103 211032
rect 143349 210974 163103 210976
rect 143349 210971 143415 210974
rect 163037 210971 163103 210974
rect 102041 210490 102107 210493
rect 213177 210490 213243 210493
rect 102041 210488 213243 210490
rect 102041 210432 102046 210488
rect 102102 210432 213182 210488
rect 213238 210432 213243 210488
rect 102041 210430 213243 210432
rect 102041 210427 102107 210430
rect 213177 210427 213243 210430
rect 213729 210490 213795 210493
rect 289905 210490 289971 210493
rect 213729 210488 289971 210490
rect 213729 210432 213734 210488
rect 213790 210432 289910 210488
rect 289966 210432 289971 210488
rect 213729 210430 289971 210432
rect 213729 210427 213795 210430
rect 289905 210427 289971 210430
rect 88241 210354 88307 210357
rect 322933 210354 322999 210357
rect 88241 210352 322999 210354
rect 88241 210296 88246 210352
rect 88302 210296 322938 210352
rect 322994 210296 322999 210352
rect 88241 210294 322999 210296
rect 88241 210291 88307 210294
rect 322933 210291 322999 210294
rect 76557 209674 76623 209677
rect 218697 209674 218763 209677
rect 76557 209672 218763 209674
rect 76557 209616 76562 209672
rect 76618 209616 218702 209672
rect 218758 209616 218763 209672
rect 76557 209614 218763 209616
rect 76557 209611 76623 209614
rect 218697 209611 218763 209614
rect 154389 209130 154455 209133
rect 178677 209130 178743 209133
rect 154389 209128 178743 209130
rect 154389 209072 154394 209128
rect 154450 209072 178682 209128
rect 178738 209072 178743 209128
rect 154389 209070 178743 209072
rect 154389 209067 154455 209070
rect 178677 209067 178743 209070
rect 194501 209130 194567 209133
rect 241513 209130 241579 209133
rect 194501 209128 241579 209130
rect 194501 209072 194506 209128
rect 194562 209072 241518 209128
rect 241574 209072 241579 209128
rect 194501 209070 241579 209072
rect 194501 209067 194567 209070
rect 241513 209067 241579 209070
rect 115841 208994 115907 208997
rect 151077 208994 151143 208997
rect 115841 208992 151143 208994
rect 115841 208936 115846 208992
rect 115902 208936 151082 208992
rect 151138 208936 151143 208992
rect 115841 208934 151143 208936
rect 115841 208931 115907 208934
rect 151077 208931 151143 208934
rect 156689 208994 156755 208997
rect 353293 208994 353359 208997
rect 156689 208992 353359 208994
rect 156689 208936 156694 208992
rect 156750 208936 353298 208992
rect 353354 208936 353359 208992
rect 156689 208934 353359 208936
rect 156689 208931 156755 208934
rect 353293 208931 353359 208934
rect 122833 208314 122899 208317
rect 122833 208312 200130 208314
rect 122833 208256 122838 208312
rect 122894 208256 200130 208312
rect 122833 208254 200130 208256
rect 122833 208251 122899 208254
rect 200070 207906 200130 208254
rect 210734 207906 210740 207908
rect 200070 207846 210740 207906
rect 210734 207844 210740 207846
rect 210804 207906 210810 207908
rect 235441 207906 235507 207909
rect 210804 207904 235507 207906
rect 210804 207848 235446 207904
rect 235502 207848 235507 207904
rect 210804 207846 235507 207848
rect 210804 207844 210810 207846
rect 235441 207843 235507 207846
rect 3509 207634 3575 207637
rect 154614 207634 154620 207636
rect 3509 207632 154620 207634
rect 3509 207576 3514 207632
rect 3570 207576 154620 207632
rect 3509 207574 154620 207576
rect 3509 207571 3575 207574
rect 154614 207572 154620 207574
rect 154684 207572 154690 207636
rect 166257 207634 166323 207637
rect 345013 207634 345079 207637
rect 166257 207632 345079 207634
rect 166257 207576 166262 207632
rect 166318 207576 345018 207632
rect 345074 207576 345079 207632
rect 166257 207574 345079 207576
rect 166257 207571 166323 207574
rect 345013 207571 345079 207574
rect 157333 207090 157399 207093
rect 205909 207090 205975 207093
rect 157333 207088 205975 207090
rect 157333 207032 157338 207088
rect 157394 207032 205914 207088
rect 205970 207032 205975 207088
rect 157333 207030 205975 207032
rect 157333 207027 157399 207030
rect 205909 207027 205975 207030
rect 53557 206954 53623 206957
rect 233877 206954 233943 206957
rect 53557 206952 233943 206954
rect 53557 206896 53562 206952
rect 53618 206896 233882 206952
rect 233938 206896 233943 206952
rect 53557 206894 233943 206896
rect 53557 206891 53623 206894
rect 233877 206891 233943 206894
rect 133781 206410 133847 206413
rect 316033 206410 316099 206413
rect 133781 206408 316099 206410
rect 133781 206352 133786 206408
rect 133842 206352 316038 206408
rect 316094 206352 316099 206408
rect 133781 206350 316099 206352
rect 133781 206347 133847 206350
rect 316033 206347 316099 206350
rect 79869 206274 79935 206277
rect 298134 206274 298140 206276
rect 79869 206272 298140 206274
rect 79869 206216 79874 206272
rect 79930 206216 298140 206272
rect 79869 206214 298140 206216
rect 79869 206211 79935 206214
rect 298134 206212 298140 206214
rect 298204 206212 298210 206276
rect 233325 205730 233391 205733
rect 233877 205730 233943 205733
rect 233325 205728 233943 205730
rect 233325 205672 233330 205728
rect 233386 205672 233882 205728
rect 233938 205672 233943 205728
rect 233325 205670 233943 205672
rect 233325 205667 233391 205670
rect 233877 205667 233943 205670
rect 583385 205730 583451 205733
rect 583520 205730 584960 205820
rect 583385 205728 584960 205730
rect 583385 205672 583390 205728
rect 583446 205672 584960 205728
rect 583385 205670 584960 205672
rect 583385 205667 583451 205670
rect 115289 205594 115355 205597
rect 210417 205594 210483 205597
rect 210693 205594 210759 205597
rect 115289 205592 210759 205594
rect 115289 205536 115294 205592
rect 115350 205536 210422 205592
rect 210478 205536 210698 205592
rect 210754 205536 210759 205592
rect 583520 205580 584960 205670
rect 115289 205534 210759 205536
rect 115289 205531 115355 205534
rect 210417 205531 210483 205534
rect 210693 205531 210759 205534
rect 242985 205186 243051 205189
rect 244038 205186 244044 205188
rect 242985 205184 244044 205186
rect 242985 205128 242990 205184
rect 243046 205128 244044 205184
rect 242985 205126 244044 205128
rect 242985 205123 243051 205126
rect 244038 205124 244044 205126
rect 244108 205124 244114 205188
rect 132401 205050 132467 205053
rect 171869 205050 171935 205053
rect 132401 205048 171935 205050
rect 132401 204992 132406 205048
rect 132462 204992 171874 205048
rect 171930 204992 171935 205048
rect 132401 204990 171935 204992
rect 132401 204987 132467 204990
rect 171869 204987 171935 204990
rect 207749 205050 207815 205053
rect 301129 205050 301195 205053
rect 207749 205048 301195 205050
rect 207749 204992 207754 205048
rect 207810 204992 301134 205048
rect 301190 204992 301195 205048
rect 207749 204990 301195 204992
rect 207749 204987 207815 204990
rect 301129 204987 301195 204990
rect 66662 204852 66668 204916
rect 66732 204914 66738 204916
rect 583385 204914 583451 204917
rect 66732 204912 583451 204914
rect 66732 204856 583390 204912
rect 583446 204856 583451 204912
rect 66732 204854 583451 204856
rect 66732 204852 66738 204854
rect 583385 204851 583451 204854
rect 114461 204234 114527 204237
rect 220997 204234 221063 204237
rect 221457 204234 221523 204237
rect 245837 204234 245903 204237
rect 246389 204234 246455 204237
rect 114461 204232 221523 204234
rect 114461 204176 114466 204232
rect 114522 204176 221002 204232
rect 221058 204176 221462 204232
rect 221518 204176 221523 204232
rect 114461 204174 221523 204176
rect 114461 204171 114527 204174
rect 220997 204171 221063 204174
rect 221457 204171 221523 204174
rect 238710 204232 246455 204234
rect 238710 204176 245842 204232
rect 245898 204176 246394 204232
rect 246450 204176 246455 204232
rect 238710 204174 246455 204176
rect 153009 204098 153075 204101
rect 238710 204098 238770 204174
rect 245837 204171 245903 204174
rect 246389 204171 246455 204174
rect 153009 204096 238770 204098
rect 153009 204040 153014 204096
rect 153070 204040 238770 204096
rect 153009 204038 238770 204040
rect 153009 204035 153075 204038
rect 83958 203492 83964 203556
rect 84028 203554 84034 203556
rect 251766 203554 251772 203556
rect 84028 203494 251772 203554
rect 84028 203492 84034 203494
rect 251766 203492 251772 203494
rect 251836 203492 251842 203556
rect 52361 202874 52427 202877
rect 215385 202874 215451 202877
rect 52361 202872 215451 202874
rect 52361 202816 52366 202872
rect 52422 202816 215390 202872
rect 215446 202816 215451 202872
rect 52361 202814 215451 202816
rect 52361 202811 52427 202814
rect 215385 202811 215451 202814
rect 205909 202330 205975 202333
rect 282177 202330 282243 202333
rect 205909 202328 282243 202330
rect 205909 202272 205914 202328
rect 205970 202272 282182 202328
rect 282238 202272 282243 202328
rect 205909 202270 282243 202272
rect 205909 202267 205975 202270
rect 282177 202267 282243 202270
rect 154481 202194 154547 202197
rect 299473 202194 299539 202197
rect 154481 202192 299539 202194
rect 154481 202136 154486 202192
rect 154542 202136 299478 202192
rect 299534 202136 299539 202192
rect 154481 202134 299539 202136
rect 154481 202131 154547 202134
rect 299473 202131 299539 202134
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 119337 201378 119403 201381
rect 166206 201378 166212 201380
rect 119337 201376 166212 201378
rect 119337 201320 119342 201376
rect 119398 201320 166212 201376
rect 119337 201318 166212 201320
rect 119337 201315 119403 201318
rect 166206 201316 166212 201318
rect 166276 201316 166282 201380
rect 129641 200834 129707 200837
rect 288382 200834 288388 200836
rect 129641 200832 288388 200834
rect 129641 200776 129646 200832
rect 129702 200776 288388 200832
rect 129641 200774 288388 200776
rect 129641 200771 129707 200774
rect 288382 200772 288388 200774
rect 288452 200772 288458 200836
rect 67081 200698 67147 200701
rect 583477 200698 583543 200701
rect 67081 200696 583543 200698
rect 67081 200640 67086 200696
rect 67142 200640 583482 200696
rect 583538 200640 583543 200696
rect 67081 200638 583543 200640
rect 67081 200635 67147 200638
rect 583477 200635 583543 200638
rect 239397 199610 239463 199613
rect 252502 199610 252508 199612
rect 239397 199608 252508 199610
rect 239397 199552 239402 199608
rect 239458 199552 252508 199608
rect 239397 199550 252508 199552
rect 239397 199547 239463 199550
rect 252502 199548 252508 199550
rect 252572 199548 252578 199612
rect 118601 199474 118667 199477
rect 202137 199474 202203 199477
rect 118601 199472 202203 199474
rect 118601 199416 118606 199472
rect 118662 199416 202142 199472
rect 202198 199416 202203 199472
rect 118601 199414 202203 199416
rect 118601 199411 118667 199414
rect 202137 199411 202203 199414
rect 213821 199474 213887 199477
rect 240358 199474 240364 199476
rect 213821 199472 240364 199474
rect 213821 199416 213826 199472
rect 213882 199416 240364 199472
rect 213821 199414 240364 199416
rect 213821 199411 213887 199414
rect 240358 199412 240364 199414
rect 240428 199412 240434 199476
rect 61929 199338 61995 199341
rect 311893 199338 311959 199341
rect 61929 199336 311959 199338
rect 61929 199280 61934 199336
rect 61990 199280 311898 199336
rect 311954 199280 311959 199336
rect 61929 199278 311959 199280
rect 61929 199275 61995 199278
rect 311893 199275 311959 199278
rect 135161 198658 135227 198661
rect 204989 198658 205055 198661
rect 135161 198656 205055 198658
rect 135161 198600 135166 198656
rect 135222 198600 204994 198656
rect 205050 198600 205055 198656
rect 135161 198598 205055 198600
rect 135161 198595 135227 198598
rect 204989 198595 205055 198598
rect 104157 198522 104223 198525
rect 157977 198522 158043 198525
rect 104157 198520 158043 198522
rect 104157 198464 104162 198520
rect 104218 198464 157982 198520
rect 158038 198464 158043 198520
rect 104157 198462 158043 198464
rect 104157 198459 104223 198462
rect 157977 198459 158043 198462
rect 222694 198188 222700 198252
rect 222764 198250 222770 198252
rect 241605 198250 241671 198253
rect 222764 198248 241671 198250
rect 222764 198192 241610 198248
rect 241666 198192 241671 198248
rect 222764 198190 241671 198192
rect 222764 198188 222770 198190
rect 241605 198187 241671 198190
rect 173341 198114 173407 198117
rect 289997 198114 290063 198117
rect 173341 198112 290063 198114
rect 173341 198056 173346 198112
rect 173402 198056 290002 198112
rect 290058 198056 290063 198112
rect 173341 198054 290063 198056
rect 173341 198051 173407 198054
rect 289997 198051 290063 198054
rect 73061 197978 73127 197981
rect 358813 197978 358879 197981
rect 73061 197976 358879 197978
rect 73061 197920 73066 197976
rect 73122 197920 358818 197976
rect 358874 197920 358879 197976
rect 73061 197918 358879 197920
rect 73061 197915 73127 197918
rect 358813 197915 358879 197918
rect 77937 197298 78003 197301
rect 220169 197298 220235 197301
rect 77937 197296 220235 197298
rect 77937 197240 77942 197296
rect 77998 197240 220174 197296
rect 220230 197240 220235 197296
rect 77937 197238 220235 197240
rect 77937 197235 78003 197238
rect 220169 197235 220235 197238
rect 224718 196692 224724 196756
rect 224788 196754 224794 196756
rect 232037 196754 232103 196757
rect 224788 196752 232103 196754
rect 224788 196696 232042 196752
rect 232098 196696 232103 196752
rect 224788 196694 232103 196696
rect 224788 196692 224794 196694
rect 232037 196691 232103 196694
rect 140681 196618 140747 196621
rect 332685 196618 332751 196621
rect 140681 196616 332751 196618
rect 140681 196560 140686 196616
rect 140742 196560 332690 196616
rect 332746 196560 332751 196616
rect 140681 196558 332751 196560
rect 140681 196555 140747 196558
rect 332685 196555 332751 196558
rect 225689 196346 225755 196349
rect 228633 196346 228699 196349
rect 225689 196344 228699 196346
rect 225689 196288 225694 196344
rect 225750 196288 228638 196344
rect 228694 196288 228699 196344
rect 225689 196286 228699 196288
rect 225689 196283 225755 196286
rect 228633 196283 228699 196286
rect 130377 195938 130443 195941
rect 248597 195938 248663 195941
rect 130377 195936 248663 195938
rect 130377 195880 130382 195936
rect 130438 195880 248602 195936
rect 248658 195880 248663 195936
rect 130377 195878 248663 195880
rect 130377 195875 130443 195878
rect 248597 195875 248663 195878
rect 107469 195802 107535 195805
rect 158713 195802 158779 195805
rect 107469 195800 158779 195802
rect 107469 195744 107474 195800
rect 107530 195744 158718 195800
rect 158774 195744 158779 195800
rect 107469 195742 158779 195744
rect 107469 195739 107535 195742
rect 158713 195739 158779 195742
rect 151721 195258 151787 195261
rect 316125 195258 316191 195261
rect 151721 195256 316191 195258
rect 151721 195200 151726 195256
rect 151782 195200 316130 195256
rect 316186 195200 316191 195256
rect 151721 195198 316191 195200
rect 151721 195195 151787 195198
rect 316125 195195 316191 195198
rect 168373 194442 168439 194445
rect 169518 194442 169524 194444
rect 168373 194440 169524 194442
rect 168373 194384 168378 194440
rect 168434 194384 169524 194440
rect 168373 194382 169524 194384
rect 168373 194379 168439 194382
rect 169518 194380 169524 194382
rect 169588 194380 169594 194444
rect 156597 194170 156663 194173
rect 233877 194170 233943 194173
rect 156597 194168 233943 194170
rect 156597 194112 156602 194168
rect 156658 194112 233882 194168
rect 233938 194112 233943 194168
rect 156597 194110 233943 194112
rect 156597 194107 156663 194110
rect 233877 194107 233943 194110
rect 65926 193972 65932 194036
rect 65996 194034 66002 194036
rect 180333 194034 180399 194037
rect 65996 194032 180399 194034
rect 65996 193976 180338 194032
rect 180394 193976 180399 194032
rect 65996 193974 180399 193976
rect 65996 193972 66002 193974
rect 180333 193971 180399 193974
rect 266997 194034 267063 194037
rect 283782 194034 283788 194036
rect 266997 194032 283788 194034
rect 266997 193976 267002 194032
rect 267058 193976 283788 194032
rect 266997 193974 283788 193976
rect 266997 193971 267063 193974
rect 283782 193972 283788 193974
rect 283852 193972 283858 194036
rect 107561 193898 107627 193901
rect 287094 193898 287100 193900
rect 107561 193896 287100 193898
rect 107561 193840 107566 193896
rect 107622 193840 287100 193896
rect 107561 193838 287100 193840
rect 107561 193835 107627 193838
rect 287094 193836 287100 193838
rect 287164 193836 287170 193900
rect 111057 193218 111123 193221
rect 212717 193218 212783 193221
rect 111057 193216 212783 193218
rect 111057 193160 111062 193216
rect 111118 193160 212722 193216
rect 212778 193160 212783 193216
rect 111057 193158 212783 193160
rect 111057 193155 111123 193158
rect 212717 193155 212783 193158
rect 218697 192674 218763 192677
rect 280470 192674 280476 192676
rect 218697 192672 280476 192674
rect 218697 192616 218702 192672
rect 218758 192616 280476 192672
rect 218697 192614 280476 192616
rect 218697 192611 218763 192614
rect 280470 192612 280476 192614
rect 280540 192612 280546 192676
rect 85481 192538 85547 192541
rect 255814 192538 255820 192540
rect 85481 192536 255820 192538
rect 85481 192480 85486 192536
rect 85542 192480 255820 192536
rect 85481 192478 255820 192480
rect 85481 192475 85547 192478
rect 255814 192476 255820 192478
rect 255884 192476 255890 192540
rect 580257 192538 580323 192541
rect 583520 192538 584960 192628
rect 580257 192536 584960 192538
rect 580257 192480 580262 192536
rect 580318 192480 584960 192536
rect 580257 192478 584960 192480
rect 580257 192475 580323 192478
rect 583520 192388 584960 192478
rect 97901 191178 97967 191181
rect 249006 191178 249012 191180
rect 97901 191176 249012 191178
rect 97901 191120 97906 191176
rect 97962 191120 249012 191176
rect 97901 191118 249012 191120
rect 97901 191115 97967 191118
rect 249006 191116 249012 191118
rect 249076 191116 249082 191180
rect 133137 191042 133203 191045
rect 318793 191042 318859 191045
rect 133137 191040 318859 191042
rect 133137 190984 133142 191040
rect 133198 190984 318798 191040
rect 318854 190984 318859 191040
rect 133137 190982 318859 190984
rect 133137 190979 133203 190982
rect 318793 190979 318859 190982
rect 148961 189954 149027 189957
rect 181437 189954 181503 189957
rect 148961 189952 181503 189954
rect 148961 189896 148966 189952
rect 149022 189896 181442 189952
rect 181498 189896 181503 189952
rect 148961 189894 181503 189896
rect 148961 189891 149027 189894
rect 181437 189891 181503 189894
rect 195421 189954 195487 189957
rect 300853 189954 300919 189957
rect 195421 189952 300919 189954
rect 195421 189896 195426 189952
rect 195482 189896 300858 189952
rect 300914 189896 300919 189952
rect 195421 189894 300919 189896
rect 195421 189891 195487 189894
rect 300853 189891 300919 189894
rect 89621 189818 89687 189821
rect 196709 189818 196775 189821
rect 89621 189816 196775 189818
rect 89621 189760 89626 189816
rect 89682 189760 196714 189816
rect 196770 189760 196775 189816
rect 89621 189758 196775 189760
rect 89621 189755 89687 189758
rect 196709 189755 196775 189758
rect 161974 189620 161980 189684
rect 162044 189682 162050 189684
rect 335353 189682 335419 189685
rect 162044 189680 335419 189682
rect 162044 189624 335358 189680
rect 335414 189624 335419 189680
rect 162044 189622 335419 189624
rect 162044 189620 162050 189622
rect 335353 189619 335419 189622
rect 221549 189138 221615 189141
rect 248505 189138 248571 189141
rect 221549 189136 248571 189138
rect 221549 189080 221554 189136
rect 221610 189080 248510 189136
rect 248566 189080 248571 189136
rect 221549 189078 248571 189080
rect 221549 189075 221615 189078
rect 248505 189075 248571 189078
rect -960 188866 480 188956
rect 3509 188866 3575 188869
rect -960 188864 3575 188866
rect -960 188808 3514 188864
rect 3570 188808 3575 188864
rect -960 188806 3575 188808
rect -960 188716 480 188806
rect 3509 188803 3575 188806
rect 221222 188532 221228 188596
rect 221292 188594 221298 188596
rect 279141 188594 279207 188597
rect 221292 188592 279207 188594
rect 221292 188536 279146 188592
rect 279202 188536 279207 188592
rect 221292 188534 279207 188536
rect 221292 188532 221298 188534
rect 279141 188531 279207 188534
rect 160829 188458 160895 188461
rect 180241 188458 180307 188461
rect 160829 188456 180307 188458
rect 160829 188400 160834 188456
rect 160890 188400 180246 188456
rect 180302 188400 180307 188456
rect 160829 188398 180307 188400
rect 160829 188395 160895 188398
rect 180241 188395 180307 188398
rect 184749 188458 184815 188461
rect 242934 188458 242940 188460
rect 184749 188456 242940 188458
rect 184749 188400 184754 188456
rect 184810 188400 242940 188456
rect 184749 188398 242940 188400
rect 184749 188395 184815 188398
rect 242934 188396 242940 188398
rect 243004 188396 243010 188460
rect 99281 188322 99347 188325
rect 305085 188322 305151 188325
rect 99281 188320 305151 188322
rect 99281 188264 99286 188320
rect 99342 188264 305090 188320
rect 305146 188264 305151 188320
rect 99281 188262 305151 188264
rect 99281 188259 99347 188262
rect 305085 188259 305151 188262
rect 180333 187642 180399 187645
rect 209773 187642 209839 187645
rect 211061 187642 211127 187645
rect 180333 187640 211127 187642
rect 180333 187584 180338 187640
rect 180394 187584 209778 187640
rect 209834 187584 211066 187640
rect 211122 187584 211127 187640
rect 180333 187582 211127 187584
rect 180333 187579 180399 187582
rect 209773 187579 209839 187582
rect 211061 187579 211127 187582
rect 203517 187234 203583 187237
rect 238845 187234 238911 187237
rect 203517 187232 238911 187234
rect 203517 187176 203522 187232
rect 203578 187176 238850 187232
rect 238906 187176 238911 187232
rect 203517 187174 238911 187176
rect 203517 187171 203583 187174
rect 238845 187171 238911 187174
rect 151077 187098 151143 187101
rect 293953 187098 294019 187101
rect 151077 187096 294019 187098
rect 151077 187040 151082 187096
rect 151138 187040 293958 187096
rect 294014 187040 294019 187096
rect 151077 187038 294019 187040
rect 151077 187035 151143 187038
rect 293953 187035 294019 187038
rect 153101 186962 153167 186965
rect 167637 186962 167703 186965
rect 153101 186960 167703 186962
rect 153101 186904 153106 186960
rect 153162 186904 167642 186960
rect 167698 186904 167703 186960
rect 153101 186902 167703 186904
rect 153101 186899 153167 186902
rect 167637 186899 167703 186902
rect 211061 186962 211127 186965
rect 580257 186962 580323 186965
rect 211061 186960 580323 186962
rect 211061 186904 211066 186960
rect 211122 186904 580262 186960
rect 580318 186904 580323 186960
rect 211061 186902 580323 186904
rect 211061 186899 211127 186902
rect 580257 186899 580323 186902
rect 240726 186356 240732 186420
rect 240796 186418 240802 186420
rect 242157 186418 242223 186421
rect 240796 186416 242223 186418
rect 240796 186360 242162 186416
rect 242218 186360 242223 186416
rect 240796 186358 242223 186360
rect 240796 186356 240802 186358
rect 242157 186355 242223 186358
rect 91001 185738 91067 185741
rect 246246 185738 246252 185740
rect 91001 185736 246252 185738
rect 91001 185680 91006 185736
rect 91062 185680 246252 185736
rect 91001 185678 246252 185680
rect 91001 185675 91067 185678
rect 246246 185676 246252 185678
rect 246316 185676 246322 185740
rect 271137 185738 271203 185741
rect 291326 185738 291332 185740
rect 271137 185736 291332 185738
rect 271137 185680 271142 185736
rect 271198 185680 291332 185736
rect 271137 185678 291332 185680
rect 271137 185675 271203 185678
rect 291326 185676 291332 185678
rect 291396 185676 291402 185740
rect 168966 185540 168972 185604
rect 169036 185602 169042 185604
rect 329833 185602 329899 185605
rect 169036 185600 329899 185602
rect 169036 185544 329838 185600
rect 329894 185544 329899 185600
rect 169036 185542 329899 185544
rect 169036 185540 169042 185542
rect 329833 185539 329899 185542
rect 193029 184378 193095 184381
rect 241697 184378 241763 184381
rect 193029 184376 241763 184378
rect 193029 184320 193034 184376
rect 193090 184320 241702 184376
rect 241758 184320 241763 184376
rect 193029 184318 241763 184320
rect 193029 184315 193095 184318
rect 241697 184315 241763 184318
rect 145414 184180 145420 184244
rect 145484 184242 145490 184244
rect 197997 184242 198063 184245
rect 145484 184240 198063 184242
rect 145484 184184 198002 184240
rect 198058 184184 198063 184240
rect 145484 184182 198063 184184
rect 145484 184180 145490 184182
rect 197997 184179 198063 184182
rect 210417 184242 210483 184245
rect 288566 184242 288572 184244
rect 210417 184240 288572 184242
rect 210417 184184 210422 184240
rect 210478 184184 288572 184240
rect 210417 184182 288572 184184
rect 210417 184179 210483 184182
rect 288566 184180 288572 184182
rect 288636 184180 288642 184244
rect 100661 183698 100727 183701
rect 180333 183698 180399 183701
rect 100661 183696 180399 183698
rect 100661 183640 100666 183696
rect 100722 183640 180338 183696
rect 180394 183640 180399 183696
rect 100661 183638 180399 183640
rect 100661 183635 100727 183638
rect 180333 183635 180399 183638
rect 196801 183154 196867 183157
rect 237598 183154 237604 183156
rect 196801 183152 237604 183154
rect 196801 183096 196806 183152
rect 196862 183096 237604 183152
rect 196801 183094 237604 183096
rect 196801 183091 196867 183094
rect 237598 183092 237604 183094
rect 237668 183092 237674 183156
rect 226926 182956 226932 183020
rect 226996 183018 227002 183020
rect 233417 183018 233483 183021
rect 226996 183016 233483 183018
rect 226996 182960 233422 183016
rect 233478 182960 233483 183016
rect 226996 182958 233483 182960
rect 226996 182956 227002 182958
rect 233417 182955 233483 182958
rect 233877 183018 233943 183021
rect 284518 183018 284524 183020
rect 233877 183016 284524 183018
rect 233877 182960 233882 183016
rect 233938 182960 284524 183016
rect 233877 182958 284524 182960
rect 233877 182955 233943 182958
rect 284518 182956 284524 182958
rect 284588 182956 284594 183020
rect 160737 182882 160803 182885
rect 285806 182882 285812 182884
rect 160737 182880 285812 182882
rect 160737 182824 160742 182880
rect 160798 182824 285812 182880
rect 160737 182822 285812 182824
rect 160737 182819 160803 182822
rect 285806 182820 285812 182822
rect 285876 182820 285882 182884
rect 119521 182338 119587 182341
rect 169109 182338 169175 182341
rect 119521 182336 169175 182338
rect 119521 182280 119526 182336
rect 119582 182280 169114 182336
rect 169170 182280 169175 182336
rect 119521 182278 169175 182280
rect 119521 182275 119587 182278
rect 169109 182275 169175 182278
rect 98913 182202 98979 182205
rect 178861 182202 178927 182205
rect 98913 182200 178927 182202
rect 98913 182144 98918 182200
rect 98974 182144 178866 182200
rect 178922 182144 178927 182200
rect 98913 182142 178927 182144
rect 98913 182139 98979 182142
rect 178861 182139 178927 182142
rect 231761 182066 231827 182069
rect 233182 182066 233188 182068
rect 231761 182064 233188 182066
rect 231761 182008 231766 182064
rect 231822 182008 233188 182064
rect 231761 182006 233188 182008
rect 231761 182003 231827 182006
rect 233182 182004 233188 182006
rect 233252 182004 233258 182068
rect 226977 181658 227043 181661
rect 236177 181658 236243 181661
rect 226977 181656 236243 181658
rect 226977 181600 226982 181656
rect 227038 181600 236182 181656
rect 236238 181600 236243 181656
rect 226977 181598 236243 181600
rect 226977 181595 227043 181598
rect 236177 181595 236243 181598
rect 196893 181522 196959 181525
rect 230606 181522 230612 181524
rect 196893 181520 230612 181522
rect 196893 181464 196898 181520
rect 196954 181464 230612 181520
rect 196893 181462 230612 181464
rect 196893 181459 196959 181462
rect 230606 181460 230612 181462
rect 230676 181460 230682 181524
rect 269757 181522 269823 181525
rect 281574 181522 281580 181524
rect 269757 181520 281580 181522
rect 269757 181464 269762 181520
rect 269818 181464 281580 181520
rect 269757 181462 281580 181464
rect 269757 181459 269823 181462
rect 281574 181460 281580 181462
rect 281644 181460 281650 181524
rect 166349 181386 166415 181389
rect 229277 181386 229343 181389
rect 166349 181384 229343 181386
rect 166349 181328 166354 181384
rect 166410 181328 229282 181384
rect 229338 181328 229343 181384
rect 166349 181326 229343 181328
rect 166349 181323 166415 181326
rect 229277 181323 229343 181326
rect 235349 181386 235415 181389
rect 281717 181386 281783 181389
rect 235349 181384 281783 181386
rect 235349 181328 235354 181384
rect 235410 181328 281722 181384
rect 281778 181328 281783 181384
rect 235349 181326 281783 181328
rect 235349 181323 235415 181326
rect 281717 181323 281783 181326
rect 100753 180978 100819 180981
rect 166533 180978 166599 180981
rect 100753 180976 166599 180978
rect 100753 180920 100758 180976
rect 100814 180920 166538 180976
rect 166594 180920 166599 180976
rect 100753 180918 166599 180920
rect 100753 180915 100819 180918
rect 166533 180915 166599 180918
rect 115841 180842 115907 180845
rect 191281 180842 191347 180845
rect 115841 180840 191347 180842
rect 115841 180784 115846 180840
rect 115902 180784 191286 180840
rect 191342 180784 191347 180840
rect 115841 180782 191347 180784
rect 115841 180779 115907 180782
rect 191281 180779 191347 180782
rect 226333 180706 226399 180709
rect 229870 180706 229876 180708
rect 226333 180704 229876 180706
rect 226333 180648 226338 180704
rect 226394 180648 229876 180704
rect 226333 180646 229876 180648
rect 226333 180643 226399 180646
rect 229870 180644 229876 180646
rect 229940 180644 229946 180708
rect 221457 180162 221523 180165
rect 283097 180162 283163 180165
rect 221457 180160 283163 180162
rect 221457 180104 221462 180160
rect 221518 180104 283102 180160
rect 283158 180104 283163 180160
rect 221457 180102 283163 180104
rect 221457 180099 221523 180102
rect 283097 180099 283163 180102
rect 160001 180026 160067 180029
rect 233877 180026 233943 180029
rect 160001 180024 233943 180026
rect 160001 179968 160006 180024
rect 160062 179968 233882 180024
rect 233938 179968 233943 180024
rect 160001 179966 233943 179968
rect 160001 179963 160067 179966
rect 233877 179963 233943 179966
rect 110229 179482 110295 179485
rect 185669 179482 185735 179485
rect 110229 179480 185735 179482
rect 110229 179424 110234 179480
rect 110290 179424 185674 179480
rect 185730 179424 185735 179480
rect 110229 179422 185735 179424
rect 110229 179419 110295 179422
rect 185669 179419 185735 179422
rect 278037 179482 278103 179485
rect 280429 179482 280495 179485
rect 278037 179480 280495 179482
rect 278037 179424 278042 179480
rect 278098 179424 280434 179480
rect 280490 179424 280495 179480
rect 278037 179422 280495 179424
rect 278037 179419 278103 179422
rect 280429 179419 280495 179422
rect 181621 179346 181687 179349
rect 221549 179346 221615 179349
rect 181621 179344 221615 179346
rect 181621 179288 181626 179344
rect 181682 179288 221554 179344
rect 221610 179288 221615 179344
rect 181621 179286 221615 179288
rect 181621 179283 181687 179286
rect 221549 179283 221615 179286
rect 580165 179210 580231 179213
rect 583520 179210 584960 179300
rect 580165 179208 584960 179210
rect 580165 179152 580170 179208
rect 580226 179152 584960 179208
rect 580165 179150 584960 179152
rect 580165 179147 580231 179150
rect 274582 179012 274588 179076
rect 274652 179074 274658 179076
rect 279417 179074 279483 179077
rect 274652 179072 279483 179074
rect 274652 179016 279422 179072
rect 279478 179016 279483 179072
rect 583520 179060 584960 179150
rect 274652 179014 279483 179016
rect 274652 179012 274658 179014
rect 279417 179011 279483 179014
rect 276749 178938 276815 178941
rect 288709 178938 288775 178941
rect 276749 178936 288775 178938
rect 276749 178880 276754 178936
rect 276810 178880 288714 178936
rect 288770 178880 288775 178936
rect 276749 178878 288775 178880
rect 276749 178875 276815 178878
rect 288709 178875 288775 178878
rect 247677 178802 247743 178805
rect 292757 178802 292823 178805
rect 247677 178800 292823 178802
rect 247677 178744 247682 178800
rect 247738 178744 292762 178800
rect 292818 178744 292823 178800
rect 247677 178742 292823 178744
rect 247677 178739 247743 178742
rect 292757 178739 292823 178742
rect 183461 178666 183527 178669
rect 226333 178666 226399 178669
rect 278814 178666 278820 178668
rect 183461 178664 219450 178666
rect 183461 178608 183466 178664
rect 183522 178608 219450 178664
rect 183461 178606 219450 178608
rect 183461 178603 183527 178606
rect 219390 178530 219450 178606
rect 226333 178664 278820 178666
rect 226333 178608 226338 178664
rect 226394 178608 278820 178664
rect 226333 178606 278820 178608
rect 226333 178603 226399 178606
rect 278814 178604 278820 178606
rect 278884 178604 278890 178668
rect 226333 178530 226399 178533
rect 219390 178528 226399 178530
rect 219390 178472 226338 178528
rect 226394 178472 226399 178528
rect 219390 178470 226399 178472
rect 226333 178467 226399 178470
rect 231710 178332 231716 178396
rect 231780 178394 231786 178396
rect 236085 178394 236151 178397
rect 231780 178392 236151 178394
rect 231780 178336 236090 178392
rect 236146 178336 236151 178392
rect 231780 178334 236151 178336
rect 231780 178332 231786 178334
rect 236085 178331 236151 178334
rect 113214 178196 113220 178260
rect 113284 178258 113290 178260
rect 177481 178258 177547 178261
rect 113284 178256 177547 178258
rect 113284 178200 177486 178256
rect 177542 178200 177547 178256
rect 113284 178198 177547 178200
rect 113284 178196 113290 178198
rect 177481 178195 177547 178198
rect 223481 178258 223547 178261
rect 231761 178258 231827 178261
rect 223481 178256 231827 178258
rect 223481 178200 223486 178256
rect 223542 178200 231766 178256
rect 231822 178200 231827 178256
rect 223481 178198 231827 178200
rect 223481 178195 223547 178198
rect 231761 178195 231827 178198
rect 166206 178122 166212 178124
rect 97030 178062 166212 178122
rect 97030 177988 97090 178062
rect 166206 178060 166212 178062
rect 166276 178060 166282 178124
rect 215293 178122 215359 178125
rect 244549 178122 244615 178125
rect 215293 178120 244615 178122
rect 215293 178064 215298 178120
rect 215354 178064 244554 178120
rect 244610 178064 244615 178120
rect 215293 178062 244615 178064
rect 215293 178059 215359 178062
rect 244549 178059 244615 178062
rect 97022 177924 97028 177988
rect 97092 177924 97098 177988
rect 222837 177986 222903 177989
rect 229369 177986 229435 177989
rect 222837 177984 229435 177986
rect 222837 177928 222842 177984
rect 222898 177928 229374 177984
rect 229430 177928 229435 177984
rect 222837 177926 229435 177928
rect 222837 177923 222903 177926
rect 229369 177923 229435 177926
rect 98310 177516 98316 177580
rect 98380 177578 98386 177580
rect 98913 177578 98979 177581
rect 100753 177580 100819 177581
rect 100702 177578 100708 177580
rect 98380 177576 98979 177578
rect 98380 177520 98918 177576
rect 98974 177520 98979 177576
rect 98380 177518 98979 177520
rect 100662 177518 100708 177578
rect 100772 177576 100819 177580
rect 100814 177520 100819 177576
rect 98380 177516 98386 177518
rect 98913 177515 98979 177518
rect 100702 177516 100708 177518
rect 100772 177516 100819 177520
rect 105670 177516 105676 177580
rect 105740 177578 105746 177580
rect 106181 177578 106247 177581
rect 105740 177576 106247 177578
rect 105740 177520 106186 177576
rect 106242 177520 106247 177576
rect 105740 177518 106247 177520
rect 105740 177516 105746 177518
rect 100753 177515 100819 177516
rect 106181 177515 106247 177518
rect 108062 177516 108068 177580
rect 108132 177578 108138 177580
rect 108941 177578 109007 177581
rect 115841 177580 115907 177581
rect 119521 177580 119587 177581
rect 115790 177578 115796 177580
rect 108132 177576 109007 177578
rect 108132 177520 108946 177576
rect 109002 177520 109007 177576
rect 108132 177518 109007 177520
rect 115750 177518 115796 177578
rect 115860 177576 115907 177580
rect 119470 177578 119476 177580
rect 115902 177520 115907 177576
rect 108132 177516 108138 177518
rect 108941 177515 109007 177518
rect 115790 177516 115796 177518
rect 115860 177516 115907 177520
rect 119430 177518 119476 177578
rect 119540 177576 119587 177580
rect 119582 177520 119587 177576
rect 119470 177516 119476 177518
rect 119540 177516 119587 177520
rect 121862 177516 121868 177580
rect 121932 177578 121938 177580
rect 122741 177578 122807 177581
rect 121932 177576 122807 177578
rect 121932 177520 122746 177576
rect 122802 177520 122807 177576
rect 121932 177518 122807 177520
rect 121932 177516 121938 177518
rect 115841 177515 115907 177516
rect 119521 177515 119587 177516
rect 122741 177515 122807 177518
rect 123150 177516 123156 177580
rect 123220 177578 123226 177580
rect 124121 177578 124187 177581
rect 123220 177576 124187 177578
rect 123220 177520 124126 177576
rect 124182 177520 124187 177576
rect 123220 177518 124187 177520
rect 123220 177516 123226 177518
rect 124121 177515 124187 177518
rect 125726 177516 125732 177580
rect 125796 177578 125802 177580
rect 125961 177578 126027 177581
rect 125796 177576 126027 177578
rect 125796 177520 125966 177576
rect 126022 177520 126027 177576
rect 125796 177518 126027 177520
rect 125796 177516 125802 177518
rect 125961 177515 126027 177518
rect 127014 177516 127020 177580
rect 127084 177578 127090 177580
rect 128261 177578 128327 177581
rect 127084 177576 128327 177578
rect 127084 177520 128266 177576
rect 128322 177520 128327 177576
rect 127084 177518 128327 177520
rect 127084 177516 127090 177518
rect 128261 177515 128327 177518
rect 129406 177516 129412 177580
rect 129476 177578 129482 177580
rect 129641 177578 129707 177581
rect 132401 177580 132467 177581
rect 133137 177580 133203 177581
rect 132350 177578 132356 177580
rect 129476 177576 129707 177578
rect 129476 177520 129646 177576
rect 129702 177520 129707 177576
rect 129476 177518 129707 177520
rect 132310 177518 132356 177578
rect 132420 177576 132467 177580
rect 133086 177578 133092 177580
rect 132462 177520 132467 177576
rect 129476 177516 129482 177518
rect 129641 177515 129707 177518
rect 132350 177516 132356 177518
rect 132420 177516 132467 177520
rect 133046 177518 133092 177578
rect 133156 177576 133203 177580
rect 133198 177520 133203 177576
rect 133086 177516 133092 177518
rect 133156 177516 133203 177520
rect 134374 177516 134380 177580
rect 134444 177578 134450 177580
rect 135161 177578 135227 177581
rect 148225 177580 148291 177581
rect 148174 177578 148180 177580
rect 134444 177576 135227 177578
rect 134444 177520 135166 177576
rect 135222 177520 135227 177576
rect 134444 177518 135227 177520
rect 148134 177518 148180 177578
rect 148244 177576 148291 177580
rect 148286 177520 148291 177576
rect 134444 177516 134450 177518
rect 132401 177515 132467 177516
rect 133137 177515 133203 177516
rect 135161 177515 135227 177518
rect 148174 177516 148180 177518
rect 148244 177516 148291 177520
rect 148225 177515 148291 177516
rect 195329 177442 195395 177445
rect 230422 177442 230428 177444
rect 195329 177440 230428 177442
rect 195329 177384 195334 177440
rect 195390 177384 230428 177440
rect 195329 177382 230428 177384
rect 195329 177379 195395 177382
rect 230422 177380 230428 177382
rect 230492 177380 230498 177444
rect 272517 177442 272583 177445
rect 287278 177442 287284 177444
rect 272517 177440 287284 177442
rect 272517 177384 272522 177440
rect 272578 177384 287284 177440
rect 272517 177382 287284 177384
rect 272517 177379 272583 177382
rect 287278 177380 287284 177382
rect 287348 177380 287354 177444
rect 104566 177244 104572 177308
rect 104636 177306 104642 177308
rect 223389 177306 223455 177309
rect 298369 177306 298435 177309
rect 104636 177246 113190 177306
rect 104636 177244 104642 177246
rect 106958 177108 106964 177172
rect 107028 177170 107034 177172
rect 113130 177170 113190 177246
rect 223389 177304 298435 177306
rect 223389 177248 223394 177304
rect 223450 177248 298374 177304
rect 298430 177248 298435 177304
rect 223389 177246 298435 177248
rect 223389 177243 223455 177246
rect 298369 177243 298435 177246
rect 195513 177170 195579 177173
rect 107028 177110 112546 177170
rect 113130 177168 195579 177170
rect 113130 177112 195518 177168
rect 195574 177112 195579 177168
rect 113130 177110 195579 177112
rect 107028 177108 107034 177110
rect 109534 176972 109540 177036
rect 109604 177034 109610 177036
rect 110229 177034 110295 177037
rect 109604 177032 110295 177034
rect 109604 176976 110234 177032
rect 110290 176976 110295 177032
rect 109604 176974 110295 176976
rect 109604 176972 109610 176974
rect 110229 176971 110295 176974
rect 112110 176972 112116 177036
rect 112180 177034 112186 177036
rect 112253 177034 112319 177037
rect 112180 177032 112319 177034
rect 112180 176976 112258 177032
rect 112314 176976 112319 177032
rect 112180 176974 112319 176976
rect 112486 177034 112546 177110
rect 195513 177107 195579 177110
rect 169201 177034 169267 177037
rect 112486 177032 169267 177034
rect 112486 176976 169206 177032
rect 169262 176976 169267 177032
rect 112486 176974 169267 176976
rect 112180 176972 112186 176974
rect 112253 176971 112319 176974
rect 169201 176971 169267 176974
rect 278773 177034 278839 177037
rect 279366 177034 279372 177036
rect 278773 177032 279372 177034
rect 278773 176976 278778 177032
rect 278834 176976 279372 177032
rect 278773 176974 279372 176976
rect 278773 176971 278839 176974
rect 279366 176972 279372 176974
rect 279436 176972 279442 177036
rect 101990 176836 101996 176900
rect 102060 176898 102066 176900
rect 181529 176898 181595 176901
rect 229185 176900 229251 176901
rect 229134 176898 229140 176900
rect 102060 176896 181595 176898
rect 102060 176840 181534 176896
rect 181590 176840 181595 176896
rect 102060 176838 181595 176840
rect 229094 176838 229140 176898
rect 229204 176896 229251 176900
rect 229246 176840 229251 176896
rect 102060 176836 102066 176838
rect 181529 176835 181595 176838
rect 229134 176836 229140 176838
rect 229204 176836 229251 176840
rect 229185 176835 229251 176836
rect 100661 176762 100727 176765
rect 103421 176762 103487 176765
rect 116945 176764 117011 176765
rect 116894 176762 116900 176764
rect 99422 176760 100727 176762
rect 99422 176704 100666 176760
rect 100722 176704 100727 176760
rect 99422 176702 100727 176704
rect 99422 176492 99482 176702
rect 100661 176699 100727 176702
rect 103286 176760 103487 176762
rect 103286 176704 103426 176760
rect 103482 176704 103487 176760
rect 103286 176702 103487 176704
rect 116854 176702 116900 176762
rect 116964 176760 117011 176764
rect 117006 176704 117011 176760
rect 103286 176492 103346 176702
rect 103421 176699 103487 176702
rect 116894 176700 116900 176702
rect 116964 176700 117011 176704
rect 120758 176700 120764 176764
rect 120828 176762 120834 176764
rect 120993 176762 121059 176765
rect 124489 176764 124555 176765
rect 124438 176762 124444 176764
rect 120828 176760 121059 176762
rect 120828 176704 120998 176760
rect 121054 176704 121059 176760
rect 120828 176702 121059 176704
rect 124398 176702 124444 176762
rect 124508 176760 124555 176764
rect 128169 176762 128235 176765
rect 136081 176764 136147 176765
rect 136030 176762 136036 176764
rect 124550 176704 124555 176760
rect 120828 176700 120834 176702
rect 116945 176699 117011 176700
rect 120993 176699 121059 176702
rect 124438 176700 124444 176702
rect 124508 176700 124555 176704
rect 124489 176699 124555 176700
rect 128126 176760 128235 176762
rect 128126 176704 128174 176760
rect 128230 176704 128235 176760
rect 128126 176699 128235 176704
rect 135990 176702 136036 176762
rect 136100 176760 136147 176764
rect 136142 176704 136147 176760
rect 136030 176700 136036 176702
rect 136100 176700 136147 176704
rect 158846 176700 158852 176764
rect 158916 176762 158922 176764
rect 158989 176762 159055 176765
rect 158916 176760 159055 176762
rect 158916 176704 158994 176760
rect 159050 176704 159055 176760
rect 158916 176702 159055 176704
rect 158916 176700 158922 176702
rect 136081 176699 136147 176700
rect 158989 176699 159055 176702
rect 227805 176762 227871 176765
rect 279233 176762 279299 176765
rect 227805 176760 279299 176762
rect 227805 176704 227810 176760
rect 227866 176704 279238 176760
rect 279294 176704 279299 176760
rect 227805 176702 279299 176704
rect 227805 176699 227871 176702
rect 279233 176699 279299 176702
rect 128126 176492 128186 176699
rect 226190 176564 226196 176628
rect 226260 176626 226266 176628
rect 229185 176626 229251 176629
rect 226260 176624 229251 176626
rect 226260 176568 229190 176624
rect 229246 176568 229251 176624
rect 226260 176566 229251 176568
rect 226260 176564 226266 176566
rect 229185 176563 229251 176566
rect 230606 176564 230612 176628
rect 230676 176626 230682 176628
rect 231485 176626 231551 176629
rect 254025 176626 254091 176629
rect 230676 176624 254091 176626
rect 230676 176568 231490 176624
rect 231546 176568 254030 176624
rect 254086 176568 254091 176624
rect 230676 176566 254091 176568
rect 230676 176564 230682 176566
rect 231485 176563 231551 176566
rect 254025 176563 254091 176566
rect 99414 176428 99420 176492
rect 99484 176428 99490 176492
rect 103278 176428 103284 176492
rect 103348 176428 103354 176492
rect 128118 176428 128124 176492
rect 128188 176428 128194 176492
rect 227713 176218 227779 176221
rect 227713 176216 228282 176218
rect 227713 176160 227718 176216
rect 227774 176160 228282 176216
rect 227713 176158 228282 176160
rect 227713 176155 227779 176158
rect -960 175796 480 176036
rect 118366 175884 118372 175948
rect 118436 175946 118442 175948
rect 214925 175946 214991 175949
rect 223665 175948 223731 175949
rect 223614 175946 223620 175948
rect 118436 175944 214991 175946
rect 118436 175888 214930 175944
rect 214986 175888 214991 175944
rect 118436 175886 214991 175888
rect 223574 175886 223620 175946
rect 223684 175944 223731 175948
rect 223726 175888 223731 175944
rect 118436 175884 118442 175886
rect 214925 175883 214991 175886
rect 223614 175884 223620 175886
rect 223684 175884 223731 175888
rect 223665 175883 223731 175884
rect 130745 175676 130811 175677
rect 130694 175674 130700 175676
rect 130654 175614 130700 175674
rect 130764 175672 130811 175676
rect 130806 175616 130811 175672
rect 130694 175612 130700 175614
rect 130764 175612 130811 175616
rect 130745 175611 130811 175612
rect 213913 175674 213979 175677
rect 213913 175672 217028 175674
rect 213913 175616 213918 175672
rect 213974 175616 217028 175672
rect 228222 175644 228282 176158
rect 228357 175946 228423 175949
rect 228541 175946 228607 175949
rect 232078 175946 232084 175948
rect 228357 175944 228466 175946
rect 228357 175888 228362 175944
rect 228418 175888 228466 175944
rect 228357 175883 228466 175888
rect 228541 175944 232084 175946
rect 228541 175888 228546 175944
rect 228602 175888 232084 175944
rect 228541 175886 232084 175888
rect 228541 175883 228607 175886
rect 232078 175884 232084 175886
rect 232148 175884 232154 175948
rect 228406 175810 228466 175883
rect 234654 175810 234660 175812
rect 228406 175750 234660 175810
rect 234654 175748 234660 175750
rect 234724 175748 234730 175812
rect 264973 175674 265039 175677
rect 264973 175672 268180 175674
rect 213913 175614 217028 175616
rect 264973 175616 264978 175672
rect 265034 175616 268180 175672
rect 264973 175614 268180 175616
rect 213913 175611 213979 175614
rect 264973 175611 265039 175614
rect 114318 175476 114324 175540
rect 114388 175538 114394 175540
rect 166349 175538 166415 175541
rect 114388 175536 166415 175538
rect 114388 175480 166354 175536
rect 166410 175480 166415 175536
rect 114388 175478 166415 175480
rect 114388 175476 114394 175478
rect 166349 175475 166415 175478
rect 110638 175340 110644 175404
rect 110708 175402 110714 175404
rect 171961 175402 172027 175405
rect 110708 175400 172027 175402
rect 110708 175344 171966 175400
rect 172022 175344 172027 175400
rect 110708 175342 172027 175344
rect 110708 175340 110714 175342
rect 171961 175339 172027 175342
rect 279374 175269 279434 175508
rect 164877 175266 164943 175269
rect 169293 175266 169359 175269
rect 164877 175264 169359 175266
rect 164877 175208 164882 175264
rect 164938 175208 169298 175264
rect 169354 175208 169359 175264
rect 164877 175206 169359 175208
rect 164877 175203 164943 175206
rect 169293 175203 169359 175206
rect 178769 175266 178835 175269
rect 214097 175266 214163 175269
rect 231761 175266 231827 175269
rect 178769 175264 214163 175266
rect 178769 175208 178774 175264
rect 178830 175208 214102 175264
rect 214158 175208 214163 175264
rect 178769 175206 214163 175208
rect 228988 175264 231827 175266
rect 228988 175208 231766 175264
rect 231822 175208 231827 175264
rect 228988 175206 231827 175208
rect 178769 175203 178835 175206
rect 214097 175203 214163 175206
rect 231761 175203 231827 175206
rect 265065 175266 265131 175269
rect 265065 175264 268180 175266
rect 265065 175208 265070 175264
rect 265126 175208 268180 175264
rect 265065 175206 268180 175208
rect 279325 175264 279434 175269
rect 279325 175208 279330 175264
rect 279386 175208 279434 175264
rect 279325 175206 279434 175208
rect 265065 175203 265131 175206
rect 279325 175203 279391 175206
rect 213913 174994 213979 174997
rect 213913 174992 217028 174994
rect 213913 174936 213918 174992
rect 213974 174936 217028 174992
rect 213913 174934 217028 174936
rect 213913 174931 213979 174934
rect 264973 174858 265039 174861
rect 264973 174856 268180 174858
rect 264973 174800 264978 174856
rect 265034 174800 268180 174856
rect 264973 174798 268180 174800
rect 264973 174795 265039 174798
rect 231485 174722 231551 174725
rect 280337 174722 280403 174725
rect 228988 174720 231551 174722
rect 228988 174664 231490 174720
rect 231546 174664 231551 174720
rect 228988 174662 231551 174664
rect 279956 174720 280403 174722
rect 279956 174664 280342 174720
rect 280398 174664 280403 174720
rect 279956 174662 280403 174664
rect 231485 174659 231551 174662
rect 280337 174659 280403 174662
rect 229277 174586 229343 174589
rect 232037 174586 232103 174589
rect 229277 174584 232103 174586
rect 229277 174528 229282 174584
rect 229338 174528 232042 174584
rect 232098 174528 232103 174584
rect 229277 174526 232103 174528
rect 229277 174523 229343 174526
rect 232037 174523 232103 174526
rect 260097 174450 260163 174453
rect 279417 174450 279483 174453
rect 260097 174448 268180 174450
rect 260097 174392 260102 174448
rect 260158 174392 268180 174448
rect 260097 174390 268180 174392
rect 279374 174448 279483 174450
rect 279374 174392 279422 174448
rect 279478 174392 279483 174448
rect 260097 174387 260163 174390
rect 279374 174387 279483 174392
rect 214005 174314 214071 174317
rect 256693 174314 256759 174317
rect 214005 174312 217028 174314
rect 214005 174256 214010 174312
rect 214066 174256 217028 174312
rect 214005 174254 217028 174256
rect 228988 174312 256759 174314
rect 228988 174256 256698 174312
rect 256754 174256 256759 174312
rect 228988 174254 256759 174256
rect 214005 174251 214071 174254
rect 256693 174251 256759 174254
rect 238293 174042 238359 174045
rect 238293 174040 268180 174042
rect 238293 173984 238298 174040
rect 238354 173984 268180 174040
rect 279374 174012 279434 174387
rect 238293 173982 268180 173984
rect 238293 173979 238359 173982
rect 229870 173844 229876 173908
rect 229940 173906 229946 173908
rect 230841 173906 230907 173909
rect 229940 173904 230907 173906
rect 229940 173848 230846 173904
rect 230902 173848 230907 173904
rect 229940 173846 230907 173848
rect 229940 173844 229946 173846
rect 230841 173843 230907 173846
rect 230749 173770 230815 173773
rect 228988 173768 230815 173770
rect 228988 173712 230754 173768
rect 230810 173712 230815 173768
rect 228988 173710 230815 173712
rect 230749 173707 230815 173710
rect 279366 173708 279372 173772
rect 279436 173708 279442 173772
rect 213913 173634 213979 173637
rect 265065 173634 265131 173637
rect 213913 173632 217028 173634
rect 213913 173576 213918 173632
rect 213974 173576 217028 173632
rect 213913 173574 217028 173576
rect 265065 173632 268180 173634
rect 265065 173576 265070 173632
rect 265126 173576 268180 173632
rect 265065 173574 268180 173576
rect 213913 173571 213979 173574
rect 265065 173571 265131 173574
rect 229185 173362 229251 173365
rect 228988 173360 229251 173362
rect 228988 173304 229190 173360
rect 229246 173304 229251 173360
rect 228988 173302 229251 173304
rect 229185 173299 229251 173302
rect 279374 173196 279434 173708
rect 214005 172954 214071 172957
rect 214005 172952 217028 172954
rect 214005 172896 214010 172952
rect 214066 172896 217028 172952
rect 214005 172894 217028 172896
rect 214005 172891 214071 172894
rect 231577 172818 231643 172821
rect 228988 172816 231643 172818
rect 228988 172760 231582 172816
rect 231638 172760 231643 172816
rect 228988 172758 231643 172760
rect 231577 172755 231643 172758
rect 254669 172818 254735 172821
rect 268150 172818 268210 173060
rect 254669 172816 268210 172818
rect 254669 172760 254674 172816
rect 254730 172760 268210 172816
rect 254669 172758 268210 172760
rect 254669 172755 254735 172758
rect 264973 172682 265039 172685
rect 264973 172680 268180 172682
rect 264973 172624 264978 172680
rect 265034 172624 268180 172680
rect 264973 172622 268180 172624
rect 264973 172619 265039 172622
rect 282821 172546 282887 172549
rect 279956 172544 282887 172546
rect 279956 172488 282826 172544
rect 282882 172488 282887 172544
rect 279956 172486 282887 172488
rect 282821 172483 282887 172486
rect 244365 172410 244431 172413
rect 228988 172408 244431 172410
rect 228988 172352 244370 172408
rect 244426 172352 244431 172408
rect 228988 172350 244431 172352
rect 244365 172347 244431 172350
rect 213913 172274 213979 172277
rect 265065 172274 265131 172277
rect 213913 172272 217028 172274
rect 213913 172216 213918 172272
rect 213974 172216 217028 172272
rect 213913 172214 217028 172216
rect 265065 172272 268180 172274
rect 265065 172216 265070 172272
rect 265126 172216 268180 172272
rect 265065 172214 268180 172216
rect 213913 172211 213979 172214
rect 265065 172211 265131 172214
rect 231761 171866 231827 171869
rect 228988 171864 231827 171866
rect 228988 171808 231766 171864
rect 231822 171808 231827 171864
rect 228988 171806 231827 171808
rect 231761 171803 231827 171806
rect 164724 171594 165354 171600
rect 167729 171594 167795 171597
rect 164724 171592 167795 171594
rect 164724 171540 167734 171592
rect 165294 171536 167734 171540
rect 167790 171536 167795 171592
rect 165294 171534 167795 171536
rect 167729 171531 167795 171534
rect 214005 171594 214071 171597
rect 257429 171594 257495 171597
rect 268150 171594 268210 171836
rect 281533 171730 281599 171733
rect 279956 171728 281599 171730
rect 279956 171672 281538 171728
rect 281594 171672 281599 171728
rect 279956 171670 281599 171672
rect 281533 171667 281599 171670
rect 214005 171592 217028 171594
rect 214005 171536 214010 171592
rect 214066 171536 217028 171592
rect 214005 171534 217028 171536
rect 257429 171592 268210 171594
rect 257429 171536 257434 171592
rect 257490 171536 268210 171592
rect 257429 171534 268210 171536
rect 214005 171531 214071 171534
rect 257429 171531 257495 171534
rect 231117 171458 231183 171461
rect 228988 171456 231183 171458
rect 228988 171400 231122 171456
rect 231178 171400 231183 171456
rect 228988 171398 231183 171400
rect 231117 171395 231183 171398
rect 264973 171458 265039 171461
rect 264973 171456 268180 171458
rect 264973 171400 264978 171456
rect 265034 171400 268180 171456
rect 264973 171398 268180 171400
rect 264973 171395 265039 171398
rect 214649 171050 214715 171053
rect 265065 171050 265131 171053
rect 214649 171048 217028 171050
rect 214649 170992 214654 171048
rect 214710 170992 217028 171048
rect 214649 170990 217028 170992
rect 265065 171048 268180 171050
rect 265065 170992 265070 171048
rect 265126 170992 268180 171048
rect 265065 170990 268180 170992
rect 214649 170987 214715 170990
rect 265065 170987 265131 170990
rect 232078 170914 232084 170916
rect 228988 170854 232084 170914
rect 232078 170852 232084 170854
rect 232148 170852 232154 170916
rect 281574 170914 281580 170916
rect 279956 170854 281580 170914
rect 281574 170852 281580 170854
rect 281644 170852 281650 170916
rect 230657 170506 230723 170509
rect 228988 170504 230723 170506
rect 228988 170448 230662 170504
rect 230718 170448 230723 170504
rect 228988 170446 230723 170448
rect 230657 170443 230723 170446
rect 213913 170370 213979 170373
rect 235993 170370 236059 170373
rect 251541 170370 251607 170373
rect 213913 170368 217028 170370
rect 213913 170312 213918 170368
rect 213974 170312 217028 170368
rect 213913 170310 217028 170312
rect 235993 170368 251607 170370
rect 235993 170312 235998 170368
rect 236054 170312 251546 170368
rect 251602 170312 251607 170368
rect 235993 170310 251607 170312
rect 213913 170307 213979 170310
rect 235993 170307 236059 170310
rect 251541 170307 251607 170310
rect 254577 170234 254643 170237
rect 268150 170234 268210 170476
rect 280429 170234 280495 170237
rect 254577 170232 268210 170234
rect 254577 170176 254582 170232
rect 254638 170176 268210 170232
rect 254577 170174 268210 170176
rect 279956 170232 280495 170234
rect 279956 170176 280434 170232
rect 280490 170176 280495 170232
rect 279956 170174 280495 170176
rect 254577 170171 254643 170174
rect 280429 170171 280495 170174
rect 264973 170098 265039 170101
rect 264973 170096 268180 170098
rect 264973 170040 264978 170096
rect 265034 170040 268180 170096
rect 264973 170038 268180 170040
rect 264973 170035 265039 170038
rect 231209 169962 231275 169965
rect 228988 169960 231275 169962
rect 228988 169904 231214 169960
rect 231270 169904 231275 169960
rect 228988 169902 231275 169904
rect 231209 169899 231275 169902
rect 213913 169690 213979 169693
rect 264973 169690 265039 169693
rect 213913 169688 217028 169690
rect 213913 169632 213918 169688
rect 213974 169632 217028 169688
rect 213913 169630 217028 169632
rect 264973 169688 268180 169690
rect 264973 169632 264978 169688
rect 265034 169632 268180 169688
rect 264973 169630 268180 169632
rect 213913 169627 213979 169630
rect 264973 169627 265039 169630
rect 230933 169554 230999 169557
rect 228988 169552 230999 169554
rect 228988 169496 230938 169552
rect 230994 169496 230999 169552
rect 228988 169494 230999 169496
rect 230933 169491 230999 169494
rect 281533 169418 281599 169421
rect 279956 169416 281599 169418
rect 279956 169360 281538 169416
rect 281594 169360 281599 169416
rect 279956 169358 281599 169360
rect 281533 169355 281599 169358
rect 264237 169282 264303 169285
rect 264237 169280 268180 169282
rect 264237 169224 264242 169280
rect 264298 169224 268180 169280
rect 264237 169222 268180 169224
rect 264237 169219 264303 169222
rect 214005 169010 214071 169013
rect 231669 169010 231735 169013
rect 214005 169008 217028 169010
rect 214005 168952 214010 169008
rect 214066 168952 217028 169008
rect 214005 168950 217028 168952
rect 228988 169008 231735 169010
rect 228988 168952 231674 169008
rect 231730 168952 231735 169008
rect 228988 168950 231735 168952
rect 214005 168947 214071 168950
rect 231669 168947 231735 168950
rect 265157 168874 265223 168877
rect 265157 168872 268180 168874
rect 265157 168816 265162 168872
rect 265218 168816 268180 168872
rect 265157 168814 268180 168816
rect 265157 168811 265223 168814
rect 281809 168738 281875 168741
rect 279956 168736 281875 168738
rect 279956 168680 281814 168736
rect 281870 168680 281875 168736
rect 279956 168678 281875 168680
rect 281809 168675 281875 168678
rect 241605 168602 241671 168605
rect 228988 168600 241671 168602
rect 228988 168544 241610 168600
rect 241666 168544 241671 168600
rect 228988 168542 241671 168544
rect 241605 168539 241671 168542
rect 253197 168466 253263 168469
rect 253197 168464 268180 168466
rect 253197 168408 253202 168464
rect 253258 168408 268180 168464
rect 253197 168406 268180 168408
rect 253197 168403 253263 168406
rect 213913 168330 213979 168333
rect 213913 168328 217028 168330
rect 213913 168272 213918 168328
rect 213974 168272 217028 168328
rect 213913 168270 217028 168272
rect 213913 168267 213979 168270
rect 237414 168058 237420 168060
rect 228988 167998 237420 168058
rect 237414 167996 237420 167998
rect 237484 167996 237490 168060
rect 264973 167922 265039 167925
rect 284518 167922 284524 167924
rect 264973 167920 268180 167922
rect 264973 167864 264978 167920
rect 265034 167864 268180 167920
rect 264973 167862 268180 167864
rect 279956 167862 284524 167922
rect 264973 167859 265039 167862
rect 284518 167860 284524 167862
rect 284588 167860 284594 167924
rect 214005 167650 214071 167653
rect 230933 167650 230999 167653
rect 214005 167648 217028 167650
rect 214005 167592 214010 167648
rect 214066 167592 217028 167648
rect 214005 167590 217028 167592
rect 228988 167648 230999 167650
rect 228988 167592 230938 167648
rect 230994 167592 230999 167648
rect 228988 167590 230999 167592
rect 214005 167587 214071 167590
rect 230933 167587 230999 167590
rect 279366 167588 279372 167652
rect 279436 167588 279442 167652
rect 265065 167514 265131 167517
rect 265065 167512 268180 167514
rect 265065 167456 265070 167512
rect 265126 167456 268180 167512
rect 265065 167454 268180 167456
rect 265065 167451 265131 167454
rect 231669 167106 231735 167109
rect 228988 167104 231735 167106
rect 228988 167048 231674 167104
rect 231730 167048 231735 167104
rect 228988 167046 231735 167048
rect 231669 167043 231735 167046
rect 239397 167106 239463 167109
rect 239397 167104 268180 167106
rect 239397 167048 239402 167104
rect 239458 167048 268180 167104
rect 279374 167076 279434 167588
rect 239397 167046 268180 167048
rect 239397 167043 239463 167046
rect 213913 166970 213979 166973
rect 234061 166970 234127 166973
rect 240358 166970 240364 166972
rect 213913 166968 217028 166970
rect 213913 166912 213918 166968
rect 213974 166912 217028 166968
rect 213913 166910 217028 166912
rect 234061 166968 240364 166970
rect 234061 166912 234066 166968
rect 234122 166912 240364 166968
rect 234061 166910 240364 166912
rect 213913 166907 213979 166910
rect 234061 166907 234127 166910
rect 240358 166908 240364 166910
rect 240428 166908 240434 166972
rect 236361 166698 236427 166701
rect 228988 166696 236427 166698
rect 228988 166640 236366 166696
rect 236422 166640 236427 166696
rect 228988 166638 236427 166640
rect 236361 166635 236427 166638
rect 265065 166698 265131 166701
rect 265065 166696 268180 166698
rect 265065 166640 265070 166696
rect 265126 166640 268180 166696
rect 265065 166638 268180 166640
rect 265065 166635 265131 166638
rect 214925 166426 214991 166429
rect 282821 166426 282887 166429
rect 583569 166426 583635 166429
rect 214925 166424 217028 166426
rect 214925 166368 214930 166424
rect 214986 166368 217028 166424
rect 214925 166366 217028 166368
rect 279956 166424 282887 166426
rect 279956 166368 282826 166424
rect 282882 166368 282887 166424
rect 279956 166366 282887 166368
rect 214925 166363 214991 166366
rect 282821 166363 282887 166366
rect 583526 166424 583635 166426
rect 583526 166368 583574 166424
rect 583630 166368 583635 166424
rect 583526 166363 583635 166368
rect 264973 166290 265039 166293
rect 264973 166288 268180 166290
rect 264973 166232 264978 166288
rect 265034 166232 268180 166288
rect 264973 166230 268180 166232
rect 264973 166227 265039 166230
rect 231301 166154 231367 166157
rect 228988 166152 231367 166154
rect 228988 166096 231306 166152
rect 231362 166096 231367 166152
rect 228988 166094 231367 166096
rect 231301 166091 231367 166094
rect 583526 166018 583586 166363
rect 583342 165972 583586 166018
rect 583342 165958 584960 165972
rect 279325 165882 279391 165885
rect 583342 165882 583402 165958
rect 583520 165882 584960 165958
rect 258030 165822 268180 165882
rect 279325 165880 279434 165882
rect 279325 165824 279330 165880
rect 279386 165824 279434 165880
rect 214005 165746 214071 165749
rect 231669 165746 231735 165749
rect 214005 165744 217028 165746
rect 214005 165688 214010 165744
rect 214066 165688 217028 165744
rect 214005 165686 217028 165688
rect 228988 165744 231735 165746
rect 228988 165688 231674 165744
rect 231730 165688 231735 165744
rect 228988 165686 231735 165688
rect 214005 165683 214071 165686
rect 231669 165683 231735 165686
rect 251817 165746 251883 165749
rect 258030 165746 258090 165822
rect 279325 165819 279434 165824
rect 583342 165822 584960 165882
rect 251817 165744 258090 165746
rect 251817 165688 251822 165744
rect 251878 165688 258090 165744
rect 251817 165686 258090 165688
rect 251817 165683 251883 165686
rect 232497 165610 232563 165613
rect 238937 165610 239003 165613
rect 232497 165608 239003 165610
rect 232497 165552 232502 165608
rect 232558 165552 238942 165608
rect 238998 165552 239003 165608
rect 279374 165580 279434 165819
rect 583520 165732 584960 165822
rect 232497 165550 239003 165552
rect 232497 165547 232563 165550
rect 238937 165547 239003 165550
rect 264973 165338 265039 165341
rect 264973 165336 268180 165338
rect 264973 165280 264978 165336
rect 265034 165280 268180 165336
rect 264973 165278 268180 165280
rect 264973 165275 265039 165278
rect 236494 165202 236500 165204
rect 228988 165142 236500 165202
rect 236494 165140 236500 165142
rect 236564 165140 236570 165204
rect 213913 165066 213979 165069
rect 213913 165064 217028 165066
rect 213913 165008 213918 165064
rect 213974 165008 217028 165064
rect 213913 165006 217028 165008
rect 213913 165003 213979 165006
rect 230013 164930 230079 164933
rect 246021 164930 246087 164933
rect 282821 164930 282887 164933
rect 230013 164928 246087 164930
rect 230013 164872 230018 164928
rect 230074 164872 246026 164928
rect 246082 164872 246087 164928
rect 279956 164928 282887 164930
rect 230013 164870 246087 164872
rect 230013 164867 230079 164870
rect 246021 164867 246087 164870
rect 231945 164794 232011 164797
rect 228988 164792 232011 164794
rect 228988 164736 231950 164792
rect 232006 164736 232011 164792
rect 228988 164734 232011 164736
rect 231945 164731 232011 164734
rect 267825 164658 267891 164661
rect 268150 164658 268210 164900
rect 279956 164872 282826 164928
rect 282882 164872 282887 164928
rect 279956 164870 282887 164872
rect 282821 164867 282887 164870
rect 267825 164656 268210 164658
rect 267825 164600 267830 164656
rect 267886 164600 268210 164656
rect 267825 164598 268210 164600
rect 267825 164595 267891 164598
rect 261753 164522 261819 164525
rect 261753 164520 268180 164522
rect 261753 164464 261758 164520
rect 261814 164464 268180 164520
rect 261753 164462 268180 164464
rect 261753 164459 261819 164462
rect 214005 164386 214071 164389
rect 231117 164386 231183 164389
rect 214005 164384 217028 164386
rect 214005 164328 214010 164384
rect 214066 164328 217028 164384
rect 214005 164326 217028 164328
rect 228988 164384 231183 164386
rect 228988 164328 231122 164384
rect 231178 164328 231183 164384
rect 228988 164326 231183 164328
rect 214005 164323 214071 164326
rect 231117 164323 231183 164326
rect 265617 164386 265683 164389
rect 267825 164386 267891 164389
rect 265617 164384 267891 164386
rect 265617 164328 265622 164384
rect 265678 164328 267830 164384
rect 267886 164328 267891 164384
rect 265617 164326 267891 164328
rect 265617 164323 265683 164326
rect 267825 164323 267891 164326
rect 265065 164114 265131 164117
rect 282821 164114 282887 164117
rect 265065 164112 268180 164114
rect 265065 164056 265070 164112
rect 265126 164056 268180 164112
rect 265065 164054 268180 164056
rect 279956 164112 282887 164114
rect 279956 164056 282826 164112
rect 282882 164056 282887 164112
rect 279956 164054 282887 164056
rect 265065 164051 265131 164054
rect 282821 164051 282887 164054
rect 231485 163842 231551 163845
rect 228988 163840 231551 163842
rect 228988 163784 231490 163840
rect 231546 163784 231551 163840
rect 228988 163782 231551 163784
rect 231485 163779 231551 163782
rect 213913 163706 213979 163709
rect 264973 163706 265039 163709
rect 213913 163704 217028 163706
rect 213913 163648 213918 163704
rect 213974 163648 217028 163704
rect 213913 163646 217028 163648
rect 264973 163704 268180 163706
rect 264973 163648 264978 163704
rect 265034 163648 268180 163704
rect 264973 163646 268180 163648
rect 213913 163643 213979 163646
rect 264973 163643 265039 163646
rect 232037 163434 232103 163437
rect 228988 163432 232103 163434
rect 228988 163376 232042 163432
rect 232098 163376 232103 163432
rect 228988 163374 232103 163376
rect 232037 163371 232103 163374
rect 282821 163298 282887 163301
rect 258030 163238 268180 163298
rect 279956 163296 282887 163298
rect 279956 163240 282826 163296
rect 282882 163240 282887 163296
rect 279956 163238 282887 163240
rect 235533 163162 235599 163165
rect 258030 163162 258090 163238
rect 282821 163235 282887 163238
rect 235533 163160 258090 163162
rect 235533 163104 235538 163160
rect 235594 163104 258090 163160
rect 235533 163102 258090 163104
rect 235533 163099 235599 163102
rect 214005 163026 214071 163029
rect 214005 163024 217028 163026
rect -960 162890 480 162980
rect 214005 162968 214010 163024
rect 214066 162968 217028 163024
rect 214005 162966 217028 162968
rect 214005 162963 214071 162966
rect 3233 162890 3299 162893
rect 231577 162890 231643 162893
rect -960 162888 3299 162890
rect -960 162832 3238 162888
rect 3294 162832 3299 162888
rect -960 162830 3299 162832
rect 228988 162888 231643 162890
rect 228988 162832 231582 162888
rect 231638 162832 231643 162888
rect 228988 162830 231643 162832
rect -960 162740 480 162830
rect 3233 162827 3299 162830
rect 231577 162827 231643 162830
rect 263041 162890 263107 162893
rect 263041 162888 268180 162890
rect 263041 162832 263046 162888
rect 263102 162832 268180 162888
rect 263041 162830 268180 162832
rect 263041 162827 263107 162830
rect 282821 162618 282887 162621
rect 279956 162616 282887 162618
rect 279956 162560 282826 162616
rect 282882 162560 282887 162616
rect 279956 162558 282887 162560
rect 282821 162555 282887 162558
rect 256785 162482 256851 162485
rect 228988 162480 256851 162482
rect 228988 162424 256790 162480
rect 256846 162424 256851 162480
rect 228988 162422 256851 162424
rect 256785 162419 256851 162422
rect 213913 162346 213979 162349
rect 265157 162346 265223 162349
rect 213913 162344 217028 162346
rect 213913 162288 213918 162344
rect 213974 162288 217028 162344
rect 213913 162286 217028 162288
rect 265157 162344 268180 162346
rect 265157 162288 265162 162344
rect 265218 162288 268180 162344
rect 265157 162286 268180 162288
rect 213913 162283 213979 162286
rect 265157 162283 265223 162286
rect 231761 161938 231827 161941
rect 228988 161936 231827 161938
rect 228988 161880 231766 161936
rect 231822 161880 231827 161936
rect 228988 161878 231827 161880
rect 231761 161875 231827 161878
rect 265065 161938 265131 161941
rect 265065 161936 268180 161938
rect 265065 161880 265070 161936
rect 265126 161880 268180 161936
rect 265065 161878 268180 161880
rect 265065 161875 265131 161878
rect 214005 161802 214071 161805
rect 282729 161802 282795 161805
rect 214005 161800 217028 161802
rect 214005 161744 214010 161800
rect 214066 161744 217028 161800
rect 214005 161742 217028 161744
rect 279956 161800 282795 161802
rect 279956 161744 282734 161800
rect 282790 161744 282795 161800
rect 279956 161742 282795 161744
rect 214005 161739 214071 161742
rect 282729 161739 282795 161742
rect 245929 161530 245995 161533
rect 228988 161528 245995 161530
rect 228988 161472 245934 161528
rect 245990 161472 245995 161528
rect 228988 161470 245995 161472
rect 245929 161467 245995 161470
rect 264973 161530 265039 161533
rect 264973 161528 268180 161530
rect 264973 161472 264978 161528
rect 265034 161472 268180 161528
rect 264973 161470 268180 161472
rect 264973 161467 265039 161470
rect 213913 161122 213979 161125
rect 265065 161122 265131 161125
rect 282821 161122 282887 161125
rect 213913 161120 217028 161122
rect 213913 161064 213918 161120
rect 213974 161064 217028 161120
rect 213913 161062 217028 161064
rect 265065 161120 268180 161122
rect 265065 161064 265070 161120
rect 265126 161064 268180 161120
rect 265065 161062 268180 161064
rect 279956 161120 282887 161122
rect 279956 161064 282826 161120
rect 282882 161064 282887 161120
rect 279956 161062 282887 161064
rect 213913 161059 213979 161062
rect 265065 161059 265131 161062
rect 282821 161059 282887 161062
rect 231761 160986 231827 160989
rect 228988 160984 231827 160986
rect 228988 160928 231766 160984
rect 231822 160928 231827 160984
rect 228988 160926 231827 160928
rect 231761 160923 231827 160926
rect 231577 160714 231643 160717
rect 244222 160714 244228 160716
rect 231577 160712 244228 160714
rect 231577 160656 231582 160712
rect 231638 160656 244228 160712
rect 231577 160654 244228 160656
rect 231577 160651 231643 160654
rect 244222 160652 244228 160654
rect 244292 160652 244298 160716
rect 231301 160578 231367 160581
rect 228988 160576 231367 160578
rect 228988 160520 231306 160576
rect 231362 160520 231367 160576
rect 228988 160518 231367 160520
rect 231301 160515 231367 160518
rect 214005 160442 214071 160445
rect 243629 160442 243695 160445
rect 268150 160442 268210 160684
rect 214005 160440 217028 160442
rect 214005 160384 214010 160440
rect 214066 160384 217028 160440
rect 214005 160382 217028 160384
rect 243629 160440 268210 160442
rect 243629 160384 243634 160440
rect 243690 160384 268210 160440
rect 243629 160382 268210 160384
rect 214005 160379 214071 160382
rect 243629 160379 243695 160382
rect 264973 160306 265039 160309
rect 282729 160306 282795 160309
rect 264973 160304 268180 160306
rect 264973 160248 264978 160304
rect 265034 160248 268180 160304
rect 264973 160246 268180 160248
rect 279956 160304 282795 160306
rect 279956 160248 282734 160304
rect 282790 160248 282795 160304
rect 279956 160246 282795 160248
rect 264973 160243 265039 160246
rect 282729 160243 282795 160246
rect 231761 160034 231827 160037
rect 228988 160032 231827 160034
rect 228988 159976 231766 160032
rect 231822 159976 231827 160032
rect 228988 159974 231827 159976
rect 231761 159971 231827 159974
rect 213913 159762 213979 159765
rect 265065 159762 265131 159765
rect 213913 159760 217028 159762
rect 213913 159704 213918 159760
rect 213974 159704 217028 159760
rect 213913 159702 217028 159704
rect 265065 159760 268180 159762
rect 265065 159704 265070 159760
rect 265126 159704 268180 159760
rect 265065 159702 268180 159704
rect 213913 159699 213979 159702
rect 265065 159699 265131 159702
rect 231669 159626 231735 159629
rect 228988 159624 231735 159626
rect 228988 159568 231674 159624
rect 231730 159568 231735 159624
rect 228988 159566 231735 159568
rect 231669 159563 231735 159566
rect 282545 159490 282611 159493
rect 279956 159488 282611 159490
rect 279956 159432 282550 159488
rect 282606 159432 282611 159488
rect 279956 159430 282611 159432
rect 282545 159427 282611 159430
rect 214005 159082 214071 159085
rect 231577 159082 231643 159085
rect 214005 159080 217028 159082
rect 214005 159024 214010 159080
rect 214066 159024 217028 159080
rect 214005 159022 217028 159024
rect 228988 159080 231643 159082
rect 228988 159024 231582 159080
rect 231638 159024 231643 159080
rect 228988 159022 231643 159024
rect 214005 159019 214071 159022
rect 231577 159019 231643 159022
rect 233734 159020 233740 159084
rect 233804 159082 233810 159084
rect 268150 159082 268210 159324
rect 233804 159022 268210 159082
rect 233804 159020 233810 159022
rect 264973 158946 265039 158949
rect 264973 158944 268180 158946
rect 264973 158888 264978 158944
rect 265034 158888 268180 158944
rect 264973 158886 268180 158888
rect 264973 158883 265039 158886
rect 282453 158810 282519 158813
rect 279956 158808 282519 158810
rect 279956 158752 282458 158808
rect 282514 158752 282519 158808
rect 279956 158750 282519 158752
rect 282453 158747 282519 158750
rect 230933 158674 230999 158677
rect 228988 158672 230999 158674
rect 228988 158616 230938 158672
rect 230994 158616 230999 158672
rect 228988 158614 230999 158616
rect 230933 158611 230999 158614
rect 264973 158538 265039 158541
rect 264973 158536 268180 158538
rect 264973 158480 264978 158536
rect 265034 158480 268180 158536
rect 264973 158478 268180 158480
rect 264973 158475 265039 158478
rect 213913 158402 213979 158405
rect 213913 158400 217028 158402
rect 213913 158344 213918 158400
rect 213974 158344 217028 158400
rect 213913 158342 217028 158344
rect 213913 158339 213979 158342
rect 229737 158130 229803 158133
rect 228988 158128 229803 158130
rect 228988 158072 229742 158128
rect 229798 158072 229803 158128
rect 228988 158070 229803 158072
rect 229737 158067 229803 158070
rect 265157 158130 265223 158133
rect 265157 158128 268180 158130
rect 265157 158072 265162 158128
rect 265218 158072 268180 158128
rect 265157 158070 268180 158072
rect 265157 158067 265223 158070
rect 232630 157932 232636 157996
rect 232700 157994 232706 157996
rect 252553 157994 252619 157997
rect 282085 157994 282151 157997
rect 232700 157992 252619 157994
rect 232700 157936 252558 157992
rect 252614 157936 252619 157992
rect 232700 157934 252619 157936
rect 279956 157992 282151 157994
rect 279956 157936 282090 157992
rect 282146 157936 282151 157992
rect 279956 157934 282151 157936
rect 232700 157932 232706 157934
rect 252553 157931 252619 157934
rect 282085 157931 282151 157934
rect 214005 157722 214071 157725
rect 231485 157722 231551 157725
rect 214005 157720 217028 157722
rect 214005 157664 214010 157720
rect 214066 157664 217028 157720
rect 214005 157662 217028 157664
rect 228988 157720 231551 157722
rect 228988 157664 231490 157720
rect 231546 157664 231551 157720
rect 228988 157662 231551 157664
rect 214005 157659 214071 157662
rect 231485 157659 231551 157662
rect 258030 157662 268180 157722
rect 236821 157586 236887 157589
rect 258030 157586 258090 157662
rect 236821 157584 258090 157586
rect 236821 157528 236826 157584
rect 236882 157528 258090 157584
rect 236821 157526 258090 157528
rect 236821 157523 236887 157526
rect 231117 157450 231183 157453
rect 231894 157450 231900 157452
rect 231117 157448 231900 157450
rect 231117 157392 231122 157448
rect 231178 157392 231900 157448
rect 231117 157390 231900 157392
rect 231117 157387 231183 157390
rect 231894 157388 231900 157390
rect 231964 157388 231970 157452
rect 281901 157314 281967 157317
rect 279956 157312 281967 157314
rect 279956 157256 281906 157312
rect 281962 157256 281967 157312
rect 279956 157254 281967 157256
rect 281901 157251 281967 157254
rect 213913 157178 213979 157181
rect 234613 157178 234679 157181
rect 213913 157176 217028 157178
rect 213913 157120 213918 157176
rect 213974 157120 217028 157176
rect 213913 157118 217028 157120
rect 228988 157176 234679 157178
rect 228988 157120 234618 157176
rect 234674 157120 234679 157176
rect 228988 157118 234679 157120
rect 213913 157115 213979 157118
rect 234613 157115 234679 157118
rect 265065 157178 265131 157181
rect 265065 157176 268180 157178
rect 265065 157120 265070 157176
rect 265126 157120 268180 157176
rect 265065 157118 268180 157120
rect 265065 157115 265131 157118
rect 231761 156770 231827 156773
rect 228988 156768 231827 156770
rect 228988 156712 231766 156768
rect 231822 156712 231827 156768
rect 228988 156710 231827 156712
rect 231761 156707 231827 156710
rect 264973 156770 265039 156773
rect 264973 156768 268180 156770
rect 264973 156712 264978 156768
rect 265034 156712 268180 156768
rect 264973 156710 268180 156712
rect 264973 156707 265039 156710
rect 242249 156634 242315 156637
rect 265157 156634 265223 156637
rect 242249 156632 265223 156634
rect 242249 156576 242254 156632
rect 242310 156576 265162 156632
rect 265218 156576 265223 156632
rect 242249 156574 265223 156576
rect 242249 156571 242315 156574
rect 265157 156571 265223 156574
rect 214005 156498 214071 156501
rect 214005 156496 217028 156498
rect 214005 156440 214010 156496
rect 214066 156440 217028 156496
rect 214005 156438 217028 156440
rect 214005 156435 214071 156438
rect 265709 156362 265775 156365
rect 265709 156360 268180 156362
rect 265709 156304 265714 156360
rect 265770 156304 268180 156360
rect 265709 156302 268180 156304
rect 265709 156299 265775 156302
rect 248505 156226 248571 156229
rect 228988 156224 248571 156226
rect 228988 156168 248510 156224
rect 248566 156168 248571 156224
rect 228988 156166 248571 156168
rect 248505 156163 248571 156166
rect 279926 156090 279986 156468
rect 291326 156090 291332 156092
rect 279926 156030 291332 156090
rect 291326 156028 291332 156030
rect 291396 156028 291402 156092
rect 265157 155954 265223 155957
rect 265157 155952 268180 155954
rect 265157 155896 265162 155952
rect 265218 155896 268180 155952
rect 265157 155894 268180 155896
rect 265157 155891 265223 155894
rect 213913 155818 213979 155821
rect 231485 155818 231551 155821
rect 213913 155816 217028 155818
rect 213913 155760 213918 155816
rect 213974 155760 217028 155816
rect 213913 155758 217028 155760
rect 228988 155816 231551 155818
rect 228988 155760 231490 155816
rect 231546 155760 231551 155816
rect 228988 155758 231551 155760
rect 213913 155755 213979 155758
rect 231485 155755 231551 155758
rect 282821 155682 282887 155685
rect 279956 155680 282887 155682
rect 279956 155624 282826 155680
rect 282882 155624 282887 155680
rect 279956 155622 282887 155624
rect 282821 155619 282887 155622
rect 265801 155546 265867 155549
rect 265801 155544 268180 155546
rect 265801 155488 265806 155544
rect 265862 155488 268180 155544
rect 265801 155486 268180 155488
rect 265801 155483 265867 155486
rect 230749 155274 230815 155277
rect 228988 155272 230815 155274
rect 228988 155216 230754 155272
rect 230810 155216 230815 155272
rect 228988 155214 230815 155216
rect 230749 155211 230815 155214
rect 166206 154532 166212 154596
rect 166276 154594 166282 154596
rect 216998 154594 217058 155108
rect 258030 155078 268180 155138
rect 232681 155002 232747 155005
rect 258030 155002 258090 155078
rect 282177 155002 282243 155005
rect 232681 155000 258090 155002
rect 232681 154944 232686 155000
rect 232742 154944 258090 155000
rect 232681 154942 258090 154944
rect 279956 155000 282243 155002
rect 279956 154944 282182 155000
rect 282238 154944 282243 155000
rect 279956 154942 282243 154944
rect 232681 154939 232747 154942
rect 282177 154939 282243 154942
rect 233877 154866 233943 154869
rect 228988 154864 233943 154866
rect 228988 154808 233882 154864
rect 233938 154808 233943 154864
rect 228988 154806 233943 154808
rect 233877 154803 233943 154806
rect 166276 154534 217058 154594
rect 264973 154594 265039 154597
rect 264973 154592 268180 154594
rect 264973 154536 264978 154592
rect 265034 154536 268180 154592
rect 264973 154534 268180 154536
rect 166276 154532 166282 154534
rect 264973 154531 265039 154534
rect 214833 154458 214899 154461
rect 214833 154456 217028 154458
rect 214833 154400 214838 154456
rect 214894 154400 217028 154456
rect 214833 154398 217028 154400
rect 214833 154395 214899 154398
rect 231669 154322 231735 154325
rect 228988 154320 231735 154322
rect 228988 154264 231674 154320
rect 231730 154264 231735 154320
rect 228988 154262 231735 154264
rect 231669 154259 231735 154262
rect 266261 154186 266327 154189
rect 282085 154186 282151 154189
rect 266261 154184 268180 154186
rect 266261 154128 266266 154184
rect 266322 154128 268180 154184
rect 266261 154126 268180 154128
rect 279956 154184 282151 154186
rect 279956 154128 282090 154184
rect 282146 154128 282151 154184
rect 279956 154126 282151 154128
rect 266261 154123 266327 154126
rect 282085 154123 282151 154126
rect 231761 153914 231827 153917
rect 228988 153912 231827 153914
rect 228988 153856 231766 153912
rect 231822 153856 231827 153912
rect 228988 153854 231827 153856
rect 231761 153851 231827 153854
rect 213913 153778 213979 153781
rect 229737 153778 229803 153781
rect 238886 153778 238892 153780
rect 213913 153776 217028 153778
rect 213913 153720 213918 153776
rect 213974 153720 217028 153776
rect 213913 153718 217028 153720
rect 229737 153776 238892 153778
rect 229737 153720 229742 153776
rect 229798 153720 238892 153776
rect 229737 153718 238892 153720
rect 213913 153715 213979 153718
rect 229737 153715 229803 153718
rect 238886 153716 238892 153718
rect 238956 153716 238962 153780
rect 265249 153778 265315 153781
rect 265249 153776 268180 153778
rect 265249 153720 265254 153776
rect 265310 153720 268180 153776
rect 265249 153718 268180 153720
rect 265249 153715 265315 153718
rect 282361 153506 282427 153509
rect 279956 153504 282427 153506
rect 279956 153448 282366 153504
rect 282422 153448 282427 153504
rect 279956 153446 282427 153448
rect 282361 153443 282427 153446
rect 231577 153370 231643 153373
rect 228988 153368 231643 153370
rect 228988 153312 231582 153368
rect 231638 153312 231643 153368
rect 228988 153310 231643 153312
rect 231577 153307 231643 153310
rect 258030 153310 268180 153370
rect 235441 153234 235507 153237
rect 258030 153234 258090 153310
rect 235441 153232 258090 153234
rect 235441 153176 235446 153232
rect 235502 153176 258090 153232
rect 235441 153174 258090 153176
rect 235441 153171 235507 153174
rect 213913 153098 213979 153101
rect 231761 153098 231827 153101
rect 259453 153098 259519 153101
rect 213913 153096 217028 153098
rect 213913 153040 213918 153096
rect 213974 153040 217028 153096
rect 213913 153038 217028 153040
rect 231761 153096 259519 153098
rect 231761 153040 231766 153096
rect 231822 153040 259458 153096
rect 259514 153040 259519 153096
rect 231761 153038 259519 153040
rect 213913 153035 213979 153038
rect 231761 153035 231827 153038
rect 259453 153035 259519 153038
rect 231853 152962 231919 152965
rect 228988 152960 231919 152962
rect 228988 152904 231858 152960
rect 231914 152904 231919 152960
rect 228988 152902 231919 152904
rect 231853 152899 231919 152902
rect 265065 152962 265131 152965
rect 265065 152960 268180 152962
rect 265065 152904 265070 152960
rect 265126 152904 268180 152960
rect 265065 152902 268180 152904
rect 265065 152899 265131 152902
rect 281717 152690 281783 152693
rect 279956 152688 281783 152690
rect 279956 152632 281722 152688
rect 281778 152632 281783 152688
rect 279956 152630 281783 152632
rect 281717 152627 281783 152630
rect 583293 152690 583359 152693
rect 583520 152690 584960 152780
rect 583293 152688 584960 152690
rect 583293 152632 583298 152688
rect 583354 152632 584960 152688
rect 583293 152630 584960 152632
rect 583293 152627 583359 152630
rect 214005 152554 214071 152557
rect 230657 152554 230723 152557
rect 214005 152552 217028 152554
rect 214005 152496 214010 152552
rect 214066 152496 217028 152552
rect 214005 152494 217028 152496
rect 228988 152552 230723 152554
rect 228988 152496 230662 152552
rect 230718 152496 230723 152552
rect 228988 152494 230723 152496
rect 214005 152491 214071 152494
rect 230657 152491 230723 152494
rect 264973 152554 265039 152557
rect 264973 152552 268180 152554
rect 264973 152496 264978 152552
rect 265034 152496 268180 152552
rect 583520 152540 584960 152630
rect 264973 152494 268180 152496
rect 264973 152491 265039 152494
rect 230974 152356 230980 152420
rect 231044 152418 231050 152420
rect 240869 152418 240935 152421
rect 231044 152416 240935 152418
rect 231044 152360 240874 152416
rect 240930 152360 240935 152416
rect 231044 152358 240935 152360
rect 231044 152356 231050 152358
rect 240869 152355 240935 152358
rect 231761 152010 231827 152013
rect 228988 152008 231827 152010
rect 228988 151952 231766 152008
rect 231822 151952 231827 152008
rect 228988 151950 231827 151952
rect 231761 151947 231827 151950
rect 258809 152010 258875 152013
rect 258809 152008 268180 152010
rect 258809 151952 258814 152008
rect 258870 151952 268180 152008
rect 258809 151950 268180 151952
rect 258809 151947 258875 151950
rect 215937 151874 216003 151877
rect 215937 151872 217028 151874
rect 215937 151816 215942 151872
rect 215998 151816 217028 151872
rect 215937 151814 217028 151816
rect 215937 151811 216003 151814
rect 244774 151812 244780 151876
rect 244844 151874 244850 151876
rect 249742 151874 249748 151876
rect 244844 151814 249748 151874
rect 244844 151812 244850 151814
rect 249742 151812 249748 151814
rect 249812 151812 249818 151876
rect 281625 151874 281691 151877
rect 279956 151872 281691 151874
rect 279956 151816 281630 151872
rect 281686 151816 281691 151872
rect 279956 151814 281691 151816
rect 281625 151811 281691 151814
rect 231117 151602 231183 151605
rect 228988 151600 231183 151602
rect 228988 151544 231122 151600
rect 231178 151544 231183 151600
rect 228988 151542 231183 151544
rect 231117 151539 231183 151542
rect 264973 151602 265039 151605
rect 264973 151600 268180 151602
rect 264973 151544 264978 151600
rect 265034 151544 268180 151600
rect 264973 151542 268180 151544
rect 264973 151539 265039 151542
rect 214005 151194 214071 151197
rect 214005 151192 217028 151194
rect 214005 151136 214010 151192
rect 214066 151136 217028 151192
rect 214005 151134 217028 151136
rect 214005 151131 214071 151134
rect 232998 151132 233004 151196
rect 233068 151194 233074 151196
rect 242014 151194 242020 151196
rect 233068 151134 242020 151194
rect 233068 151132 233074 151134
rect 242014 151132 242020 151134
rect 242084 151132 242090 151196
rect 265065 151194 265131 151197
rect 282821 151194 282887 151197
rect 265065 151192 268180 151194
rect 265065 151136 265070 151192
rect 265126 151136 268180 151192
rect 265065 151134 268180 151136
rect 279956 151192 282887 151194
rect 279956 151136 282826 151192
rect 282882 151136 282887 151192
rect 279956 151134 282887 151136
rect 265065 151131 265131 151134
rect 282821 151131 282887 151134
rect 231761 151058 231827 151061
rect 248597 151058 248663 151061
rect 228988 151056 231827 151058
rect 228988 151000 231766 151056
rect 231822 151000 231827 151056
rect 228988 150998 231827 151000
rect 231761 150995 231827 150998
rect 238710 151056 248663 151058
rect 238710 151000 248602 151056
rect 248658 151000 248663 151056
rect 238710 150998 248663 151000
rect 231669 150922 231735 150925
rect 238710 150922 238770 150998
rect 248597 150995 248663 150998
rect 231669 150920 238770 150922
rect 231669 150864 231674 150920
rect 231730 150864 238770 150920
rect 231669 150862 238770 150864
rect 231669 150859 231735 150862
rect 249149 150786 249215 150789
rect 249149 150784 268180 150786
rect 249149 150728 249154 150784
rect 249210 150728 268180 150784
rect 249149 150726 268180 150728
rect 249149 150723 249215 150726
rect 229369 150650 229435 150653
rect 228988 150648 229435 150650
rect 228988 150592 229374 150648
rect 229430 150592 229435 150648
rect 228988 150590 229435 150592
rect 229369 150587 229435 150590
rect 279325 150650 279391 150653
rect 279325 150648 279434 150650
rect 279325 150592 279330 150648
rect 279386 150592 279434 150648
rect 279325 150587 279434 150592
rect 213913 150514 213979 150517
rect 213913 150512 217028 150514
rect 213913 150456 213918 150512
rect 213974 150456 217028 150512
rect 213913 150454 217028 150456
rect 213913 150451 213979 150454
rect 264973 150378 265039 150381
rect 264973 150376 268180 150378
rect 264973 150320 264978 150376
rect 265034 150320 268180 150376
rect 279374 150348 279434 150587
rect 264973 150318 268180 150320
rect 264973 150315 265039 150318
rect 231761 150106 231827 150109
rect 228988 150104 231827 150106
rect 228988 150048 231766 150104
rect 231822 150048 231827 150104
rect 228988 150046 231827 150048
rect 231761 150043 231827 150046
rect 265157 149970 265223 149973
rect 265157 149968 268180 149970
rect -960 149834 480 149924
rect 265157 149912 265162 149968
rect 265218 149912 268180 149968
rect 265157 149910 268180 149912
rect 265157 149907 265223 149910
rect 2773 149834 2839 149837
rect -960 149832 2839 149834
rect -960 149776 2778 149832
rect 2834 149776 2839 149832
rect -960 149774 2839 149776
rect -960 149684 480 149774
rect 2773 149771 2839 149774
rect 214557 149834 214623 149837
rect 214557 149832 217028 149834
rect 214557 149776 214562 149832
rect 214618 149776 217028 149832
rect 214557 149774 217028 149776
rect 214557 149771 214623 149774
rect 229134 149698 229140 149700
rect 228988 149638 229140 149698
rect 229134 149636 229140 149638
rect 229204 149636 229210 149700
rect 258030 149502 268180 149562
rect 240869 149426 240935 149429
rect 258030 149426 258090 149502
rect 240869 149424 258090 149426
rect 240869 149368 240874 149424
rect 240930 149368 258090 149424
rect 240869 149366 258090 149368
rect 240869 149363 240935 149366
rect 214005 149154 214071 149157
rect 231485 149154 231551 149157
rect 214005 149152 217028 149154
rect 214005 149096 214010 149152
rect 214066 149096 217028 149152
rect 214005 149094 217028 149096
rect 228988 149152 231551 149154
rect 228988 149096 231490 149152
rect 231546 149096 231551 149152
rect 228988 149094 231551 149096
rect 279926 149154 279986 149668
rect 287278 149154 287284 149156
rect 279926 149094 287284 149154
rect 214005 149091 214071 149094
rect 231485 149091 231551 149094
rect 287278 149092 287284 149094
rect 287348 149092 287354 149156
rect 264973 149018 265039 149021
rect 264973 149016 268180 149018
rect 264973 148960 264978 149016
rect 265034 148960 268180 149016
rect 264973 148958 268180 148960
rect 264973 148955 265039 148958
rect 281533 148882 281599 148885
rect 279956 148880 281599 148882
rect 279956 148824 281538 148880
rect 281594 148824 281599 148880
rect 279956 148822 281599 148824
rect 281533 148819 281599 148822
rect 230749 148746 230815 148749
rect 228988 148744 230815 148746
rect 228988 148688 230754 148744
rect 230810 148688 230815 148744
rect 228988 148686 230815 148688
rect 230749 148683 230815 148686
rect 265617 148610 265683 148613
rect 265617 148608 268180 148610
rect 265617 148552 265622 148608
rect 265678 148552 268180 148608
rect 265617 148550 268180 148552
rect 265617 148547 265683 148550
rect 213913 148474 213979 148477
rect 213913 148472 217028 148474
rect 213913 148416 213918 148472
rect 213974 148416 217028 148472
rect 213913 148414 217028 148416
rect 213913 148411 213979 148414
rect 229921 148338 229987 148341
rect 259085 148338 259151 148341
rect 229921 148336 259151 148338
rect 229921 148280 229926 148336
rect 229982 148280 259090 148336
rect 259146 148280 259151 148336
rect 229921 148278 259151 148280
rect 229921 148275 229987 148278
rect 259085 148275 259151 148278
rect 231761 148202 231827 148205
rect 228988 148200 231827 148202
rect 228988 148144 231766 148200
rect 231822 148144 231827 148200
rect 228988 148142 231827 148144
rect 231761 148139 231827 148142
rect 258030 148142 268180 148202
rect 242014 148004 242020 148068
rect 242084 148066 242090 148068
rect 258030 148066 258090 148142
rect 282821 148066 282887 148069
rect 242084 148006 258090 148066
rect 279956 148064 282887 148066
rect 279956 148008 282826 148064
rect 282882 148008 282887 148064
rect 279956 148006 282887 148008
rect 242084 148004 242090 148006
rect 282821 148003 282887 148006
rect 213913 147930 213979 147933
rect 259085 147930 259151 147933
rect 213913 147928 217028 147930
rect 213913 147872 213918 147928
rect 213974 147872 217028 147928
rect 213913 147870 217028 147872
rect 259085 147928 268210 147930
rect 259085 147872 259090 147928
rect 259146 147872 268210 147928
rect 259085 147870 268210 147872
rect 213913 147867 213979 147870
rect 259085 147867 259151 147870
rect 230841 147794 230907 147797
rect 228988 147792 230907 147794
rect 228988 147736 230846 147792
rect 230902 147736 230907 147792
rect 268150 147764 268210 147870
rect 228988 147734 230907 147736
rect 230841 147731 230907 147734
rect 265893 147386 265959 147389
rect 282821 147386 282887 147389
rect 265893 147384 268180 147386
rect 265893 147328 265898 147384
rect 265954 147328 268180 147384
rect 265893 147326 268180 147328
rect 279956 147384 282887 147386
rect 279956 147328 282826 147384
rect 282882 147328 282887 147384
rect 279956 147326 282887 147328
rect 265893 147323 265959 147326
rect 282821 147323 282887 147326
rect 213913 147250 213979 147253
rect 231669 147250 231735 147253
rect 213913 147248 217028 147250
rect 213913 147192 213918 147248
rect 213974 147192 217028 147248
rect 213913 147190 217028 147192
rect 228988 147248 231735 147250
rect 228988 147192 231674 147248
rect 231730 147192 231735 147248
rect 228988 147190 231735 147192
rect 213913 147187 213979 147190
rect 231669 147187 231735 147190
rect 279417 147114 279483 147117
rect 279374 147112 279483 147114
rect 279374 147056 279422 147112
rect 279478 147056 279483 147112
rect 279374 147051 279483 147056
rect 231393 146978 231459 146981
rect 241513 146978 241579 146981
rect 231393 146976 241579 146978
rect 231393 146920 231398 146976
rect 231454 146920 241518 146976
rect 241574 146920 241579 146976
rect 231393 146918 241579 146920
rect 231393 146915 231459 146918
rect 241513 146915 241579 146918
rect 229093 146842 229159 146845
rect 228988 146840 229159 146842
rect 228988 146784 229098 146840
rect 229154 146784 229159 146840
rect 228988 146782 229159 146784
rect 229093 146779 229159 146782
rect 216029 146570 216095 146573
rect 257521 146570 257587 146573
rect 268150 146570 268210 146948
rect 216029 146568 217028 146570
rect 216029 146512 216034 146568
rect 216090 146512 217028 146568
rect 216029 146510 217028 146512
rect 257521 146568 268210 146570
rect 257521 146512 257526 146568
rect 257582 146512 268210 146568
rect 279374 146540 279434 147051
rect 257521 146510 268210 146512
rect 216029 146507 216095 146510
rect 257521 146507 257587 146510
rect 265157 146434 265223 146437
rect 265157 146432 268180 146434
rect 265157 146376 265162 146432
rect 265218 146376 268180 146432
rect 265157 146374 268180 146376
rect 265157 146371 265223 146374
rect 231761 146298 231827 146301
rect 228988 146296 231827 146298
rect 228988 146240 231766 146296
rect 231822 146240 231827 146296
rect 228988 146238 231827 146240
rect 231761 146235 231827 146238
rect 265065 146026 265131 146029
rect 265065 146024 268180 146026
rect 265065 145968 265070 146024
rect 265126 145968 268180 146024
rect 265065 145966 268180 145968
rect 265065 145963 265131 145966
rect 213913 145890 213979 145893
rect 230749 145890 230815 145893
rect 280153 145890 280219 145893
rect 213913 145888 217028 145890
rect 213913 145832 213918 145888
rect 213974 145832 217028 145888
rect 213913 145830 217028 145832
rect 228988 145888 230815 145890
rect 228988 145832 230754 145888
rect 230810 145832 230815 145888
rect 228988 145830 230815 145832
rect 279956 145888 280219 145890
rect 279956 145832 280158 145888
rect 280214 145832 280219 145888
rect 279956 145830 280219 145832
rect 213913 145827 213979 145830
rect 230749 145827 230815 145830
rect 280153 145827 280219 145830
rect 230422 145346 230428 145348
rect 228988 145286 230428 145346
rect 230422 145284 230428 145286
rect 230492 145284 230498 145348
rect 242341 145346 242407 145349
rect 268150 145346 268210 145588
rect 242341 145344 268210 145346
rect 242341 145288 242346 145344
rect 242402 145288 268210 145344
rect 242341 145286 268210 145288
rect 242341 145283 242407 145286
rect 214465 145210 214531 145213
rect 264973 145210 265039 145213
rect 214465 145208 217028 145210
rect 214465 145152 214470 145208
rect 214526 145152 217028 145208
rect 214465 145150 217028 145152
rect 264973 145208 268180 145210
rect 264973 145152 264978 145208
rect 265034 145152 268180 145208
rect 264973 145150 268180 145152
rect 214465 145147 214531 145150
rect 264973 145147 265039 145150
rect 282269 145074 282335 145077
rect 279956 145072 282335 145074
rect 279956 145016 282274 145072
rect 282330 145016 282335 145072
rect 279956 145014 282335 145016
rect 282269 145011 282335 145014
rect 238753 144938 238819 144941
rect 228988 144936 238819 144938
rect 228988 144880 238758 144936
rect 238814 144880 238819 144936
rect 228988 144878 238819 144880
rect 238753 144875 238819 144878
rect 231761 144802 231827 144805
rect 245745 144802 245811 144805
rect 231761 144800 245811 144802
rect 231761 144744 231766 144800
rect 231822 144744 245750 144800
rect 245806 144744 245811 144800
rect 231761 144742 245811 144744
rect 231761 144739 231827 144742
rect 245745 144739 245811 144742
rect 264973 144802 265039 144805
rect 264973 144800 268180 144802
rect 264973 144744 264978 144800
rect 265034 144744 268180 144800
rect 264973 144742 268180 144744
rect 264973 144739 265039 144742
rect 230749 144666 230815 144669
rect 240726 144666 240732 144668
rect 230749 144664 240732 144666
rect 230749 144608 230754 144664
rect 230810 144608 240732 144664
rect 230749 144606 240732 144608
rect 230749 144603 230815 144606
rect 240726 144604 240732 144606
rect 240796 144604 240802 144668
rect 214005 144530 214071 144533
rect 214005 144528 217028 144530
rect 214005 144472 214010 144528
rect 214066 144472 217028 144528
rect 214005 144470 217028 144472
rect 214005 144467 214071 144470
rect 231301 144394 231367 144397
rect 228988 144392 231367 144394
rect 228988 144336 231306 144392
rect 231362 144336 231367 144392
rect 228988 144334 231367 144336
rect 231301 144331 231367 144334
rect 230749 143986 230815 143989
rect 228988 143984 230815 143986
rect 228988 143928 230754 143984
rect 230810 143928 230815 143984
rect 228988 143926 230815 143928
rect 230749 143923 230815 143926
rect 250478 143924 250484 143988
rect 250548 143986 250554 143988
rect 268150 143986 268210 144364
rect 281901 144258 281967 144261
rect 279956 144256 281967 144258
rect 279956 144200 281906 144256
rect 281962 144200 281967 144256
rect 279956 144198 281967 144200
rect 281901 144195 281967 144198
rect 250548 143926 268210 143986
rect 250548 143924 250554 143926
rect 213913 143850 213979 143853
rect 265249 143850 265315 143853
rect 213913 143848 217028 143850
rect 213913 143792 213918 143848
rect 213974 143792 217028 143848
rect 213913 143790 217028 143792
rect 265249 143848 268180 143850
rect 265249 143792 265254 143848
rect 265310 143792 268180 143848
rect 265249 143790 268180 143792
rect 213913 143787 213979 143790
rect 265249 143787 265315 143790
rect 282453 143578 282519 143581
rect 279956 143576 282519 143578
rect 279956 143520 282458 143576
rect 282514 143520 282519 143576
rect 279956 143518 282519 143520
rect 282453 143515 282519 143518
rect 230289 143442 230355 143445
rect 228988 143440 230355 143442
rect 228988 143384 230294 143440
rect 230350 143384 230355 143440
rect 228988 143382 230355 143384
rect 230289 143379 230355 143382
rect 264973 143442 265039 143445
rect 264973 143440 268180 143442
rect 264973 143384 264978 143440
rect 265034 143384 268180 143440
rect 264973 143382 268180 143384
rect 264973 143379 265039 143382
rect 213913 143306 213979 143309
rect 213913 143304 217028 143306
rect 213913 143248 213918 143304
rect 213974 143248 217028 143304
rect 213913 143246 217028 143248
rect 213913 143243 213979 143246
rect 231761 143034 231827 143037
rect 228988 143032 231827 143034
rect 228988 142976 231766 143032
rect 231822 142976 231827 143032
rect 228988 142974 231827 142976
rect 231761 142971 231827 142974
rect 265157 143034 265223 143037
rect 265157 143032 268180 143034
rect 265157 142976 265162 143032
rect 265218 142976 268180 143032
rect 265157 142974 268180 142976
rect 265157 142971 265223 142974
rect 169518 142700 169524 142764
rect 169588 142762 169594 142764
rect 202229 142762 202295 142765
rect 169588 142760 202295 142762
rect 169588 142704 202234 142760
rect 202290 142704 202295 142760
rect 169588 142702 202295 142704
rect 169588 142700 169594 142702
rect 202229 142699 202295 142702
rect 231158 142700 231164 142764
rect 231228 142762 231234 142764
rect 245193 142762 245259 142765
rect 282085 142762 282151 142765
rect 231228 142760 245259 142762
rect 231228 142704 245198 142760
rect 245254 142704 245259 142760
rect 231228 142702 245259 142704
rect 279956 142760 282151 142762
rect 279956 142704 282090 142760
rect 282146 142704 282151 142760
rect 279956 142702 282151 142704
rect 231228 142700 231234 142702
rect 245193 142699 245259 142702
rect 282085 142699 282151 142702
rect 214005 142626 214071 142629
rect 214005 142624 217028 142626
rect 214005 142568 214010 142624
rect 214066 142568 217028 142624
rect 214005 142566 217028 142568
rect 258030 142566 268180 142626
rect 214005 142563 214071 142566
rect 232998 142490 233004 142492
rect 228988 142430 233004 142490
rect 232998 142428 233004 142430
rect 233068 142428 233074 142492
rect 245009 142490 245075 142493
rect 258030 142490 258090 142566
rect 245009 142488 258090 142490
rect 245009 142432 245014 142488
rect 245070 142432 258090 142488
rect 245009 142430 258090 142432
rect 245009 142427 245075 142430
rect 265065 142218 265131 142221
rect 265065 142216 268180 142218
rect 265065 142160 265070 142216
rect 265126 142160 268180 142216
rect 265065 142158 268180 142160
rect 265065 142155 265131 142158
rect 232630 142082 232636 142084
rect 228988 142022 232636 142082
rect 232630 142020 232636 142022
rect 232700 142020 232706 142084
rect 281901 142082 281967 142085
rect 279956 142080 281967 142082
rect 279956 142024 281906 142080
rect 281962 142024 281967 142080
rect 279956 142022 281967 142024
rect 281901 142019 281967 142022
rect 213269 141946 213335 141949
rect 213269 141944 217028 141946
rect 213269 141888 213274 141944
rect 213330 141888 217028 141944
rect 213269 141886 217028 141888
rect 213269 141883 213335 141886
rect 265341 141810 265407 141813
rect 265341 141808 268180 141810
rect 265341 141752 265346 141808
rect 265402 141752 268180 141808
rect 265341 141750 268180 141752
rect 265341 141747 265407 141750
rect 231301 141674 231367 141677
rect 228988 141672 231367 141674
rect 228988 141616 231306 141672
rect 231362 141616 231367 141672
rect 228988 141614 231367 141616
rect 231301 141611 231367 141614
rect 282269 141266 282335 141269
rect 170397 140858 170463 140861
rect 216998 140858 217058 141236
rect 258030 141206 268180 141266
rect 279956 141264 282335 141266
rect 279956 141208 282274 141264
rect 282330 141208 282335 141264
rect 279956 141206 282335 141208
rect 229737 141130 229803 141133
rect 228988 141128 229803 141130
rect 228988 141072 229742 141128
rect 229798 141072 229803 141128
rect 228988 141070 229803 141072
rect 229737 141067 229803 141070
rect 232446 141068 232452 141132
rect 232516 141130 232522 141132
rect 258030 141130 258090 141206
rect 282269 141203 282335 141206
rect 232516 141070 258090 141130
rect 232516 141068 232522 141070
rect 170397 140856 217058 140858
rect 170397 140800 170402 140856
rect 170458 140800 217058 140856
rect 170397 140798 217058 140800
rect 264973 140858 265039 140861
rect 264973 140856 268180 140858
rect 264973 140800 264978 140856
rect 265034 140800 268180 140856
rect 264973 140798 268180 140800
rect 170397 140795 170463 140798
rect 264973 140795 265039 140798
rect 230657 140722 230723 140725
rect 228988 140720 230723 140722
rect 228988 140664 230662 140720
rect 230718 140664 230723 140720
rect 228988 140662 230723 140664
rect 230657 140659 230723 140662
rect 214005 140586 214071 140589
rect 214005 140584 217028 140586
rect 214005 140528 214010 140584
rect 214066 140528 217028 140584
rect 214005 140526 217028 140528
rect 214005 140523 214071 140526
rect 281717 140450 281783 140453
rect 279956 140448 281783 140450
rect 252502 140178 252508 140180
rect 228988 140118 252508 140178
rect 252502 140116 252508 140118
rect 252572 140116 252578 140180
rect 268150 140178 268210 140420
rect 279956 140392 281722 140448
rect 281778 140392 281783 140448
rect 279956 140390 281783 140392
rect 281717 140387 281783 140390
rect 258030 140118 268210 140178
rect 213913 139906 213979 139909
rect 213913 139904 217028 139906
rect 213913 139848 213918 139904
rect 213974 139848 217028 139904
rect 213913 139846 217028 139848
rect 213913 139843 213979 139846
rect 231301 139770 231367 139773
rect 228988 139768 231367 139770
rect 228988 139712 231306 139768
rect 231362 139712 231367 139768
rect 228988 139710 231367 139712
rect 231301 139707 231367 139710
rect 237966 139708 237972 139772
rect 238036 139770 238042 139772
rect 258030 139770 258090 140118
rect 265801 140042 265867 140045
rect 265801 140040 268180 140042
rect 265801 139984 265806 140040
rect 265862 139984 268180 140040
rect 265801 139982 268180 139984
rect 265801 139979 265867 139982
rect 282269 139770 282335 139773
rect 238036 139710 258090 139770
rect 279956 139768 282335 139770
rect 279956 139712 282274 139768
rect 282330 139712 282335 139768
rect 279956 139710 282335 139712
rect 238036 139708 238042 139710
rect 282269 139707 282335 139710
rect 264973 139634 265039 139637
rect 264973 139632 268180 139634
rect 264973 139576 264978 139632
rect 265034 139576 268180 139632
rect 264973 139574 268180 139576
rect 264973 139571 265039 139574
rect 583109 139362 583175 139365
rect 583520 139362 584960 139452
rect 583109 139360 584960 139362
rect 583109 139304 583114 139360
rect 583170 139304 584960 139360
rect 583109 139302 584960 139304
rect 583109 139299 583175 139302
rect 213913 139226 213979 139229
rect 233182 139226 233188 139228
rect 213913 139224 217028 139226
rect 213913 139168 213918 139224
rect 213974 139168 217028 139224
rect 213913 139166 217028 139168
rect 228988 139166 233188 139226
rect 213913 139163 213979 139166
rect 233182 139164 233188 139166
rect 233252 139164 233258 139228
rect 583520 139212 584960 139302
rect 237598 138818 237604 138820
rect 228988 138758 237604 138818
rect 237598 138756 237604 138758
rect 237668 138756 237674 138820
rect 268150 138818 268210 139196
rect 282269 138954 282335 138957
rect 279956 138952 282335 138954
rect 279956 138896 282274 138952
rect 282330 138896 282335 138952
rect 279956 138894 282335 138896
rect 282269 138891 282335 138894
rect 258030 138758 268210 138818
rect 204989 138138 205055 138141
rect 216998 138138 217058 138652
rect 238150 138348 238156 138412
rect 238220 138410 238226 138412
rect 258030 138410 258090 138758
rect 264973 138682 265039 138685
rect 264973 138680 268180 138682
rect 264973 138624 264978 138680
rect 265034 138624 268180 138680
rect 264973 138622 268180 138624
rect 264973 138619 265039 138622
rect 238220 138350 258090 138410
rect 238220 138348 238226 138350
rect 231761 138274 231827 138277
rect 228988 138272 231827 138274
rect 228988 138216 231766 138272
rect 231822 138216 231827 138272
rect 228988 138214 231827 138216
rect 231761 138211 231827 138214
rect 262857 138274 262923 138277
rect 282821 138274 282887 138277
rect 262857 138272 268180 138274
rect 262857 138216 262862 138272
rect 262918 138216 268180 138272
rect 262857 138214 268180 138216
rect 279956 138272 282887 138274
rect 279956 138216 282826 138272
rect 282882 138216 282887 138272
rect 279956 138214 282887 138216
rect 262857 138211 262923 138214
rect 282821 138211 282887 138214
rect 204989 138136 217058 138138
rect 204989 138080 204994 138136
rect 205050 138080 217058 138136
rect 204989 138078 217058 138080
rect 204989 138075 205055 138078
rect 214741 138002 214807 138005
rect 214741 138000 217028 138002
rect 214741 137944 214746 138000
rect 214802 137944 217028 138000
rect 214741 137942 217028 137944
rect 214741 137939 214807 137942
rect 234654 137866 234660 137868
rect 228988 137806 234660 137866
rect 234654 137804 234660 137806
rect 234724 137804 234730 137868
rect 268150 137594 268210 137836
rect 258030 137534 268210 137594
rect 213913 137322 213979 137325
rect 230013 137322 230079 137325
rect 213913 137320 217028 137322
rect 213913 137264 213918 137320
rect 213974 137264 217028 137320
rect 213913 137262 217028 137264
rect 228988 137320 230079 137322
rect 228988 137264 230018 137320
rect 230074 137264 230079 137320
rect 228988 137262 230079 137264
rect 213913 137259 213979 137262
rect 230013 137259 230079 137262
rect 229737 137186 229803 137189
rect 258030 137186 258090 137534
rect 264973 137458 265039 137461
rect 281717 137458 281783 137461
rect 264973 137456 268180 137458
rect 264973 137400 264978 137456
rect 265034 137400 268180 137456
rect 264973 137398 268180 137400
rect 279956 137456 281783 137458
rect 279956 137400 281722 137456
rect 281778 137400 281783 137456
rect 279956 137398 281783 137400
rect 264973 137395 265039 137398
rect 281717 137395 281783 137398
rect 229737 137184 258090 137186
rect 229737 137128 229742 137184
rect 229798 137128 258090 137184
rect 229737 137126 258090 137128
rect 229737 137123 229803 137126
rect 258030 136990 268180 137050
rect 231577 136914 231643 136917
rect 228988 136912 231643 136914
rect -960 136778 480 136868
rect 228988 136856 231582 136912
rect 231638 136856 231643 136912
rect 228988 136854 231643 136856
rect 231577 136851 231643 136854
rect 236729 136914 236795 136917
rect 258030 136914 258090 136990
rect 236729 136912 258090 136914
rect 236729 136856 236734 136912
rect 236790 136856 258090 136912
rect 236729 136854 258090 136856
rect 236729 136851 236795 136854
rect 3509 136778 3575 136781
rect -960 136776 3575 136778
rect -960 136720 3514 136776
rect 3570 136720 3575 136776
rect -960 136718 3575 136720
rect -960 136628 480 136718
rect 3509 136715 3575 136718
rect 214005 136642 214071 136645
rect 265065 136642 265131 136645
rect 282821 136642 282887 136645
rect 214005 136640 217028 136642
rect 214005 136584 214010 136640
rect 214066 136584 217028 136640
rect 214005 136582 217028 136584
rect 265065 136640 268180 136642
rect 265065 136584 265070 136640
rect 265126 136584 268180 136640
rect 265065 136582 268180 136584
rect 279956 136640 282887 136642
rect 279956 136584 282826 136640
rect 282882 136584 282887 136640
rect 279956 136582 282887 136584
rect 214005 136579 214071 136582
rect 265065 136579 265131 136582
rect 282821 136579 282887 136582
rect 242934 136370 242940 136372
rect 228988 136310 242940 136370
rect 242934 136308 242940 136310
rect 243004 136308 243010 136372
rect 267089 136234 267155 136237
rect 267089 136232 268180 136234
rect 267089 136176 267094 136232
rect 267150 136176 268180 136232
rect 267089 136174 268180 136176
rect 267089 136171 267155 136174
rect 213913 135962 213979 135965
rect 231393 135962 231459 135965
rect 281901 135962 281967 135965
rect 213913 135960 217028 135962
rect 213913 135904 213918 135960
rect 213974 135904 217028 135960
rect 213913 135902 217028 135904
rect 228988 135960 231459 135962
rect 228988 135904 231398 135960
rect 231454 135904 231459 135960
rect 228988 135902 231459 135904
rect 279956 135960 281967 135962
rect 279956 135904 281906 135960
rect 281962 135904 281967 135960
rect 279956 135902 281967 135904
rect 213913 135899 213979 135902
rect 231393 135899 231459 135902
rect 281901 135899 281967 135902
rect 262949 135690 263015 135693
rect 262949 135688 268180 135690
rect 262949 135632 262954 135688
rect 263010 135632 268180 135688
rect 262949 135630 268180 135632
rect 262949 135627 263015 135630
rect 230933 135418 230999 135421
rect 228988 135416 230999 135418
rect 228988 135360 230938 135416
rect 230994 135360 230999 135416
rect 228988 135358 230999 135360
rect 230933 135355 230999 135358
rect 167637 135282 167703 135285
rect 265893 135282 265959 135285
rect 167637 135280 217028 135282
rect 167637 135224 167642 135280
rect 167698 135224 217028 135280
rect 167637 135222 217028 135224
rect 265893 135280 268180 135282
rect 265893 135224 265898 135280
rect 265954 135224 268180 135280
rect 265893 135222 268180 135224
rect 167637 135219 167703 135222
rect 265893 135219 265959 135222
rect 283782 135146 283788 135148
rect 279956 135086 283788 135146
rect 283782 135084 283788 135086
rect 283852 135084 283858 135148
rect 231761 135010 231827 135013
rect 228988 135008 231827 135010
rect 228988 134952 231766 135008
rect 231822 134952 231827 135008
rect 228988 134950 231827 134952
rect 231761 134947 231827 134950
rect 199377 134194 199443 134197
rect 216998 134194 217058 134572
rect 260046 134540 260052 134604
rect 260116 134602 260122 134604
rect 268150 134602 268210 134844
rect 260116 134542 268210 134602
rect 260116 134540 260122 134542
rect 231669 134466 231735 134469
rect 228988 134464 231735 134466
rect 228988 134408 231674 134464
rect 231730 134408 231735 134464
rect 228988 134406 231735 134408
rect 231669 134403 231735 134406
rect 246573 134466 246639 134469
rect 265341 134466 265407 134469
rect 246573 134464 265407 134466
rect 246573 134408 246578 134464
rect 246634 134408 265346 134464
rect 265402 134408 265407 134464
rect 246573 134406 265407 134408
rect 246573 134403 246639 134406
rect 265341 134403 265407 134406
rect 265617 134466 265683 134469
rect 282085 134466 282151 134469
rect 265617 134464 268180 134466
rect 265617 134408 265622 134464
rect 265678 134408 268180 134464
rect 265617 134406 268180 134408
rect 279956 134464 282151 134466
rect 279956 134408 282090 134464
rect 282146 134408 282151 134464
rect 279956 134406 282151 134408
rect 265617 134403 265683 134406
rect 282085 134403 282151 134406
rect 199377 134192 217058 134194
rect 199377 134136 199382 134192
rect 199438 134136 217058 134192
rect 199377 134134 217058 134136
rect 199377 134131 199443 134134
rect 231485 134058 231551 134061
rect 228988 134056 231551 134058
rect 228988 134000 231490 134056
rect 231546 134000 231551 134056
rect 228988 133998 231551 134000
rect 231485 133995 231551 133998
rect 264973 134058 265039 134061
rect 264973 134056 268180 134058
rect 264973 134000 264978 134056
rect 265034 134000 268180 134056
rect 264973 133998 268180 134000
rect 264973 133995 265039 133998
rect 213913 133922 213979 133925
rect 213913 133920 217028 133922
rect 213913 133864 213918 133920
rect 213974 133864 217028 133920
rect 213913 133862 217028 133864
rect 213913 133859 213979 133862
rect 250529 133650 250595 133653
rect 238710 133648 250595 133650
rect 238710 133592 250534 133648
rect 250590 133592 250595 133648
rect 238710 133590 250595 133592
rect 232865 133514 232931 133517
rect 228988 133512 232931 133514
rect 228988 133456 232870 133512
rect 232926 133456 232931 133512
rect 228988 133454 232931 133456
rect 232865 133451 232931 133454
rect 178534 133044 178540 133108
rect 178604 133106 178610 133108
rect 198089 133106 198155 133109
rect 178604 133104 198155 133106
rect 178604 133048 198094 133104
rect 198150 133048 198155 133104
rect 178604 133046 198155 133048
rect 178604 133044 178610 133046
rect 198089 133043 198155 133046
rect 166206 132772 166212 132836
rect 166276 132834 166282 132836
rect 216998 132834 217058 133348
rect 238710 133106 238770 133590
rect 250529 133587 250595 133590
rect 265065 133650 265131 133653
rect 282821 133650 282887 133653
rect 265065 133648 268180 133650
rect 265065 133592 265070 133648
rect 265126 133592 268180 133648
rect 265065 133590 268180 133592
rect 279956 133648 282887 133650
rect 279956 133592 282826 133648
rect 282882 133592 282887 133648
rect 279956 133590 282887 133592
rect 265065 133587 265131 133590
rect 282821 133587 282887 133590
rect 228988 133046 238770 133106
rect 264973 133106 265039 133109
rect 264973 133104 268180 133106
rect 264973 133048 264978 133104
rect 265034 133048 268180 133104
rect 264973 133046 268180 133048
rect 264973 133043 265039 133046
rect 282269 132834 282335 132837
rect 166276 132774 217058 132834
rect 279956 132832 282335 132834
rect 279956 132776 282274 132832
rect 282330 132776 282335 132832
rect 279956 132774 282335 132776
rect 166276 132772 166282 132774
rect 282269 132771 282335 132774
rect 213913 132698 213979 132701
rect 213913 132696 217028 132698
rect 213913 132640 213918 132696
rect 213974 132640 217028 132696
rect 213913 132638 217028 132640
rect 258030 132638 268180 132698
rect 213913 132635 213979 132638
rect 231669 132562 231735 132565
rect 228988 132560 231735 132562
rect 228988 132504 231674 132560
rect 231730 132504 231735 132560
rect 228988 132502 231735 132504
rect 231669 132499 231735 132502
rect 249057 132562 249123 132565
rect 258030 132562 258090 132638
rect 249057 132560 258090 132562
rect 249057 132504 249062 132560
rect 249118 132504 258090 132560
rect 249057 132502 258090 132504
rect 249057 132499 249123 132502
rect 231761 132154 231827 132157
rect 228988 132152 231827 132154
rect 228988 132096 231766 132152
rect 231822 132096 231827 132152
rect 228988 132094 231827 132096
rect 231761 132091 231827 132094
rect 213913 132018 213979 132021
rect 229829 132018 229895 132021
rect 268150 132018 268210 132260
rect 282821 132154 282887 132157
rect 279956 132152 282887 132154
rect 279956 132096 282826 132152
rect 282882 132096 282887 132152
rect 279956 132094 282887 132096
rect 282821 132091 282887 132094
rect 213913 132016 217028 132018
rect 213913 131960 213918 132016
rect 213974 131960 217028 132016
rect 213913 131958 217028 131960
rect 229829 132016 268210 132018
rect 229829 131960 229834 132016
rect 229890 131960 268210 132016
rect 229829 131958 268210 131960
rect 213913 131955 213979 131958
rect 229829 131955 229895 131958
rect 264973 131882 265039 131885
rect 264973 131880 268180 131882
rect 264973 131824 264978 131880
rect 265034 131824 268180 131880
rect 264973 131822 268180 131824
rect 264973 131819 265039 131822
rect 230974 131610 230980 131612
rect 228988 131550 230980 131610
rect 230974 131548 230980 131550
rect 231044 131548 231050 131612
rect 265065 131474 265131 131477
rect 265065 131472 268180 131474
rect 265065 131416 265070 131472
rect 265126 131416 268180 131472
rect 265065 131414 268180 131416
rect 265065 131411 265131 131414
rect 214557 131338 214623 131341
rect 282729 131338 282795 131341
rect 214557 131336 217028 131338
rect 214557 131280 214562 131336
rect 214618 131280 217028 131336
rect 214557 131278 217028 131280
rect 279956 131336 282795 131338
rect 279956 131280 282734 131336
rect 282790 131280 282795 131336
rect 279956 131278 282795 131280
rect 214557 131275 214623 131278
rect 282729 131275 282795 131278
rect 231117 131202 231183 131205
rect 228988 131200 231183 131202
rect 228988 131144 231122 131200
rect 231178 131144 231183 131200
rect 228988 131142 231183 131144
rect 231117 131139 231183 131142
rect 262806 131004 262812 131068
rect 262876 131066 262882 131068
rect 262876 131006 268180 131066
rect 262876 131004 262882 131006
rect 214005 130658 214071 130661
rect 231209 130658 231275 130661
rect 282269 130658 282335 130661
rect 214005 130656 217028 130658
rect 214005 130600 214010 130656
rect 214066 130600 217028 130656
rect 214005 130598 217028 130600
rect 228988 130656 231275 130658
rect 228988 130600 231214 130656
rect 231270 130600 231275 130656
rect 228988 130598 231275 130600
rect 279956 130656 282335 130658
rect 279956 130600 282274 130656
rect 282330 130600 282335 130656
rect 279956 130598 282335 130600
rect 214005 130595 214071 130598
rect 231209 130595 231275 130598
rect 282269 130595 282335 130598
rect 264973 130522 265039 130525
rect 264973 130520 268180 130522
rect 264973 130464 264978 130520
rect 265034 130464 268180 130520
rect 264973 130462 268180 130464
rect 264973 130459 265039 130462
rect 231761 130250 231827 130253
rect 228988 130248 231827 130250
rect 228988 130192 231766 130248
rect 231822 130192 231827 130248
rect 228988 130190 231827 130192
rect 231761 130187 231827 130190
rect 238109 130114 238175 130117
rect 238109 130112 268180 130114
rect 238109 130056 238114 130112
rect 238170 130056 268180 130112
rect 238109 130054 268180 130056
rect 238109 130051 238175 130054
rect 213913 129978 213979 129981
rect 213913 129976 217028 129978
rect 213913 129920 213918 129976
rect 213974 129920 217028 129976
rect 213913 129918 217028 129920
rect 213913 129915 213979 129918
rect 230565 129842 230631 129845
rect 281533 129842 281599 129845
rect 228988 129840 230631 129842
rect 228988 129784 230570 129840
rect 230626 129784 230631 129840
rect 228988 129782 230631 129784
rect 279956 129840 281599 129842
rect 279956 129784 281538 129840
rect 281594 129784 281599 129840
rect 279956 129782 281599 129784
rect 230565 129779 230631 129782
rect 281533 129779 281599 129782
rect 264973 129706 265039 129709
rect 264973 129704 268180 129706
rect 264973 129648 264978 129704
rect 265034 129648 268180 129704
rect 264973 129646 268180 129648
rect 264973 129643 265039 129646
rect 67449 129298 67515 129301
rect 68142 129298 68816 129304
rect 67449 129296 68816 129298
rect 67449 129240 67454 129296
rect 67510 129244 68816 129296
rect 214005 129298 214071 129301
rect 231761 129298 231827 129301
rect 214005 129296 217028 129298
rect 67510 129240 68202 129244
rect 67449 129238 68202 129240
rect 214005 129240 214010 129296
rect 214066 129240 217028 129296
rect 214005 129238 217028 129240
rect 228988 129296 231827 129298
rect 228988 129240 231766 129296
rect 231822 129240 231827 129296
rect 228988 129238 231827 129240
rect 67449 129235 67515 129238
rect 214005 129235 214071 129238
rect 231761 129235 231827 129238
rect 266854 129236 266860 129300
rect 266924 129298 266930 129300
rect 266924 129238 268180 129298
rect 266924 129236 266930 129238
rect 231301 129026 231367 129029
rect 251817 129026 251883 129029
rect 282085 129026 282151 129029
rect 231301 129024 251883 129026
rect 231301 128968 231306 129024
rect 231362 128968 251822 129024
rect 251878 128968 251883 129024
rect 231301 128966 251883 128968
rect 279956 129024 282151 129026
rect 279956 128968 282090 129024
rect 282146 128968 282151 129024
rect 279956 128966 282151 128968
rect 231301 128963 231367 128966
rect 251817 128963 251883 128966
rect 282085 128963 282151 128966
rect 230749 128890 230815 128893
rect 228988 128888 230815 128890
rect 228988 128832 230754 128888
rect 230810 128832 230815 128888
rect 228988 128830 230815 128832
rect 230749 128827 230815 128830
rect 258030 128830 268180 128890
rect 213913 128754 213979 128757
rect 213913 128752 217028 128754
rect 213913 128696 213918 128752
rect 213974 128696 217028 128752
rect 213913 128694 217028 128696
rect 213913 128691 213979 128694
rect 253054 128692 253060 128756
rect 253124 128754 253130 128756
rect 258030 128754 258090 128830
rect 253124 128694 258090 128754
rect 253124 128692 253130 128694
rect 267774 128420 267780 128484
rect 267844 128482 267850 128484
rect 267844 128422 268180 128482
rect 267844 128420 267850 128422
rect 253197 128346 253263 128349
rect 282821 128346 282887 128349
rect 228988 128344 253263 128346
rect 228988 128288 253202 128344
rect 253258 128288 253263 128344
rect 228988 128286 253263 128288
rect 279956 128344 282887 128346
rect 279956 128288 282826 128344
rect 282882 128288 282887 128344
rect 279956 128286 282887 128288
rect 253197 128283 253263 128286
rect 282821 128283 282887 128286
rect 65333 128074 65399 128077
rect 68142 128074 68816 128080
rect 65333 128072 68816 128074
rect 65333 128016 65338 128072
rect 65394 128020 68816 128072
rect 214005 128074 214071 128077
rect 214005 128072 217028 128074
rect 65394 128016 68202 128020
rect 65333 128014 68202 128016
rect 214005 128016 214010 128072
rect 214066 128016 217028 128072
rect 214005 128014 217028 128016
rect 65333 128011 65399 128014
rect 214005 128011 214071 128014
rect 231761 127938 231827 127941
rect 228988 127936 231827 127938
rect 228988 127880 231766 127936
rect 231822 127880 231827 127936
rect 228988 127878 231827 127880
rect 231761 127875 231827 127878
rect 264094 127876 264100 127940
rect 264164 127938 264170 127940
rect 264164 127878 268180 127938
rect 264164 127876 264170 127878
rect 264973 127530 265039 127533
rect 282729 127530 282795 127533
rect 264973 127528 268180 127530
rect 264973 127472 264978 127528
rect 265034 127472 268180 127528
rect 264973 127470 268180 127472
rect 279956 127528 282795 127530
rect 279956 127472 282734 127528
rect 282790 127472 282795 127528
rect 279956 127470 282795 127472
rect 264973 127467 265039 127470
rect 282729 127467 282795 127470
rect 213913 127394 213979 127397
rect 231117 127394 231183 127397
rect 213913 127392 217028 127394
rect 213913 127336 213918 127392
rect 213974 127336 217028 127392
rect 213913 127334 217028 127336
rect 228988 127392 231183 127394
rect 228988 127336 231122 127392
rect 231178 127336 231183 127392
rect 228988 127334 231183 127336
rect 213913 127331 213979 127334
rect 231117 127331 231183 127334
rect 64781 127122 64847 127125
rect 65333 127122 65399 127125
rect 64781 127120 65399 127122
rect 64781 127064 64786 127120
rect 64842 127064 65338 127120
rect 65394 127064 65399 127120
rect 64781 127062 65399 127064
rect 64781 127059 64847 127062
rect 65333 127059 65399 127062
rect 258574 127060 258580 127124
rect 258644 127122 258650 127124
rect 258644 127062 268180 127122
rect 258644 127060 258650 127062
rect 231761 126986 231827 126989
rect 228988 126984 231827 126986
rect 228988 126928 231766 126984
rect 231822 126928 231827 126984
rect 228988 126926 231827 126928
rect 231761 126923 231827 126926
rect 280102 126850 280108 126852
rect 279956 126790 280108 126850
rect 280102 126788 280108 126790
rect 280172 126788 280178 126852
rect 214005 126714 214071 126717
rect 214005 126712 217028 126714
rect 214005 126656 214010 126712
rect 214066 126656 217028 126712
rect 214005 126654 217028 126656
rect 258030 126654 268180 126714
rect 214005 126651 214071 126654
rect 230974 126516 230980 126580
rect 231044 126578 231050 126580
rect 258030 126578 258090 126654
rect 231044 126518 258090 126578
rect 231044 126516 231050 126518
rect 230933 126442 230999 126445
rect 228988 126440 230999 126442
rect 228988 126384 230938 126440
rect 230994 126384 230999 126440
rect 228988 126382 230999 126384
rect 230933 126379 230999 126382
rect 67541 126306 67607 126309
rect 68142 126306 68816 126312
rect 67541 126304 68816 126306
rect 67541 126248 67546 126304
rect 67602 126252 68816 126304
rect 264973 126306 265039 126309
rect 264973 126304 268180 126306
rect 67602 126248 68202 126252
rect 67541 126246 68202 126248
rect 264973 126248 264978 126304
rect 265034 126248 268180 126304
rect 264973 126246 268180 126248
rect 67541 126243 67607 126246
rect 264973 126243 265039 126246
rect 213913 126034 213979 126037
rect 231209 126034 231275 126037
rect 282269 126034 282335 126037
rect 213913 126032 217028 126034
rect 213913 125976 213918 126032
rect 213974 125976 217028 126032
rect 213913 125974 217028 125976
rect 228988 126032 231275 126034
rect 228988 125976 231214 126032
rect 231270 125976 231275 126032
rect 228988 125974 231275 125976
rect 279956 126032 282335 126034
rect 279956 125976 282274 126032
rect 282330 125976 282335 126032
rect 279956 125974 282335 125976
rect 213913 125971 213979 125974
rect 231209 125971 231275 125974
rect 282269 125971 282335 125974
rect 580901 126034 580967 126037
rect 583520 126034 584960 126124
rect 580901 126032 584960 126034
rect 580901 125976 580906 126032
rect 580962 125976 584960 126032
rect 580901 125974 584960 125976
rect 580901 125971 580967 125974
rect 265709 125898 265775 125901
rect 265709 125896 268180 125898
rect 265709 125840 265714 125896
rect 265770 125840 268180 125896
rect 583520 125884 584960 125974
rect 265709 125838 268180 125840
rect 265709 125835 265775 125838
rect 231301 125490 231367 125493
rect 228988 125488 231367 125490
rect 228988 125432 231306 125488
rect 231362 125432 231367 125488
rect 228988 125430 231367 125432
rect 231301 125427 231367 125430
rect 213913 125354 213979 125357
rect 264605 125354 264671 125357
rect 213913 125352 217028 125354
rect 213913 125296 213918 125352
rect 213974 125296 217028 125352
rect 213913 125294 217028 125296
rect 264605 125352 268180 125354
rect 264605 125296 264610 125352
rect 264666 125296 268180 125352
rect 264605 125294 268180 125296
rect 213913 125291 213979 125294
rect 264605 125291 264671 125294
rect 66161 125218 66227 125221
rect 68142 125218 68816 125224
rect 282085 125218 282151 125221
rect 66161 125216 68816 125218
rect 66161 125160 66166 125216
rect 66222 125164 68816 125216
rect 279956 125216 282151 125218
rect 66222 125160 68202 125164
rect 66161 125158 68202 125160
rect 279956 125160 282090 125216
rect 282146 125160 282151 125216
rect 279956 125158 282151 125160
rect 66161 125155 66227 125158
rect 282085 125155 282151 125158
rect 236637 125082 236703 125085
rect 228988 125080 236703 125082
rect 228988 125024 236642 125080
rect 236698 125024 236703 125080
rect 228988 125022 236703 125024
rect 236637 125019 236703 125022
rect 264973 124946 265039 124949
rect 264973 124944 268180 124946
rect 264973 124888 264978 124944
rect 265034 124888 268180 124944
rect 264973 124886 268180 124888
rect 264973 124883 265039 124886
rect 231117 124810 231183 124813
rect 257521 124810 257587 124813
rect 231117 124808 257587 124810
rect 231117 124752 231122 124808
rect 231178 124752 257526 124808
rect 257582 124752 257587 124808
rect 231117 124750 257587 124752
rect 231117 124747 231183 124750
rect 257521 124747 257587 124750
rect 214925 124674 214991 124677
rect 214925 124672 217028 124674
rect 214925 124616 214930 124672
rect 214986 124616 217028 124672
rect 214925 124614 217028 124616
rect 214925 124611 214991 124614
rect 230473 124538 230539 124541
rect 228988 124536 230539 124538
rect 228988 124480 230478 124536
rect 230534 124480 230539 124536
rect 228988 124478 230539 124480
rect 230473 124475 230539 124478
rect 239397 124538 239463 124541
rect 282821 124538 282887 124541
rect 239397 124536 268180 124538
rect 239397 124480 239402 124536
rect 239458 124480 268180 124536
rect 239397 124478 268180 124480
rect 279956 124536 282887 124538
rect 279956 124480 282826 124536
rect 282882 124480 282887 124536
rect 279956 124478 282887 124480
rect 239397 124475 239463 124478
rect 282821 124475 282887 124478
rect 213913 124130 213979 124133
rect 231761 124130 231827 124133
rect 213913 124128 217028 124130
rect 213913 124072 213918 124128
rect 213974 124072 217028 124128
rect 213913 124070 217028 124072
rect 228988 124128 231827 124130
rect 228988 124072 231766 124128
rect 231822 124072 231827 124128
rect 228988 124070 231827 124072
rect 213913 124067 213979 124070
rect 231761 124067 231827 124070
rect 264973 124130 265039 124133
rect 264973 124128 268180 124130
rect 264973 124072 264978 124128
rect 265034 124072 268180 124128
rect 264973 124070 268180 124072
rect 264973 124067 265039 124070
rect -960 123572 480 123812
rect 282269 123722 282335 123725
rect 258030 123662 268180 123722
rect 279956 123720 282335 123722
rect 279956 123664 282274 123720
rect 282330 123664 282335 123720
rect 279956 123662 282335 123664
rect 67357 123586 67423 123589
rect 68142 123586 68816 123592
rect 231158 123586 231164 123588
rect 67357 123584 68816 123586
rect 67357 123528 67362 123584
rect 67418 123532 68816 123584
rect 67418 123528 68202 123532
rect 67357 123526 68202 123528
rect 228988 123526 231164 123586
rect 67357 123523 67423 123526
rect 231158 123524 231164 123526
rect 231228 123524 231234 123588
rect 247953 123586 248019 123589
rect 258030 123586 258090 123662
rect 282269 123659 282335 123662
rect 247953 123584 258090 123586
rect 247953 123528 247958 123584
rect 248014 123528 258090 123584
rect 247953 123526 258090 123528
rect 247953 123523 248019 123526
rect 198273 123450 198339 123453
rect 213361 123450 213427 123453
rect 198273 123448 213427 123450
rect 198273 123392 198278 123448
rect 198334 123392 213366 123448
rect 213422 123392 213427 123448
rect 198273 123390 213427 123392
rect 198273 123387 198339 123390
rect 213361 123387 213427 123390
rect 214005 123450 214071 123453
rect 234245 123450 234311 123453
rect 254577 123450 254643 123453
rect 214005 123448 217028 123450
rect 214005 123392 214010 123448
rect 214066 123392 217028 123448
rect 214005 123390 217028 123392
rect 234245 123448 254643 123450
rect 234245 123392 234250 123448
rect 234306 123392 254582 123448
rect 254638 123392 254643 123448
rect 234245 123390 254643 123392
rect 214005 123387 214071 123390
rect 234245 123387 234311 123390
rect 254577 123387 254643 123390
rect 265065 123314 265131 123317
rect 265065 123312 268180 123314
rect 265065 123256 265070 123312
rect 265126 123256 268180 123312
rect 265065 123254 268180 123256
rect 265065 123251 265131 123254
rect 231393 123178 231459 123181
rect 228988 123176 231459 123178
rect 228988 123120 231398 123176
rect 231454 123120 231459 123176
rect 228988 123118 231459 123120
rect 231393 123115 231459 123118
rect 282821 123042 282887 123045
rect 279956 123040 282887 123042
rect 279956 122984 282826 123040
rect 282882 122984 282887 123040
rect 279956 122982 282887 122984
rect 282821 122979 282887 122982
rect 266997 122906 267063 122909
rect 266997 122904 268180 122906
rect 266997 122848 267002 122904
rect 267058 122848 268180 122904
rect 266997 122846 268180 122848
rect 266997 122843 267063 122846
rect 214005 122770 214071 122773
rect 214005 122768 217028 122770
rect 214005 122712 214010 122768
rect 214066 122712 217028 122768
rect 214005 122710 217028 122712
rect 214005 122707 214071 122710
rect 66069 122634 66135 122637
rect 68142 122634 68816 122640
rect 235533 122634 235599 122637
rect 66069 122632 68816 122634
rect 66069 122576 66074 122632
rect 66130 122580 68816 122632
rect 228988 122632 235599 122634
rect 66130 122576 68202 122580
rect 66069 122574 68202 122576
rect 228988 122576 235538 122632
rect 235594 122576 235599 122632
rect 228988 122574 235599 122576
rect 66069 122571 66135 122574
rect 235533 122571 235599 122574
rect 264973 122362 265039 122365
rect 264973 122360 268180 122362
rect 264973 122304 264978 122360
rect 265034 122304 268180 122360
rect 264973 122302 268180 122304
rect 264973 122299 265039 122302
rect 231761 122226 231827 122229
rect 282453 122226 282519 122229
rect 228988 122224 231827 122226
rect 228988 122168 231766 122224
rect 231822 122168 231827 122224
rect 228988 122166 231827 122168
rect 279956 122224 282519 122226
rect 279956 122168 282458 122224
rect 282514 122168 282519 122224
rect 279956 122166 282519 122168
rect 231761 122163 231827 122166
rect 282453 122163 282519 122166
rect 213913 122090 213979 122093
rect 213913 122088 217028 122090
rect 213913 122032 213918 122088
rect 213974 122032 217028 122088
rect 213913 122030 217028 122032
rect 213913 122027 213979 122030
rect 258030 121894 268180 121954
rect 230013 121818 230079 121821
rect 258030 121818 258090 121894
rect 230013 121816 258090 121818
rect 230013 121760 230018 121816
rect 230074 121760 258090 121816
rect 230013 121758 258090 121760
rect 230013 121755 230079 121758
rect 231485 121682 231551 121685
rect 228988 121680 231551 121682
rect 228988 121624 231490 121680
rect 231546 121624 231551 121680
rect 228988 121622 231551 121624
rect 231485 121619 231551 121622
rect 260097 121682 260163 121685
rect 260097 121680 268210 121682
rect 260097 121624 260102 121680
rect 260158 121624 268210 121680
rect 260097 121622 268210 121624
rect 260097 121619 260163 121622
rect 268150 121516 268210 121622
rect 213913 121410 213979 121413
rect 282821 121410 282887 121413
rect 213913 121408 217028 121410
rect 213913 121352 213918 121408
rect 213974 121352 217028 121408
rect 213913 121350 217028 121352
rect 279956 121408 282887 121410
rect 279956 121352 282826 121408
rect 282882 121352 282887 121408
rect 279956 121350 282887 121352
rect 213913 121347 213979 121350
rect 282821 121347 282887 121350
rect 231761 121274 231827 121277
rect 228988 121272 231827 121274
rect 228988 121216 231766 121272
rect 231822 121216 231827 121272
rect 228988 121214 231827 121216
rect 231761 121211 231827 121214
rect 264973 121138 265039 121141
rect 264973 121136 268180 121138
rect 264973 121080 264978 121136
rect 265034 121080 268180 121136
rect 264973 121078 268180 121080
rect 264973 121075 265039 121078
rect 65885 120866 65951 120869
rect 68142 120866 68816 120872
rect 65885 120864 68816 120866
rect 65885 120808 65890 120864
rect 65946 120812 68816 120864
rect 65946 120808 68202 120812
rect 65885 120806 68202 120808
rect 65885 120803 65951 120806
rect 216121 120730 216187 120733
rect 231209 120730 231275 120733
rect 216121 120728 217028 120730
rect 216121 120672 216126 120728
rect 216182 120672 217028 120728
rect 216121 120670 217028 120672
rect 228988 120728 231275 120730
rect 228988 120672 231214 120728
rect 231270 120672 231275 120728
rect 228988 120670 231275 120672
rect 216121 120667 216187 120670
rect 231209 120667 231275 120670
rect 235533 120730 235599 120733
rect 262121 120730 262187 120733
rect 235533 120728 262187 120730
rect 235533 120672 235538 120728
rect 235594 120672 262126 120728
rect 262182 120672 262187 120728
rect 235533 120670 262187 120672
rect 235533 120667 235599 120670
rect 262121 120667 262187 120670
rect 267273 120730 267339 120733
rect 280286 120730 280292 120732
rect 267273 120728 268180 120730
rect 267273 120672 267278 120728
rect 267334 120672 268180 120728
rect 267273 120670 268180 120672
rect 279956 120670 280292 120730
rect 267273 120667 267339 120670
rect 280286 120668 280292 120670
rect 280356 120668 280362 120732
rect 230657 120322 230723 120325
rect 228988 120320 230723 120322
rect 228988 120264 230662 120320
rect 230718 120264 230723 120320
rect 228988 120262 230723 120264
rect 230657 120259 230723 120262
rect 258030 120262 268180 120322
rect 64689 120186 64755 120189
rect 65885 120186 65951 120189
rect 64689 120184 65951 120186
rect 64689 120128 64694 120184
rect 64750 120128 65890 120184
rect 65946 120128 65951 120184
rect 64689 120126 65951 120128
rect 64689 120123 64755 120126
rect 65885 120123 65951 120126
rect 236637 120186 236703 120189
rect 258030 120186 258090 120262
rect 236637 120184 258090 120186
rect 236637 120128 236642 120184
rect 236698 120128 258090 120184
rect 236637 120126 258090 120128
rect 236637 120123 236703 120126
rect 214005 120050 214071 120053
rect 231761 120050 231827 120053
rect 246389 120050 246455 120053
rect 214005 120048 217028 120050
rect 214005 119992 214010 120048
rect 214066 119992 217028 120048
rect 214005 119990 217028 119992
rect 231761 120048 246455 120050
rect 231761 119992 231766 120048
rect 231822 119992 246394 120048
rect 246450 119992 246455 120048
rect 231761 119990 246455 119992
rect 214005 119987 214071 119990
rect 231761 119987 231827 119990
rect 246389 119987 246455 119990
rect 282637 119914 282703 119917
rect 279956 119912 282703 119914
rect 279956 119856 282642 119912
rect 282698 119856 282703 119912
rect 279956 119854 282703 119856
rect 282637 119851 282703 119854
rect 243629 119778 243695 119781
rect 228988 119776 243695 119778
rect 228988 119720 243634 119776
rect 243690 119720 243695 119776
rect 228988 119718 243695 119720
rect 243629 119715 243695 119718
rect 213913 119506 213979 119509
rect 262305 119506 262371 119509
rect 268150 119506 268210 119748
rect 213913 119504 217028 119506
rect 213913 119448 213918 119504
rect 213974 119448 217028 119504
rect 213913 119446 217028 119448
rect 262305 119504 268210 119506
rect 262305 119448 262310 119504
rect 262366 119448 268210 119504
rect 262305 119446 268210 119448
rect 213913 119443 213979 119446
rect 262305 119443 262371 119446
rect 231761 119370 231827 119373
rect 228988 119368 231827 119370
rect 228988 119312 231766 119368
rect 231822 119312 231827 119368
rect 228988 119310 231827 119312
rect 231761 119307 231827 119310
rect 258030 119310 268180 119370
rect 250294 119172 250300 119236
rect 250364 119234 250370 119236
rect 258030 119234 258090 119310
rect 282085 119234 282151 119237
rect 250364 119174 258090 119234
rect 279956 119232 282151 119234
rect 279956 119176 282090 119232
rect 282146 119176 282151 119232
rect 279956 119174 282151 119176
rect 250364 119172 250370 119174
rect 282085 119171 282151 119174
rect 240726 119036 240732 119100
rect 240796 119098 240802 119100
rect 262305 119098 262371 119101
rect 240796 119096 262371 119098
rect 240796 119040 262310 119096
rect 262366 119040 262371 119096
rect 240796 119038 262371 119040
rect 240796 119036 240802 119038
rect 262305 119035 262371 119038
rect 231485 118962 231551 118965
rect 228988 118960 231551 118962
rect 228988 118904 231490 118960
rect 231546 118904 231551 118960
rect 228988 118902 231551 118904
rect 231485 118899 231551 118902
rect 264237 118962 264303 118965
rect 264237 118960 268180 118962
rect 264237 118904 264242 118960
rect 264298 118904 268180 118960
rect 264237 118902 268180 118904
rect 264237 118899 264303 118902
rect 193949 118826 194015 118829
rect 193949 118824 217028 118826
rect 193949 118768 193954 118824
rect 194010 118768 217028 118824
rect 193949 118766 217028 118768
rect 193949 118763 194015 118766
rect 265065 118554 265131 118557
rect 265065 118552 268180 118554
rect 265065 118496 265070 118552
rect 265126 118496 268180 118552
rect 265065 118494 268180 118496
rect 265065 118491 265131 118494
rect 217225 118418 217291 118421
rect 233734 118418 233740 118420
rect 200070 118416 217291 118418
rect 200070 118360 217230 118416
rect 217286 118360 217291 118416
rect 200070 118358 217291 118360
rect 228988 118358 233740 118418
rect 191189 118282 191255 118285
rect 200070 118282 200130 118358
rect 217225 118355 217291 118358
rect 233734 118356 233740 118358
rect 233804 118356 233810 118420
rect 281809 118418 281875 118421
rect 279956 118416 281875 118418
rect 279956 118360 281814 118416
rect 281870 118360 281875 118416
rect 279956 118358 281875 118360
rect 281809 118355 281875 118358
rect 191189 118280 200130 118282
rect 191189 118224 191194 118280
rect 191250 118224 200130 118280
rect 191189 118222 200130 118224
rect 191189 118219 191255 118222
rect 214005 118146 214071 118149
rect 264973 118146 265039 118149
rect 214005 118144 217028 118146
rect 214005 118088 214010 118144
rect 214066 118088 217028 118144
rect 214005 118086 217028 118088
rect 264973 118144 268180 118146
rect 264973 118088 264978 118144
rect 265034 118088 268180 118144
rect 264973 118086 268180 118088
rect 214005 118083 214071 118086
rect 264973 118083 265039 118086
rect 230933 118010 230999 118013
rect 228988 118008 230999 118010
rect 228988 117952 230938 118008
rect 230994 117952 230999 118008
rect 228988 117950 230999 117952
rect 230933 117947 230999 117950
rect 231669 118010 231735 118013
rect 242341 118010 242407 118013
rect 231669 118008 242407 118010
rect 231669 117952 231674 118008
rect 231730 117952 242346 118008
rect 242402 117952 242407 118008
rect 231669 117950 242407 117952
rect 231669 117947 231735 117950
rect 242341 117947 242407 117950
rect 258030 117678 268180 117738
rect 251817 117602 251883 117605
rect 258030 117602 258090 117678
rect 280245 117602 280311 117605
rect 251817 117600 258090 117602
rect 251817 117544 251822 117600
rect 251878 117544 258090 117600
rect 251817 117542 258090 117544
rect 279956 117600 280311 117602
rect 279956 117544 280250 117600
rect 280306 117544 280311 117600
rect 279956 117542 280311 117544
rect 251817 117539 251883 117542
rect 280245 117539 280311 117542
rect 213913 117466 213979 117469
rect 231577 117466 231643 117469
rect 213913 117464 217028 117466
rect 213913 117408 213918 117464
rect 213974 117408 217028 117464
rect 213913 117406 217028 117408
rect 228988 117464 231643 117466
rect 228988 117408 231582 117464
rect 231638 117408 231643 117464
rect 228988 117406 231643 117408
rect 213913 117403 213979 117406
rect 231577 117403 231643 117406
rect 264973 117194 265039 117197
rect 264973 117192 268180 117194
rect 264973 117136 264978 117192
rect 265034 117136 268180 117192
rect 264973 117134 268180 117136
rect 264973 117131 265039 117134
rect 231761 117058 231827 117061
rect 228988 117056 231827 117058
rect 228988 117000 231766 117056
rect 231822 117000 231827 117056
rect 228988 116998 231827 117000
rect 231761 116995 231827 116998
rect 238017 116922 238083 116925
rect 262213 116922 262279 116925
rect 282821 116922 282887 116925
rect 238017 116920 262279 116922
rect 238017 116864 238022 116920
rect 238078 116864 262218 116920
rect 262274 116864 262279 116920
rect 238017 116862 262279 116864
rect 279956 116920 282887 116922
rect 279956 116864 282826 116920
rect 282882 116864 282887 116920
rect 279956 116862 282887 116864
rect 238017 116859 238083 116862
rect 262213 116859 262279 116862
rect 282821 116859 282887 116862
rect 214005 116786 214071 116789
rect 214005 116784 217028 116786
rect 214005 116728 214010 116784
rect 214066 116728 217028 116784
rect 214005 116726 217028 116728
rect 214005 116723 214071 116726
rect 171869 116514 171935 116517
rect 207749 116514 207815 116517
rect 231485 116514 231551 116517
rect 171869 116512 207815 116514
rect 171869 116456 171874 116512
rect 171930 116456 207754 116512
rect 207810 116456 207815 116512
rect 171869 116454 207815 116456
rect 228988 116512 231551 116514
rect 228988 116456 231490 116512
rect 231546 116456 231551 116512
rect 228988 116454 231551 116456
rect 171869 116451 171935 116454
rect 207749 116451 207815 116454
rect 231485 116451 231551 116454
rect 232773 116514 232839 116517
rect 268150 116514 268210 116756
rect 232773 116512 268210 116514
rect 232773 116456 232778 116512
rect 232834 116456 268210 116512
rect 232773 116454 268210 116456
rect 232773 116451 232839 116454
rect 265065 116378 265131 116381
rect 265065 116376 268180 116378
rect 265065 116320 265070 116376
rect 265126 116320 268180 116376
rect 265065 116318 268180 116320
rect 265065 116315 265131 116318
rect 213913 116106 213979 116109
rect 230749 116106 230815 116109
rect 213913 116104 217028 116106
rect 213913 116048 213918 116104
rect 213974 116048 217028 116104
rect 213913 116046 217028 116048
rect 228988 116104 230815 116106
rect 228988 116048 230754 116104
rect 230810 116048 230815 116104
rect 228988 116046 230815 116048
rect 213913 116043 213979 116046
rect 230749 116043 230815 116046
rect 262213 116106 262279 116109
rect 282361 116106 282427 116109
rect 262213 116104 268210 116106
rect 262213 116048 262218 116104
rect 262274 116048 268210 116104
rect 262213 116046 268210 116048
rect 279956 116104 282427 116106
rect 279956 116048 282366 116104
rect 282422 116048 282427 116104
rect 279956 116046 282427 116048
rect 262213 116043 262279 116046
rect 268150 115940 268210 116046
rect 282361 116043 282427 116046
rect 250437 115834 250503 115837
rect 238710 115832 250503 115834
rect 238710 115776 250442 115832
rect 250498 115776 250503 115832
rect 238710 115774 250503 115776
rect 238710 115562 238770 115774
rect 250437 115771 250503 115774
rect 228988 115502 238770 115562
rect 264973 115562 265039 115565
rect 264973 115560 268180 115562
rect 264973 115504 264978 115560
rect 265034 115504 268180 115560
rect 264973 115502 268180 115504
rect 264973 115499 265039 115502
rect 214833 115426 214899 115429
rect 282821 115426 282887 115429
rect 214833 115424 217028 115426
rect 214833 115368 214838 115424
rect 214894 115368 217028 115424
rect 214833 115366 217028 115368
rect 279956 115424 282887 115426
rect 279956 115368 282826 115424
rect 282882 115368 282887 115424
rect 279956 115366 282887 115368
rect 214833 115363 214899 115366
rect 282821 115363 282887 115366
rect 231485 115154 231551 115157
rect 228988 115152 231551 115154
rect 228988 115096 231490 115152
rect 231546 115096 231551 115152
rect 228988 115094 231551 115096
rect 231485 115091 231551 115094
rect 213913 114882 213979 114885
rect 254577 114882 254643 114885
rect 268150 114882 268210 115124
rect 213913 114880 217028 114882
rect 213913 114824 213918 114880
rect 213974 114824 217028 114880
rect 213913 114822 217028 114824
rect 254577 114880 268210 114882
rect 254577 114824 254582 114880
rect 254638 114824 268210 114880
rect 254577 114822 268210 114824
rect 213913 114819 213979 114822
rect 254577 114819 254643 114822
rect 230933 114610 230999 114613
rect 228988 114608 230999 114610
rect 228988 114552 230938 114608
rect 230994 114552 230999 114608
rect 228988 114550 230999 114552
rect 230933 114547 230999 114550
rect 262070 114548 262076 114612
rect 262140 114610 262146 114612
rect 282269 114610 282335 114613
rect 262140 114550 268180 114610
rect 279956 114608 282335 114610
rect 279956 114552 282274 114608
rect 282330 114552 282335 114608
rect 279956 114550 282335 114552
rect 262140 114548 262146 114550
rect 282269 114547 282335 114550
rect 264421 114474 264487 114477
rect 238710 114472 264487 114474
rect 238710 114416 264426 114472
rect 264482 114416 264487 114472
rect 238710 114414 264487 114416
rect 214005 114202 214071 114205
rect 238710 114202 238770 114414
rect 264421 114411 264487 114414
rect 214005 114200 217028 114202
rect 214005 114144 214010 114200
rect 214066 114144 217028 114200
rect 214005 114142 217028 114144
rect 228988 114142 238770 114202
rect 265065 114202 265131 114205
rect 265065 114200 268180 114202
rect 265065 114144 265070 114200
rect 265126 114144 268180 114200
rect 265065 114142 268180 114144
rect 214005 114139 214071 114142
rect 265065 114139 265131 114142
rect 264973 113794 265039 113797
rect 282821 113794 282887 113797
rect 264973 113792 268180 113794
rect 264973 113736 264978 113792
rect 265034 113736 268180 113792
rect 264973 113734 268180 113736
rect 279956 113792 282887 113794
rect 279956 113736 282826 113792
rect 282882 113736 282887 113792
rect 279956 113734 282887 113736
rect 264973 113731 265039 113734
rect 282821 113731 282887 113734
rect 230565 113658 230631 113661
rect 228988 113656 230631 113658
rect 228988 113600 230570 113656
rect 230626 113600 230631 113656
rect 228988 113598 230631 113600
rect 230565 113595 230631 113598
rect 213913 113522 213979 113525
rect 213913 113520 217028 113522
rect 213913 113464 213918 113520
rect 213974 113464 217028 113520
rect 213913 113462 217028 113464
rect 213913 113459 213979 113462
rect 258901 113386 258967 113389
rect 258901 113384 268180 113386
rect 258901 113328 258906 113384
rect 258962 113328 268180 113384
rect 258901 113326 268180 113328
rect 258901 113323 258967 113326
rect 231669 113250 231735 113253
rect 228988 113248 231735 113250
rect 228988 113192 231674 113248
rect 231730 113192 231735 113248
rect 228988 113190 231735 113192
rect 231669 113187 231735 113190
rect 282821 113114 282887 113117
rect 279956 113112 282887 113114
rect 279956 113056 282826 113112
rect 282882 113056 282887 113112
rect 279956 113054 282887 113056
rect 282821 113051 282887 113054
rect 214741 112842 214807 112845
rect 214741 112840 217028 112842
rect 214741 112784 214746 112840
rect 214802 112784 217028 112840
rect 214741 112782 217028 112784
rect 214741 112779 214807 112782
rect 231761 112706 231827 112709
rect 268150 112706 268210 112948
rect 582925 112842 582991 112845
rect 583520 112842 584960 112932
rect 582925 112840 584960 112842
rect 582925 112784 582930 112840
rect 582986 112784 584960 112840
rect 582925 112782 584960 112784
rect 582925 112779 582991 112782
rect 228988 112704 231827 112706
rect 228988 112648 231766 112704
rect 231822 112648 231827 112704
rect 228988 112646 231827 112648
rect 231761 112643 231827 112646
rect 258030 112646 268210 112706
rect 583520 112692 584960 112782
rect 231301 112298 231367 112301
rect 228988 112296 231367 112298
rect 228988 112240 231306 112296
rect 231362 112240 231367 112296
rect 228988 112238 231367 112240
rect 231301 112235 231367 112238
rect 213913 112162 213979 112165
rect 213913 112160 217028 112162
rect 213913 112104 213918 112160
rect 213974 112104 217028 112160
rect 213913 112102 217028 112104
rect 213913 112099 213979 112102
rect 230238 112100 230244 112164
rect 230308 112162 230314 112164
rect 258030 112162 258090 112646
rect 264973 112570 265039 112573
rect 264973 112568 268180 112570
rect 264973 112512 264978 112568
rect 265034 112512 268180 112568
rect 264973 112510 268180 112512
rect 264973 112507 265039 112510
rect 281993 112298 282059 112301
rect 279956 112296 282059 112298
rect 279956 112240 281998 112296
rect 282054 112240 282059 112296
rect 279956 112238 282059 112240
rect 281993 112235 282059 112238
rect 230308 112102 258090 112162
rect 230308 112100 230314 112102
rect 254761 112026 254827 112029
rect 254761 112024 268180 112026
rect 254761 111968 254766 112024
rect 254822 111968 268180 112024
rect 254761 111966 268180 111968
rect 254761 111963 254827 111966
rect 164724 111754 165354 111760
rect 168281 111754 168347 111757
rect 231669 111754 231735 111757
rect 164724 111752 168347 111754
rect 164724 111700 168286 111752
rect 165294 111696 168286 111700
rect 168342 111696 168347 111752
rect 165294 111694 168347 111696
rect 228988 111752 231735 111754
rect 228988 111696 231674 111752
rect 231730 111696 231735 111752
rect 228988 111694 231735 111696
rect 168281 111691 168347 111694
rect 231669 111691 231735 111694
rect 265065 111618 265131 111621
rect 284334 111618 284340 111620
rect 265065 111616 268180 111618
rect 265065 111560 265070 111616
rect 265126 111560 268180 111616
rect 265065 111558 268180 111560
rect 279956 111558 284340 111618
rect 265065 111555 265131 111558
rect 284334 111556 284340 111558
rect 284404 111556 284410 111620
rect 214005 111482 214071 111485
rect 214005 111480 217028 111482
rect 214005 111424 214010 111480
rect 214066 111424 217028 111480
rect 214005 111422 217028 111424
rect 214005 111419 214071 111422
rect 231393 111346 231459 111349
rect 228988 111344 231459 111346
rect 228988 111288 231398 111344
rect 231454 111288 231459 111344
rect 228988 111286 231459 111288
rect 231393 111283 231459 111286
rect 264973 111210 265039 111213
rect 264973 111208 268180 111210
rect 264973 111152 264978 111208
rect 265034 111152 268180 111208
rect 264973 111150 268180 111152
rect 264973 111147 265039 111150
rect 231301 111074 231367 111077
rect 250478 111074 250484 111076
rect 231301 111072 250484 111074
rect 231301 111016 231306 111072
rect 231362 111016 250484 111072
rect 231301 111014 250484 111016
rect 231301 111011 231367 111014
rect 250478 111012 250484 111014
rect 250548 111012 250554 111076
rect 213913 110802 213979 110805
rect 231761 110802 231827 110805
rect 213913 110800 217028 110802
rect -960 110666 480 110756
rect 213913 110744 213918 110800
rect 213974 110744 217028 110800
rect 213913 110742 217028 110744
rect 228988 110800 231827 110802
rect 228988 110744 231766 110800
rect 231822 110744 231827 110800
rect 228988 110742 231827 110744
rect 213913 110739 213979 110742
rect 231761 110739 231827 110742
rect 247769 110802 247835 110805
rect 282821 110802 282887 110805
rect 247769 110800 268180 110802
rect 247769 110744 247774 110800
rect 247830 110744 268180 110800
rect 247769 110742 268180 110744
rect 279956 110800 282887 110802
rect 279956 110744 282826 110800
rect 282882 110744 282887 110800
rect 279956 110742 282887 110744
rect 247769 110739 247835 110742
rect 282821 110739 282887 110742
rect 3417 110666 3483 110669
rect -960 110664 3483 110666
rect -960 110608 3422 110664
rect 3478 110608 3483 110664
rect -960 110606 3483 110608
rect -960 110516 480 110606
rect 3417 110603 3483 110606
rect 258809 110394 258875 110397
rect 228988 110392 258875 110394
rect 228988 110336 258814 110392
rect 258870 110336 258875 110392
rect 228988 110334 258875 110336
rect 258809 110331 258875 110334
rect 264421 110394 264487 110397
rect 264421 110392 268180 110394
rect 264421 110336 264426 110392
rect 264482 110336 268180 110392
rect 264421 110334 268180 110336
rect 264421 110331 264487 110334
rect 213913 110258 213979 110261
rect 213913 110256 217028 110258
rect 213913 110200 213918 110256
rect 213974 110200 217028 110256
rect 213913 110198 217028 110200
rect 213913 110195 213979 110198
rect 164724 110122 165354 110128
rect 167821 110122 167887 110125
rect 164724 110120 167887 110122
rect 164724 110068 167826 110120
rect 165294 110064 167826 110068
rect 167882 110064 167887 110120
rect 165294 110062 167887 110064
rect 167821 110059 167887 110062
rect 264973 109986 265039 109989
rect 282269 109986 282335 109989
rect 264973 109984 268180 109986
rect 264973 109928 264978 109984
rect 265034 109928 268180 109984
rect 264973 109926 268180 109928
rect 279956 109984 282335 109986
rect 279956 109928 282274 109984
rect 282330 109928 282335 109984
rect 279956 109926 282335 109928
rect 264973 109923 265039 109926
rect 282269 109923 282335 109926
rect 231209 109850 231275 109853
rect 228988 109848 231275 109850
rect 228988 109792 231214 109848
rect 231270 109792 231275 109848
rect 228988 109790 231275 109792
rect 231209 109787 231275 109790
rect 182909 109170 182975 109173
rect 216998 109170 217058 109548
rect 258030 109518 268180 109578
rect 231761 109442 231827 109445
rect 228988 109440 231827 109442
rect 228988 109384 231766 109440
rect 231822 109384 231827 109440
rect 228988 109382 231827 109384
rect 231761 109379 231827 109382
rect 242249 109442 242315 109445
rect 258030 109442 258090 109518
rect 242249 109440 258090 109442
rect 242249 109384 242254 109440
rect 242310 109384 258090 109440
rect 242249 109382 258090 109384
rect 242249 109379 242315 109382
rect 282821 109306 282887 109309
rect 279956 109304 282887 109306
rect 279956 109248 282826 109304
rect 282882 109248 282887 109304
rect 279956 109246 282887 109248
rect 282821 109243 282887 109246
rect 182909 109168 217058 109170
rect 182909 109112 182914 109168
rect 182970 109112 217058 109168
rect 182909 109110 217058 109112
rect 182909 109107 182975 109110
rect 249149 109034 249215 109037
rect 238710 109032 249215 109034
rect 238710 108976 249154 109032
rect 249210 108976 249215 109032
rect 238710 108974 249215 108976
rect 214005 108898 214071 108901
rect 238710 108898 238770 108974
rect 249149 108971 249215 108974
rect 265065 109034 265131 109037
rect 265065 109032 268180 109034
rect 265065 108976 265070 109032
rect 265126 108976 268180 109032
rect 265065 108974 268180 108976
rect 265065 108971 265131 108974
rect 214005 108896 217028 108898
rect 214005 108840 214010 108896
rect 214066 108840 217028 108896
rect 214005 108838 217028 108840
rect 228988 108838 238770 108898
rect 214005 108835 214071 108838
rect 164724 108762 165354 108768
rect 167729 108762 167795 108765
rect 164724 108760 167795 108762
rect 164724 108708 167734 108760
rect 165294 108704 167734 108708
rect 167790 108704 167795 108760
rect 165294 108702 167795 108704
rect 167729 108699 167795 108702
rect 231761 108490 231827 108493
rect 228988 108488 231827 108490
rect 228988 108432 231766 108488
rect 231822 108432 231827 108488
rect 228988 108430 231827 108432
rect 231761 108427 231827 108430
rect 180149 108354 180215 108357
rect 214557 108354 214623 108357
rect 180149 108352 214623 108354
rect 180149 108296 180154 108352
rect 180210 108296 214562 108352
rect 214618 108296 214623 108352
rect 180149 108294 214623 108296
rect 180149 108291 180215 108294
rect 214557 108291 214623 108294
rect 262765 108354 262831 108357
rect 268150 108354 268210 108596
rect 281717 108490 281783 108493
rect 279956 108488 281783 108490
rect 279956 108432 281722 108488
rect 281778 108432 281783 108488
rect 279956 108430 281783 108432
rect 281717 108427 281783 108430
rect 262765 108352 268210 108354
rect 262765 108296 262770 108352
rect 262826 108296 268210 108352
rect 262765 108294 268210 108296
rect 262765 108291 262831 108294
rect 213913 108218 213979 108221
rect 213913 108216 217028 108218
rect 213913 108160 213918 108216
rect 213974 108160 217028 108216
rect 213913 108158 217028 108160
rect 258030 108158 268180 108218
rect 213913 108155 213979 108158
rect 250437 108082 250503 108085
rect 258030 108082 258090 108158
rect 250437 108080 258090 108082
rect 250437 108024 250442 108080
rect 250498 108024 258090 108080
rect 250437 108022 258090 108024
rect 250437 108019 250503 108022
rect 231393 107946 231459 107949
rect 228988 107944 231459 107946
rect 228988 107888 231398 107944
rect 231454 107888 231459 107944
rect 228988 107886 231459 107888
rect 231393 107883 231459 107886
rect 243721 107946 243787 107949
rect 262765 107946 262831 107949
rect 243721 107944 262831 107946
rect 243721 107888 243726 107944
rect 243782 107888 262770 107944
rect 262826 107888 262831 107944
rect 243721 107886 262831 107888
rect 243721 107883 243787 107886
rect 262765 107883 262831 107886
rect 264973 107810 265039 107813
rect 282177 107810 282243 107813
rect 264973 107808 268180 107810
rect 264973 107752 264978 107808
rect 265034 107752 268180 107808
rect 264973 107750 268180 107752
rect 279956 107808 282243 107810
rect 279956 107752 282182 107808
rect 282238 107752 282243 107808
rect 279956 107750 282243 107752
rect 264973 107747 265039 107750
rect 282177 107747 282243 107750
rect 214005 107538 214071 107541
rect 240869 107538 240935 107541
rect 214005 107536 217028 107538
rect 214005 107480 214010 107536
rect 214066 107480 217028 107536
rect 214005 107478 217028 107480
rect 228988 107536 240935 107538
rect 228988 107480 240874 107536
rect 240930 107480 240935 107536
rect 228988 107478 240935 107480
rect 214005 107475 214071 107478
rect 240869 107475 240935 107478
rect 265065 107402 265131 107405
rect 265065 107400 268180 107402
rect 265065 107344 265070 107400
rect 265126 107344 268180 107400
rect 265065 107342 268180 107344
rect 265065 107339 265131 107342
rect 231209 107130 231275 107133
rect 228988 107128 231275 107130
rect 228988 107072 231214 107128
rect 231270 107072 231275 107128
rect 228988 107070 231275 107072
rect 231209 107067 231275 107070
rect 264973 106994 265039 106997
rect 285622 106994 285628 106996
rect 264973 106992 268180 106994
rect 264973 106936 264978 106992
rect 265034 106936 268180 106992
rect 264973 106934 268180 106936
rect 279956 106934 285628 106994
rect 264973 106931 265039 106934
rect 285622 106932 285628 106934
rect 285692 106932 285698 106996
rect 213913 106858 213979 106861
rect 213913 106856 217028 106858
rect 213913 106800 213918 106856
rect 213974 106800 217028 106856
rect 213913 106798 217028 106800
rect 213913 106795 213979 106798
rect 231761 106586 231827 106589
rect 228988 106584 231827 106586
rect 228988 106528 231766 106584
rect 231822 106528 231827 106584
rect 228988 106526 231827 106528
rect 231761 106523 231827 106526
rect 258030 106390 268180 106450
rect 241053 106314 241119 106317
rect 258030 106314 258090 106390
rect 241053 106312 258090 106314
rect 241053 106256 241058 106312
rect 241114 106256 258090 106312
rect 241053 106254 258090 106256
rect 241053 106251 241119 106254
rect 214005 106178 214071 106181
rect 242014 106178 242020 106180
rect 214005 106176 217028 106178
rect 214005 106120 214010 106176
rect 214066 106120 217028 106176
rect 214005 106118 217028 106120
rect 228988 106118 242020 106178
rect 214005 106115 214071 106118
rect 242014 106116 242020 106118
rect 242084 106116 242090 106180
rect 264973 106042 265039 106045
rect 264973 106040 268180 106042
rect 264973 105984 264978 106040
rect 265034 105984 268180 106040
rect 264973 105982 268180 105984
rect 264973 105979 265039 105982
rect 214373 105634 214439 105637
rect 229921 105634 229987 105637
rect 214373 105632 217028 105634
rect 214373 105576 214378 105632
rect 214434 105576 217028 105632
rect 214373 105574 217028 105576
rect 228988 105632 229987 105634
rect 228988 105576 229926 105632
rect 229982 105576 229987 105632
rect 228988 105574 229987 105576
rect 214373 105571 214439 105574
rect 229921 105571 229987 105574
rect 265065 105634 265131 105637
rect 279926 105634 279986 106148
rect 265065 105632 268180 105634
rect 265065 105576 265070 105632
rect 265126 105576 268180 105632
rect 265065 105574 268180 105576
rect 279926 105574 287070 105634
rect 265065 105571 265131 105574
rect 282821 105498 282887 105501
rect 279956 105496 282887 105498
rect 279956 105440 282826 105496
rect 282882 105440 282887 105496
rect 279956 105438 282887 105440
rect 282821 105435 282887 105438
rect 231761 105226 231827 105229
rect 228988 105224 231827 105226
rect 228988 105168 231766 105224
rect 231822 105168 231827 105224
rect 228988 105166 231827 105168
rect 231761 105163 231827 105166
rect 267181 105226 267247 105229
rect 267181 105224 268180 105226
rect 267181 105168 267186 105224
rect 267242 105168 268180 105224
rect 267181 105166 268180 105168
rect 267181 105163 267247 105166
rect 213913 104954 213979 104957
rect 287010 104954 287070 105574
rect 288566 104954 288572 104956
rect 213913 104952 217028 104954
rect 213913 104896 213918 104952
rect 213974 104896 217028 104952
rect 213913 104894 217028 104896
rect 287010 104894 288572 104954
rect 213913 104891 213979 104894
rect 288566 104892 288572 104894
rect 288636 104892 288642 104956
rect 264973 104818 265039 104821
rect 264973 104816 268180 104818
rect 264973 104760 264978 104816
rect 265034 104760 268180 104816
rect 264973 104758 268180 104760
rect 264973 104755 265039 104758
rect 231117 104682 231183 104685
rect 282821 104682 282887 104685
rect 228988 104680 231183 104682
rect 228988 104624 231122 104680
rect 231178 104624 231183 104680
rect 228988 104622 231183 104624
rect 279956 104680 282887 104682
rect 279956 104624 282826 104680
rect 282882 104624 282887 104680
rect 279956 104622 282887 104624
rect 231117 104619 231183 104622
rect 282821 104619 282887 104622
rect 231301 104274 231367 104277
rect 228988 104272 231367 104274
rect 166390 103804 166396 103868
rect 166460 103866 166466 103868
rect 216998 103866 217058 104244
rect 228988 104216 231306 104272
rect 231362 104216 231367 104272
rect 228988 104214 231367 104216
rect 231301 104211 231367 104214
rect 239673 104002 239739 104005
rect 268150 104002 268210 104380
rect 281993 104002 282059 104005
rect 239673 104000 268210 104002
rect 239673 103944 239678 104000
rect 239734 103944 268210 104000
rect 239673 103942 268210 103944
rect 279956 104000 282059 104002
rect 279956 103944 281998 104000
rect 282054 103944 282059 104000
rect 279956 103942 282059 103944
rect 239673 103939 239739 103942
rect 281993 103939 282059 103942
rect 166460 103806 217058 103866
rect 258030 103806 268180 103866
rect 166460 103804 166466 103806
rect 231301 103730 231367 103733
rect 228988 103728 231367 103730
rect 228988 103672 231306 103728
rect 231362 103672 231367 103728
rect 228988 103670 231367 103672
rect 231301 103667 231367 103670
rect 245101 103730 245167 103733
rect 258030 103730 258090 103806
rect 245101 103728 258090 103730
rect 245101 103672 245106 103728
rect 245162 103672 258090 103728
rect 245101 103670 258090 103672
rect 245101 103667 245167 103670
rect 213913 103594 213979 103597
rect 213913 103592 217028 103594
rect 213913 103536 213918 103592
rect 213974 103536 217028 103592
rect 213913 103534 217028 103536
rect 213913 103531 213979 103534
rect 264973 103458 265039 103461
rect 264973 103456 268180 103458
rect 264973 103400 264978 103456
rect 265034 103400 268180 103456
rect 264973 103398 268180 103400
rect 264973 103395 265039 103398
rect 231485 103322 231551 103325
rect 228988 103320 231551 103322
rect 228988 103264 231490 103320
rect 231546 103264 231551 103320
rect 228988 103262 231551 103264
rect 231485 103259 231551 103262
rect 282821 103186 282887 103189
rect 279956 103184 282887 103186
rect 279956 103128 282826 103184
rect 282882 103128 282887 103184
rect 279956 103126 282887 103128
rect 282821 103123 282887 103126
rect 264789 103050 264855 103053
rect 264789 103048 268180 103050
rect 264789 102992 264794 103048
rect 264850 102992 268180 103048
rect 264789 102990 268180 102992
rect 264789 102987 264855 102990
rect 214005 102914 214071 102917
rect 231301 102914 231367 102917
rect 250805 102914 250871 102917
rect 214005 102912 217028 102914
rect 214005 102856 214010 102912
rect 214066 102856 217028 102912
rect 214005 102854 217028 102856
rect 231301 102912 250871 102914
rect 231301 102856 231306 102912
rect 231362 102856 250810 102912
rect 250866 102856 250871 102912
rect 231301 102854 250871 102856
rect 214005 102851 214071 102854
rect 231301 102851 231367 102854
rect 250805 102851 250871 102854
rect 230565 102778 230631 102781
rect 228988 102776 230631 102778
rect 228988 102720 230570 102776
rect 230626 102720 230631 102776
rect 228988 102718 230631 102720
rect 230565 102715 230631 102718
rect 232865 102778 232931 102781
rect 260046 102778 260052 102780
rect 232865 102776 260052 102778
rect 232865 102720 232870 102776
rect 232926 102720 260052 102776
rect 232865 102718 260052 102720
rect 232865 102715 232931 102718
rect 260046 102716 260052 102718
rect 260116 102716 260122 102780
rect 263041 102642 263107 102645
rect 263041 102640 268180 102642
rect 263041 102584 263046 102640
rect 263102 102584 268180 102640
rect 263041 102582 268180 102584
rect 263041 102579 263107 102582
rect 65977 102370 66043 102373
rect 68142 102370 68816 102376
rect 231577 102370 231643 102373
rect 282729 102370 282795 102373
rect 65977 102368 68816 102370
rect 65977 102312 65982 102368
rect 66038 102316 68816 102368
rect 228988 102368 231643 102370
rect 66038 102312 68202 102316
rect 65977 102310 68202 102312
rect 228988 102312 231582 102368
rect 231638 102312 231643 102368
rect 228988 102310 231643 102312
rect 279956 102368 282795 102370
rect 279956 102312 282734 102368
rect 282790 102312 282795 102368
rect 279956 102310 282795 102312
rect 65977 102307 66043 102310
rect 231577 102307 231643 102310
rect 282729 102307 282795 102310
rect 213913 102234 213979 102237
rect 243629 102234 243695 102237
rect 213913 102232 217028 102234
rect 213913 102176 213918 102232
rect 213974 102176 217028 102232
rect 213913 102174 217028 102176
rect 243629 102232 268180 102234
rect 243629 102176 243634 102232
rect 243690 102176 268180 102232
rect 243629 102174 268180 102176
rect 213913 102171 213979 102174
rect 243629 102171 243695 102174
rect 231209 101826 231275 101829
rect 228988 101824 231275 101826
rect 228988 101768 231214 101824
rect 231270 101768 231275 101824
rect 228988 101766 231275 101768
rect 231209 101763 231275 101766
rect 264973 101826 265039 101829
rect 264973 101824 268180 101826
rect 264973 101768 264978 101824
rect 265034 101768 268180 101824
rect 264973 101766 268180 101768
rect 264973 101763 265039 101766
rect 282821 101690 282887 101693
rect 279956 101688 282887 101690
rect 279956 101632 282826 101688
rect 282882 101632 282887 101688
rect 279956 101630 282887 101632
rect 282821 101627 282887 101630
rect 213913 101554 213979 101557
rect 213913 101552 217028 101554
rect 213913 101496 213918 101552
rect 213974 101496 217028 101552
rect 213913 101494 217028 101496
rect 213913 101491 213979 101494
rect 168966 101356 168972 101420
rect 169036 101418 169042 101420
rect 214373 101418 214439 101421
rect 231393 101418 231459 101421
rect 169036 101416 214439 101418
rect 169036 101360 214378 101416
rect 214434 101360 214439 101416
rect 169036 101358 214439 101360
rect 228988 101416 231459 101418
rect 228988 101360 231398 101416
rect 231454 101360 231459 101416
rect 228988 101358 231459 101360
rect 169036 101356 169042 101358
rect 214373 101355 214439 101358
rect 231393 101355 231459 101358
rect 231577 101418 231643 101421
rect 260281 101418 260347 101421
rect 231577 101416 260347 101418
rect 231577 101360 231582 101416
rect 231638 101360 260286 101416
rect 260342 101360 260347 101416
rect 231577 101358 260347 101360
rect 231577 101355 231643 101358
rect 260281 101355 260347 101358
rect 265065 101282 265131 101285
rect 265065 101280 268180 101282
rect 265065 101224 265070 101280
rect 265126 101224 268180 101280
rect 265065 101222 268180 101224
rect 265065 101219 265131 101222
rect 214833 101010 214899 101013
rect 214833 101008 217028 101010
rect 214833 100952 214838 101008
rect 214894 100952 217028 101008
rect 214833 100950 217028 100952
rect 214833 100947 214899 100950
rect 231669 100874 231735 100877
rect 228988 100872 231735 100874
rect 228988 100816 231674 100872
rect 231730 100816 231735 100872
rect 228988 100814 231735 100816
rect 231669 100811 231735 100814
rect 261753 100874 261819 100877
rect 281533 100874 281599 100877
rect 261753 100872 268180 100874
rect 261753 100816 261758 100872
rect 261814 100816 268180 100872
rect 261753 100814 268180 100816
rect 279956 100872 281599 100874
rect 279956 100816 281538 100872
rect 281594 100816 281599 100872
rect 279956 100814 281599 100816
rect 261753 100811 261819 100814
rect 281533 100811 281599 100814
rect 67265 100738 67331 100741
rect 68142 100738 68816 100744
rect 67265 100736 68816 100738
rect 67265 100680 67270 100736
rect 67326 100684 68816 100736
rect 67326 100680 68202 100684
rect 67265 100678 68202 100680
rect 67265 100675 67331 100678
rect 231761 100466 231827 100469
rect 228988 100464 231827 100466
rect 228988 100408 231766 100464
rect 231822 100408 231827 100464
rect 228988 100406 231827 100408
rect 231761 100403 231827 100406
rect 262990 100404 262996 100468
rect 263060 100466 263066 100468
rect 263060 100406 268180 100466
rect 263060 100404 263066 100406
rect 214005 100330 214071 100333
rect 214005 100328 217028 100330
rect 214005 100272 214010 100328
rect 214066 100272 217028 100328
rect 214005 100270 217028 100272
rect 214005 100267 214071 100270
rect 281717 100194 281783 100197
rect 279956 100192 281783 100194
rect 279956 100136 281722 100192
rect 281778 100136 281783 100192
rect 279956 100134 281783 100136
rect 281717 100131 281783 100134
rect 231669 99922 231735 99925
rect 228988 99920 231735 99922
rect 228988 99864 231674 99920
rect 231730 99864 231735 99920
rect 228988 99862 231735 99864
rect 231669 99859 231735 99862
rect 260046 99724 260052 99788
rect 260116 99786 260122 99788
rect 268150 99786 268210 100028
rect 260116 99726 268210 99786
rect 260116 99724 260122 99726
rect 213913 99650 213979 99653
rect 264973 99650 265039 99653
rect 213913 99648 217028 99650
rect 213913 99592 213918 99648
rect 213974 99592 217028 99648
rect 213913 99590 217028 99592
rect 264973 99648 268180 99650
rect 264973 99592 264978 99648
rect 265034 99592 268180 99648
rect 264973 99590 268180 99592
rect 213913 99587 213979 99590
rect 264973 99587 265039 99590
rect 231577 99514 231643 99517
rect 228988 99512 231643 99514
rect 228988 99456 231582 99512
rect 231638 99456 231643 99512
rect 228988 99454 231643 99456
rect 231577 99451 231643 99454
rect 583017 99514 583083 99517
rect 583520 99514 584960 99604
rect 583017 99512 584960 99514
rect 583017 99456 583022 99512
rect 583078 99456 584960 99512
rect 583017 99454 584960 99456
rect 583017 99451 583083 99454
rect 583520 99364 584960 99454
rect 263174 99180 263180 99244
rect 263244 99242 263250 99244
rect 263244 99182 268180 99242
rect 263244 99180 263250 99182
rect 214005 98970 214071 98973
rect 231209 98970 231275 98973
rect 214005 98968 217028 98970
rect 214005 98912 214010 98968
rect 214066 98912 217028 98968
rect 214005 98910 217028 98912
rect 228988 98968 231275 98970
rect 228988 98912 231214 98968
rect 231270 98912 231275 98968
rect 228988 98910 231275 98912
rect 214005 98907 214071 98910
rect 231209 98907 231275 98910
rect 279374 98837 279434 99348
rect 231117 98834 231183 98837
rect 238150 98834 238156 98836
rect 231117 98832 238156 98834
rect 231117 98776 231122 98832
rect 231178 98776 238156 98832
rect 231117 98774 238156 98776
rect 231117 98771 231183 98774
rect 238150 98772 238156 98774
rect 238220 98772 238226 98836
rect 245009 98834 245075 98837
rect 262990 98834 262996 98836
rect 245009 98832 262996 98834
rect 245009 98776 245014 98832
rect 245070 98776 262996 98832
rect 245009 98774 262996 98776
rect 245009 98771 245075 98774
rect 262990 98772 262996 98774
rect 263060 98772 263066 98836
rect 279374 98832 279483 98837
rect 279374 98776 279422 98832
rect 279478 98776 279483 98832
rect 279374 98774 279483 98776
rect 279417 98771 279483 98774
rect 232681 98698 232747 98701
rect 237005 98698 237071 98701
rect 232681 98696 237071 98698
rect 232681 98640 232686 98696
rect 232742 98640 237010 98696
rect 237066 98640 237071 98696
rect 232681 98638 237071 98640
rect 232681 98635 232747 98638
rect 237005 98635 237071 98638
rect 239489 98698 239555 98701
rect 264789 98698 264855 98701
rect 239489 98696 264855 98698
rect 239489 98640 239494 98696
rect 239550 98640 264794 98696
rect 264850 98640 264855 98696
rect 239489 98638 264855 98640
rect 239489 98635 239555 98638
rect 264789 98635 264855 98638
rect 264973 98698 265039 98701
rect 264973 98696 268180 98698
rect 264973 98640 264978 98696
rect 265034 98640 268180 98696
rect 264973 98638 268180 98640
rect 264973 98635 265039 98638
rect 231393 98562 231459 98565
rect 228988 98560 231459 98562
rect 228988 98504 231398 98560
rect 231454 98504 231459 98560
rect 228988 98502 231459 98504
rect 231393 98499 231459 98502
rect 213913 98290 213979 98293
rect 267733 98290 267799 98293
rect 213913 98288 217028 98290
rect 213913 98232 213918 98288
rect 213974 98232 217028 98288
rect 213913 98230 217028 98232
rect 267733 98288 268180 98290
rect 267733 98232 267738 98288
rect 267794 98232 268180 98288
rect 267733 98230 268180 98232
rect 213913 98227 213979 98230
rect 267733 98227 267799 98230
rect 279374 98157 279434 98532
rect 279325 98152 279434 98157
rect 279325 98096 279330 98152
rect 279386 98096 279434 98152
rect 279325 98094 279434 98096
rect 279325 98091 279391 98094
rect 232446 98018 232452 98020
rect 228988 97958 232452 98018
rect 232446 97956 232452 97958
rect 232516 97956 232522 98020
rect 229093 97882 229159 97885
rect 263225 97882 263291 97885
rect 282269 97882 282335 97885
rect 229093 97880 263291 97882
rect 229093 97824 229098 97880
rect 229154 97824 263230 97880
rect 263286 97824 263291 97880
rect 279956 97880 282335 97882
rect 229093 97822 263291 97824
rect 229093 97819 229159 97822
rect 263225 97819 263291 97822
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 213453 97610 213519 97613
rect 231209 97610 231275 97613
rect 268518 97612 268578 97852
rect 279956 97824 282274 97880
rect 282330 97824 282335 97880
rect 279956 97822 282335 97824
rect 282269 97819 282335 97822
rect 213453 97608 217028 97610
rect 213453 97552 213458 97608
rect 213514 97552 217028 97608
rect 213453 97550 217028 97552
rect 228988 97608 231275 97610
rect 228988 97552 231214 97608
rect 231270 97552 231275 97608
rect 228988 97550 231275 97552
rect 213453 97547 213519 97550
rect 231209 97547 231275 97550
rect 268510 97548 268516 97612
rect 268580 97548 268586 97612
rect 264973 97474 265039 97477
rect 264973 97472 268180 97474
rect 264973 97416 264978 97472
rect 265034 97416 268180 97472
rect 264973 97414 268180 97416
rect 264973 97411 265039 97414
rect 265893 97066 265959 97069
rect 281717 97066 281783 97069
rect 228988 97006 231410 97066
rect 214833 96930 214899 96933
rect 214833 96928 217028 96930
rect 214833 96872 214838 96928
rect 214894 96872 217028 96928
rect 214833 96870 217028 96872
rect 214833 96867 214899 96870
rect 168414 96596 168420 96660
rect 168484 96658 168490 96660
rect 169569 96658 169635 96661
rect 229134 96658 229140 96660
rect 168484 96656 169635 96658
rect 168484 96600 169574 96656
rect 169630 96600 169635 96656
rect 168484 96598 169635 96600
rect 228988 96598 229140 96658
rect 168484 96596 168490 96598
rect 169569 96595 169635 96598
rect 229134 96596 229140 96598
rect 229204 96658 229210 96660
rect 230749 96658 230815 96661
rect 229204 96656 230815 96658
rect 229204 96600 230754 96656
rect 230810 96600 230815 96656
rect 229204 96598 230815 96600
rect 229204 96596 229210 96598
rect 230749 96595 230815 96598
rect 231209 96522 231275 96525
rect 231350 96522 231410 97006
rect 265893 97064 268180 97066
rect 265893 97008 265898 97064
rect 265954 97008 268180 97064
rect 265893 97006 268180 97008
rect 279956 97064 281783 97066
rect 279956 97008 281722 97064
rect 281778 97008 281783 97064
rect 279956 97006 281783 97008
rect 265893 97003 265959 97006
rect 281717 97003 281783 97006
rect 265065 96658 265131 96661
rect 265065 96656 268180 96658
rect 265065 96600 265070 96656
rect 265126 96600 268180 96656
rect 265065 96598 268180 96600
rect 265065 96595 265131 96598
rect 244273 96522 244339 96525
rect 244774 96522 244780 96524
rect 231209 96520 244780 96522
rect 231209 96464 231214 96520
rect 231270 96464 244278 96520
rect 244334 96464 244780 96520
rect 231209 96462 244780 96464
rect 231209 96459 231275 96462
rect 244273 96459 244339 96462
rect 244774 96460 244780 96462
rect 244844 96460 244850 96524
rect 213913 96386 213979 96389
rect 262673 96386 262739 96389
rect 263174 96386 263180 96388
rect 213913 96384 217028 96386
rect 213913 96328 213918 96384
rect 213974 96328 217028 96384
rect 213913 96326 217028 96328
rect 262673 96384 263180 96386
rect 262673 96328 262678 96384
rect 262734 96328 263180 96384
rect 262673 96326 263180 96328
rect 213913 96323 213979 96326
rect 262673 96323 262739 96326
rect 263174 96324 263180 96326
rect 263244 96324 263250 96388
rect 230473 96250 230539 96253
rect 228988 96248 230539 96250
rect 228988 96192 230478 96248
rect 230534 96192 230539 96248
rect 228988 96190 230539 96192
rect 230473 96187 230539 96190
rect 223665 95980 223731 95981
rect 223614 95978 223620 95980
rect 223574 95918 223620 95978
rect 223684 95976 223731 95980
rect 223726 95920 223731 95976
rect 223614 95916 223620 95918
rect 223684 95916 223731 95920
rect 223665 95915 223731 95916
rect 229093 95298 229159 95301
rect 230238 95298 230244 95300
rect 229093 95296 230244 95298
rect 229093 95240 229098 95296
rect 229154 95240 230244 95296
rect 229093 95238 230244 95240
rect 229093 95235 229159 95238
rect 230238 95236 230244 95238
rect 230308 95236 230314 95300
rect 246481 95298 246547 95301
rect 268150 95298 268210 96220
rect 279926 95842 279986 96356
rect 280061 95842 280127 95845
rect 279926 95840 280127 95842
rect 279926 95784 280066 95840
rect 280122 95784 280127 95840
rect 279926 95782 280127 95784
rect 280061 95779 280127 95782
rect 246481 95296 268210 95298
rect 246481 95240 246486 95296
rect 246542 95240 268210 95296
rect 246481 95238 268210 95240
rect 246481 95235 246547 95238
rect 205398 95100 205404 95164
rect 205468 95162 205474 95164
rect 279325 95162 279391 95165
rect 205468 95160 279391 95162
rect 205468 95104 279330 95160
rect 279386 95104 279391 95160
rect 205468 95102 279391 95104
rect 205468 95100 205474 95102
rect 279325 95099 279391 95102
rect 212390 94964 212396 95028
rect 212460 95026 212466 95028
rect 279417 95026 279483 95029
rect 212460 95024 279483 95026
rect 212460 94968 279422 95024
rect 279478 94968 279483 95024
rect 212460 94966 279483 94968
rect 212460 94964 212466 94966
rect 279417 94963 279483 94966
rect 106472 94828 106478 94892
rect 106542 94890 106548 94892
rect 106774 94890 106780 94892
rect 106542 94830 106780 94890
rect 106542 94828 106548 94830
rect 106774 94828 106780 94830
rect 106844 94828 106850 94892
rect 151302 94828 151308 94892
rect 151372 94890 151378 94892
rect 151760 94890 151766 94892
rect 151372 94830 151766 94890
rect 151372 94828 151378 94830
rect 151760 94828 151766 94830
rect 151830 94828 151836 94892
rect 162117 94890 162183 94893
rect 169293 94890 169359 94893
rect 162117 94888 169359 94890
rect 162117 94832 162122 94888
rect 162178 94832 169298 94888
rect 169354 94832 169359 94888
rect 162117 94830 169359 94832
rect 162117 94827 162183 94830
rect 169293 94827 169359 94830
rect 268510 94828 268516 94892
rect 268580 94890 268586 94892
rect 269113 94890 269179 94893
rect 268580 94888 269179 94890
rect 268580 94832 269118 94888
rect 269174 94832 269179 94888
rect 268580 94830 269179 94832
rect 268580 94828 268586 94830
rect 269113 94827 269179 94830
rect 110137 94756 110203 94757
rect 125409 94756 125475 94757
rect 106222 94692 106228 94756
rect 106292 94754 106298 94756
rect 106608 94754 106614 94756
rect 106292 94694 106614 94754
rect 106292 94692 106298 94694
rect 106608 94692 106614 94694
rect 106678 94692 106684 94756
rect 110137 94754 110150 94756
rect 110058 94752 110150 94754
rect 110058 94696 110142 94752
rect 110058 94694 110150 94696
rect 110137 94692 110150 94694
rect 110214 94692 110220 94756
rect 125376 94692 125382 94756
rect 125446 94754 125475 94756
rect 125446 94752 125538 94754
rect 125470 94696 125538 94752
rect 125446 94694 125538 94696
rect 125446 94692 125475 94694
rect 110137 94691 110203 94692
rect 125409 94691 125475 94692
rect 121453 94482 121519 94485
rect 166206 94482 166212 94484
rect 121453 94480 166212 94482
rect 121453 94424 121458 94480
rect 121514 94424 166212 94480
rect 121453 94422 166212 94424
rect 121453 94419 121519 94422
rect 166206 94420 166212 94422
rect 166276 94420 166282 94484
rect 98494 93876 98500 93940
rect 98564 93938 98570 93940
rect 209129 93938 209195 93941
rect 98564 93936 209195 93938
rect 98564 93880 209134 93936
rect 209190 93880 209195 93936
rect 98564 93878 209195 93880
rect 98564 93876 98570 93878
rect 209129 93875 209195 93878
rect 131982 93740 131988 93804
rect 132052 93802 132058 93804
rect 203517 93802 203583 93805
rect 132052 93800 203583 93802
rect 132052 93744 203522 93800
rect 203578 93744 203583 93800
rect 132052 93742 203583 93744
rect 132052 93740 132058 93742
rect 203517 93739 203583 93742
rect 111926 93604 111932 93668
rect 111996 93666 112002 93668
rect 167637 93666 167703 93669
rect 111996 93664 167703 93666
rect 111996 93608 167642 93664
rect 167698 93608 167703 93664
rect 111996 93606 167703 93608
rect 111996 93604 112002 93606
rect 167637 93603 167703 93606
rect 200614 93604 200620 93668
rect 200684 93666 200690 93668
rect 280061 93666 280127 93669
rect 200684 93664 280127 93666
rect 200684 93608 280066 93664
rect 280122 93608 280127 93664
rect 200684 93606 280127 93608
rect 200684 93604 200690 93606
rect 280061 93603 280127 93606
rect 108113 93532 108179 93533
rect 121729 93532 121795 93533
rect 108062 93530 108068 93532
rect 108022 93470 108068 93530
rect 108132 93528 108179 93532
rect 121678 93530 121684 93532
rect 108174 93472 108179 93528
rect 108062 93468 108068 93470
rect 108132 93468 108179 93472
rect 121638 93470 121684 93530
rect 121748 93528 121795 93532
rect 121790 93472 121795 93528
rect 121678 93468 121684 93470
rect 121748 93468 121795 93472
rect 123150 93468 123156 93532
rect 123220 93530 123226 93532
rect 170397 93530 170463 93533
rect 123220 93528 170463 93530
rect 123220 93472 170402 93528
rect 170458 93472 170463 93528
rect 123220 93470 170463 93472
rect 123220 93468 123226 93470
rect 108113 93467 108179 93468
rect 121729 93467 121795 93468
rect 170397 93467 170463 93470
rect 66069 93122 66135 93125
rect 122097 93122 122163 93125
rect 66069 93120 122163 93122
rect 66069 93064 66074 93120
rect 66130 93064 122102 93120
rect 122158 93064 122163 93120
rect 66069 93062 122163 93064
rect 66069 93059 66135 93062
rect 122097 93059 122163 93062
rect 169201 93122 169267 93125
rect 178953 93122 179019 93125
rect 169201 93120 179019 93122
rect 169201 93064 169206 93120
rect 169262 93064 178958 93120
rect 179014 93064 179019 93120
rect 169201 93062 179019 93064
rect 169201 93059 169267 93062
rect 178953 93059 179019 93062
rect 228357 93122 228423 93125
rect 250621 93122 250687 93125
rect 228357 93120 250687 93122
rect 228357 93064 228362 93120
rect 228418 93064 250626 93120
rect 250682 93064 250687 93120
rect 228357 93062 250687 93064
rect 228357 93059 228423 93062
rect 250621 93059 250687 93062
rect 100017 92444 100083 92445
rect 105721 92444 105787 92445
rect 99966 92442 99972 92444
rect 99926 92382 99972 92442
rect 100036 92440 100083 92444
rect 105670 92442 105676 92444
rect 100078 92384 100083 92440
rect 99966 92380 99972 92382
rect 100036 92380 100083 92384
rect 105630 92382 105676 92442
rect 105740 92440 105787 92444
rect 105782 92384 105787 92440
rect 105670 92380 105676 92382
rect 105740 92380 105787 92384
rect 111190 92380 111196 92444
rect 111260 92442 111266 92444
rect 111609 92442 111675 92445
rect 111260 92440 111675 92442
rect 111260 92384 111614 92440
rect 111670 92384 111675 92440
rect 111260 92382 111675 92384
rect 111260 92380 111266 92382
rect 100017 92379 100083 92380
rect 105721 92379 105787 92380
rect 111609 92379 111675 92382
rect 113214 92380 113220 92444
rect 113284 92442 113290 92444
rect 113449 92442 113515 92445
rect 115473 92444 115539 92445
rect 118049 92444 118115 92445
rect 136081 92444 136147 92445
rect 152089 92444 152155 92445
rect 115422 92442 115428 92444
rect 113284 92440 113515 92442
rect 113284 92384 113454 92440
rect 113510 92384 113515 92440
rect 113284 92382 113515 92384
rect 115382 92382 115428 92442
rect 115492 92440 115539 92444
rect 117998 92442 118004 92444
rect 115534 92384 115539 92440
rect 113284 92380 113290 92382
rect 113449 92379 113515 92382
rect 115422 92380 115428 92382
rect 115492 92380 115539 92384
rect 117958 92382 118004 92442
rect 118068 92440 118115 92444
rect 136030 92442 136036 92444
rect 118110 92384 118115 92440
rect 117998 92380 118004 92382
rect 118068 92380 118115 92384
rect 135990 92382 136036 92442
rect 136100 92440 136147 92444
rect 152038 92442 152044 92444
rect 136142 92384 136147 92440
rect 136030 92380 136036 92382
rect 136100 92380 136147 92384
rect 151998 92382 152044 92442
rect 152108 92440 152155 92444
rect 152150 92384 152155 92440
rect 152038 92380 152044 92382
rect 152108 92380 152155 92384
rect 115473 92379 115539 92380
rect 118049 92379 118115 92380
rect 136081 92379 136147 92380
rect 152089 92379 152155 92380
rect 125726 92244 125732 92308
rect 125796 92306 125802 92308
rect 192569 92306 192635 92309
rect 125796 92304 192635 92306
rect 125796 92248 192574 92304
rect 192630 92248 192635 92304
rect 125796 92246 192635 92248
rect 125796 92244 125802 92246
rect 192569 92243 192635 92246
rect 127566 92108 127572 92172
rect 127636 92170 127642 92172
rect 166533 92170 166599 92173
rect 127636 92168 166599 92170
rect 127636 92112 166538 92168
rect 166594 92112 166599 92168
rect 127636 92110 166599 92112
rect 127636 92108 127642 92110
rect 166533 92107 166599 92110
rect 106222 91972 106228 92036
rect 106292 92034 106298 92036
rect 124857 92034 124923 92037
rect 106292 92032 124923 92034
rect 106292 91976 124862 92032
rect 124918 91976 124923 92032
rect 106292 91974 124923 91976
rect 106292 91972 106298 91974
rect 124857 91971 124923 91974
rect 85798 91700 85804 91764
rect 85868 91762 85874 91764
rect 86493 91762 86559 91765
rect 85868 91760 86559 91762
rect 85868 91704 86498 91760
rect 86554 91704 86559 91760
rect 85868 91702 86559 91704
rect 85868 91700 85874 91702
rect 86493 91699 86559 91702
rect 104198 91700 104204 91764
rect 104268 91762 104274 91764
rect 104525 91762 104591 91765
rect 104268 91760 104591 91762
rect 104268 91704 104530 91760
rect 104586 91704 104591 91760
rect 104268 91702 104591 91704
rect 104268 91700 104274 91702
rect 104525 91699 104591 91702
rect 112294 91700 112300 91764
rect 112364 91762 112370 91764
rect 112621 91762 112687 91765
rect 112364 91760 112687 91762
rect 112364 91704 112626 91760
rect 112682 91704 112687 91760
rect 112364 91702 112687 91704
rect 112364 91700 112370 91702
rect 112621 91699 112687 91702
rect 114870 91700 114876 91764
rect 114940 91762 114946 91764
rect 115565 91762 115631 91765
rect 114940 91760 115631 91762
rect 114940 91704 115570 91760
rect 115626 91704 115631 91760
rect 114940 91702 115631 91704
rect 114940 91700 114946 91702
rect 115565 91699 115631 91702
rect 120574 91700 120580 91764
rect 120644 91762 120650 91764
rect 121177 91762 121243 91765
rect 120644 91760 121243 91762
rect 120644 91704 121182 91760
rect 121238 91704 121243 91760
rect 120644 91702 121243 91704
rect 120644 91700 120650 91702
rect 121177 91699 121243 91702
rect 195237 91762 195303 91765
rect 277393 91762 277459 91765
rect 195237 91760 277459 91762
rect 195237 91704 195242 91760
rect 195298 91704 277398 91760
rect 277454 91704 277459 91760
rect 195237 91702 277459 91704
rect 195237 91699 195303 91702
rect 277393 91699 277459 91702
rect 100886 91564 100892 91628
rect 100956 91626 100962 91628
rect 209221 91626 209287 91629
rect 100956 91624 209287 91626
rect 100956 91568 209226 91624
rect 209282 91568 209287 91624
rect 100956 91566 209287 91568
rect 100956 91564 100962 91566
rect 209221 91563 209287 91566
rect 122782 91428 122788 91492
rect 122852 91490 122858 91492
rect 124029 91490 124095 91493
rect 151537 91492 151603 91493
rect 151486 91490 151492 91492
rect 122852 91488 124095 91490
rect 122852 91432 124034 91488
rect 124090 91432 124095 91488
rect 122852 91430 124095 91432
rect 151446 91430 151492 91490
rect 151556 91488 151603 91492
rect 151598 91432 151603 91488
rect 122852 91428 122858 91430
rect 124029 91427 124095 91430
rect 151486 91428 151492 91430
rect 151556 91428 151603 91432
rect 151537 91427 151603 91428
rect 93894 91292 93900 91356
rect 93964 91354 93970 91356
rect 95141 91354 95207 91357
rect 93964 91352 95207 91354
rect 93964 91296 95146 91352
rect 95202 91296 95207 91352
rect 93964 91294 95207 91296
rect 93964 91292 93970 91294
rect 95141 91291 95207 91294
rect 96654 91292 96660 91356
rect 96724 91354 96730 91356
rect 97901 91354 97967 91357
rect 96724 91352 97967 91354
rect 96724 91296 97906 91352
rect 97962 91296 97967 91352
rect 96724 91294 97967 91296
rect 96724 91292 96730 91294
rect 97901 91291 97967 91294
rect 101949 91356 102015 91357
rect 101949 91352 101996 91356
rect 102060 91354 102066 91356
rect 101949 91296 101954 91352
rect 101949 91292 101996 91296
rect 102060 91294 102106 91354
rect 102060 91292 102066 91294
rect 109166 91292 109172 91356
rect 109236 91354 109242 91356
rect 110321 91354 110387 91357
rect 109236 91352 110387 91354
rect 109236 91296 110326 91352
rect 110382 91296 110387 91352
rect 109236 91294 110387 91296
rect 109236 91292 109242 91294
rect 101949 91291 102015 91292
rect 110321 91291 110387 91294
rect 116710 91292 116716 91356
rect 116780 91354 116786 91356
rect 117129 91354 117195 91357
rect 119705 91356 119771 91357
rect 119654 91354 119660 91356
rect 116780 91352 117195 91354
rect 116780 91296 117134 91352
rect 117190 91296 117195 91352
rect 116780 91294 117195 91296
rect 119614 91294 119660 91354
rect 119724 91352 119771 91356
rect 119766 91296 119771 91352
rect 116780 91292 116786 91294
rect 117129 91291 117195 91294
rect 119654 91292 119660 91294
rect 119724 91292 119771 91296
rect 151302 91292 151308 91356
rect 151372 91354 151378 91356
rect 151721 91354 151787 91357
rect 151372 91352 151787 91354
rect 151372 91296 151726 91352
rect 151782 91296 151787 91352
rect 151372 91294 151787 91296
rect 151372 91292 151378 91294
rect 119705 91291 119771 91292
rect 151721 91291 151787 91294
rect 74758 91156 74764 91220
rect 74828 91218 74834 91220
rect 75269 91218 75335 91221
rect 74828 91216 75335 91218
rect 74828 91160 75274 91216
rect 75330 91160 75335 91216
rect 74828 91158 75335 91160
rect 74828 91156 74834 91158
rect 75269 91155 75335 91158
rect 84326 91156 84332 91220
rect 84396 91218 84402 91220
rect 85481 91218 85547 91221
rect 86769 91220 86835 91221
rect 86718 91218 86724 91220
rect 84396 91216 85547 91218
rect 84396 91160 85486 91216
rect 85542 91160 85547 91216
rect 84396 91158 85547 91160
rect 86678 91158 86724 91218
rect 86788 91216 86835 91220
rect 86830 91160 86835 91216
rect 84396 91156 84402 91158
rect 85481 91155 85547 91158
rect 86718 91156 86724 91158
rect 86788 91156 86835 91160
rect 88006 91156 88012 91220
rect 88076 91218 88082 91220
rect 88241 91218 88307 91221
rect 88076 91216 88307 91218
rect 88076 91160 88246 91216
rect 88302 91160 88307 91216
rect 88076 91158 88307 91160
rect 88076 91156 88082 91158
rect 86769 91155 86835 91156
rect 88241 91155 88307 91158
rect 88926 91156 88932 91220
rect 88996 91218 89002 91220
rect 89621 91218 89687 91221
rect 88996 91216 89687 91218
rect 88996 91160 89626 91216
rect 89682 91160 89687 91216
rect 88996 91158 89687 91160
rect 88996 91156 89002 91158
rect 89621 91155 89687 91158
rect 90214 91156 90220 91220
rect 90284 91218 90290 91220
rect 91001 91218 91067 91221
rect 90284 91216 91067 91218
rect 90284 91160 91006 91216
rect 91062 91160 91067 91216
rect 90284 91158 91067 91160
rect 90284 91156 90290 91158
rect 91001 91155 91067 91158
rect 91318 91156 91324 91220
rect 91388 91218 91394 91220
rect 91921 91218 91987 91221
rect 91388 91216 91987 91218
rect 91388 91160 91926 91216
rect 91982 91160 91987 91216
rect 91388 91158 91987 91160
rect 91388 91156 91394 91158
rect 91921 91155 91987 91158
rect 92606 91156 92612 91220
rect 92676 91218 92682 91220
rect 93209 91218 93275 91221
rect 95049 91220 95115 91221
rect 94998 91218 95004 91220
rect 92676 91216 93275 91218
rect 92676 91160 93214 91216
rect 93270 91160 93275 91216
rect 92676 91158 93275 91160
rect 94958 91158 95004 91218
rect 95068 91216 95115 91220
rect 95110 91160 95115 91216
rect 92676 91156 92682 91158
rect 93209 91155 93275 91158
rect 94998 91156 95004 91158
rect 95068 91156 95115 91160
rect 96286 91156 96292 91220
rect 96356 91218 96362 91220
rect 96521 91218 96587 91221
rect 96356 91216 96587 91218
rect 96356 91160 96526 91216
rect 96582 91160 96587 91216
rect 96356 91158 96587 91160
rect 96356 91156 96362 91158
rect 95049 91155 95115 91156
rect 96521 91155 96587 91158
rect 97206 91156 97212 91220
rect 97276 91218 97282 91220
rect 97809 91218 97875 91221
rect 97276 91216 97875 91218
rect 97276 91160 97814 91216
rect 97870 91160 97875 91216
rect 97276 91158 97875 91160
rect 97276 91156 97282 91158
rect 97809 91155 97875 91158
rect 98126 91156 98132 91220
rect 98196 91156 98202 91220
rect 99046 91156 99052 91220
rect 99116 91218 99122 91220
rect 99189 91218 99255 91221
rect 100569 91220 100635 91221
rect 100518 91218 100524 91220
rect 99116 91216 99255 91218
rect 99116 91160 99194 91216
rect 99250 91160 99255 91216
rect 99116 91158 99255 91160
rect 100478 91158 100524 91218
rect 100588 91216 100635 91220
rect 100630 91160 100635 91216
rect 99116 91156 99122 91158
rect 98134 91082 98194 91156
rect 99189 91155 99255 91158
rect 100518 91156 100524 91158
rect 100588 91156 100635 91160
rect 101806 91156 101812 91220
rect 101876 91218 101882 91220
rect 102041 91218 102107 91221
rect 101876 91216 102107 91218
rect 101876 91160 102046 91216
rect 102102 91160 102107 91216
rect 101876 91158 102107 91160
rect 101876 91156 101882 91158
rect 100569 91155 100635 91156
rect 102041 91155 102107 91158
rect 102726 91156 102732 91220
rect 102796 91218 102802 91220
rect 103329 91218 103395 91221
rect 102796 91216 103395 91218
rect 102796 91160 103334 91216
rect 103390 91160 103395 91216
rect 102796 91158 103395 91160
rect 102796 91156 102802 91158
rect 103329 91155 103395 91158
rect 104566 91156 104572 91220
rect 104636 91218 104642 91220
rect 104709 91218 104775 91221
rect 105537 91220 105603 91221
rect 105486 91218 105492 91220
rect 104636 91216 104775 91218
rect 104636 91160 104714 91216
rect 104770 91160 104775 91216
rect 104636 91158 104775 91160
rect 105446 91158 105492 91218
rect 105556 91216 105603 91220
rect 105598 91160 105603 91216
rect 104636 91156 104642 91158
rect 104709 91155 104775 91158
rect 105486 91156 105492 91158
rect 105556 91156 105603 91160
rect 106774 91156 106780 91220
rect 106844 91218 106850 91220
rect 107561 91218 107627 91221
rect 106844 91216 107627 91218
rect 106844 91160 107566 91216
rect 107622 91160 107627 91216
rect 106844 91158 107627 91160
rect 106844 91156 106850 91158
rect 105537 91155 105603 91156
rect 107561 91155 107627 91158
rect 107694 91156 107700 91220
rect 107764 91218 107770 91220
rect 108021 91218 108087 91221
rect 107764 91216 108087 91218
rect 107764 91160 108026 91216
rect 108082 91160 108087 91216
rect 107764 91158 108087 91160
rect 107764 91156 107770 91158
rect 108021 91155 108087 91158
rect 109534 91156 109540 91220
rect 109604 91218 109610 91220
rect 110229 91218 110295 91221
rect 109604 91216 110295 91218
rect 109604 91160 110234 91216
rect 110290 91160 110295 91216
rect 109604 91158 110295 91160
rect 109604 91156 109610 91158
rect 110229 91155 110295 91158
rect 110638 91156 110644 91220
rect 110708 91218 110714 91220
rect 111701 91218 111767 91221
rect 110708 91216 111767 91218
rect 110708 91160 111706 91216
rect 111762 91160 111767 91216
rect 110708 91158 111767 91160
rect 110708 91156 110714 91158
rect 111701 91155 111767 91158
rect 113214 91156 113220 91220
rect 113284 91218 113290 91220
rect 113357 91218 113423 91221
rect 114277 91220 114343 91221
rect 114277 91218 114324 91220
rect 113284 91216 113423 91218
rect 113284 91160 113362 91216
rect 113418 91160 113423 91216
rect 113284 91158 113423 91160
rect 114232 91216 114324 91218
rect 114232 91160 114282 91216
rect 114232 91158 114324 91160
rect 113284 91156 113290 91158
rect 113357 91155 113423 91158
rect 114277 91156 114324 91158
rect 114388 91156 114394 91220
rect 115657 91218 115723 91221
rect 115790 91218 115796 91220
rect 115657 91216 115796 91218
rect 115657 91160 115662 91216
rect 115718 91160 115796 91216
rect 115657 91158 115796 91160
rect 114277 91155 114343 91156
rect 115657 91155 115723 91158
rect 115790 91156 115796 91158
rect 115860 91156 115866 91220
rect 117078 91156 117084 91220
rect 117148 91218 117154 91220
rect 117221 91218 117287 91221
rect 117148 91216 117287 91218
rect 117148 91160 117226 91216
rect 117282 91160 117287 91216
rect 117148 91158 117287 91160
rect 117148 91156 117154 91158
rect 117221 91155 117287 91158
rect 118182 91156 118188 91220
rect 118252 91218 118258 91220
rect 118509 91218 118575 91221
rect 118252 91216 118575 91218
rect 118252 91160 118514 91216
rect 118570 91160 118575 91216
rect 118252 91158 118575 91160
rect 118252 91156 118258 91158
rect 118509 91155 118575 91158
rect 119286 91156 119292 91220
rect 119356 91218 119362 91220
rect 119889 91218 119955 91221
rect 119356 91216 119955 91218
rect 119356 91160 119894 91216
rect 119950 91160 119955 91216
rect 119356 91158 119955 91160
rect 119356 91156 119362 91158
rect 119889 91155 119955 91158
rect 120206 91156 120212 91220
rect 120276 91218 120282 91220
rect 121361 91218 121427 91221
rect 120276 91216 121427 91218
rect 120276 91160 121366 91216
rect 121422 91160 121427 91216
rect 120276 91158 121427 91160
rect 120276 91156 120282 91158
rect 121361 91155 121427 91158
rect 122046 91156 122052 91220
rect 122116 91218 122122 91220
rect 122741 91218 122807 91221
rect 124121 91220 124187 91221
rect 124070 91218 124076 91220
rect 122116 91216 122807 91218
rect 122116 91160 122746 91216
rect 122802 91160 122807 91216
rect 122116 91158 122807 91160
rect 124030 91158 124076 91218
rect 124140 91216 124187 91220
rect 124182 91160 124187 91216
rect 122116 91156 122122 91158
rect 122741 91155 122807 91158
rect 124070 91156 124076 91158
rect 124140 91156 124187 91160
rect 124438 91156 124444 91220
rect 124508 91218 124514 91220
rect 124765 91218 124831 91221
rect 126513 91220 126579 91221
rect 126462 91218 126468 91220
rect 124508 91216 124831 91218
rect 124508 91160 124770 91216
rect 124826 91160 124831 91216
rect 124508 91158 124831 91160
rect 126422 91158 126468 91218
rect 126532 91216 126579 91220
rect 126574 91160 126579 91216
rect 124508 91156 124514 91158
rect 124121 91155 124187 91156
rect 124765 91155 124831 91158
rect 126462 91156 126468 91158
rect 126532 91156 126579 91160
rect 126646 91156 126652 91220
rect 126716 91218 126722 91220
rect 126881 91218 126947 91221
rect 126716 91216 126947 91218
rect 126716 91160 126886 91216
rect 126942 91160 126947 91216
rect 126716 91158 126947 91160
rect 126716 91156 126722 91158
rect 126513 91155 126579 91156
rect 126881 91155 126947 91158
rect 129406 91156 129412 91220
rect 129476 91218 129482 91220
rect 129641 91218 129707 91221
rect 129476 91216 129707 91218
rect 129476 91160 129646 91216
rect 129702 91160 129707 91216
rect 129476 91158 129707 91160
rect 129476 91156 129482 91158
rect 129641 91155 129707 91158
rect 130694 91156 130700 91220
rect 130764 91218 130770 91220
rect 131021 91218 131087 91221
rect 130764 91216 131087 91218
rect 130764 91160 131026 91216
rect 131082 91160 131087 91216
rect 130764 91158 131087 91160
rect 130764 91156 130770 91158
rect 131021 91155 131087 91158
rect 133086 91156 133092 91220
rect 133156 91218 133162 91220
rect 133781 91218 133847 91221
rect 133156 91216 133847 91218
rect 133156 91160 133786 91216
rect 133842 91160 133847 91216
rect 133156 91158 133847 91160
rect 133156 91156 133162 91158
rect 133781 91155 133847 91158
rect 134374 91156 134380 91220
rect 134444 91218 134450 91220
rect 134517 91218 134583 91221
rect 151629 91220 151695 91221
rect 151629 91218 151676 91220
rect 134444 91216 134583 91218
rect 134444 91160 134522 91216
rect 134578 91160 134583 91216
rect 134444 91158 134583 91160
rect 151584 91216 151676 91218
rect 151584 91160 151634 91216
rect 151584 91158 151676 91160
rect 134444 91156 134450 91158
rect 134517 91155 134583 91158
rect 151629 91156 151676 91158
rect 151740 91156 151746 91220
rect 151629 91155 151695 91156
rect 173249 91082 173315 91085
rect 98134 91080 173315 91082
rect 98134 91024 173254 91080
rect 173310 91024 173315 91080
rect 98134 91022 173315 91024
rect 173249 91019 173315 91022
rect 102542 90884 102548 90948
rect 102612 90946 102618 90948
rect 176193 90946 176259 90949
rect 102612 90944 176259 90946
rect 102612 90888 176198 90944
rect 176254 90888 176259 90944
rect 102612 90886 176259 90888
rect 102612 90884 102618 90886
rect 176193 90883 176259 90886
rect 209221 90402 209287 90405
rect 249333 90402 249399 90405
rect 209221 90400 249399 90402
rect 209221 90344 209226 90400
rect 209282 90344 249338 90400
rect 249394 90344 249399 90400
rect 209221 90342 249399 90344
rect 209221 90339 209287 90342
rect 249333 90339 249399 90342
rect 104525 89722 104591 89725
rect 188429 89722 188495 89725
rect 104525 89720 188495 89722
rect 104525 89664 104530 89720
rect 104586 89664 188434 89720
rect 188490 89664 188495 89720
rect 104525 89662 188495 89664
rect 104525 89659 104591 89662
rect 188429 89659 188495 89662
rect 86493 89586 86559 89589
rect 167913 89586 167979 89589
rect 86493 89584 167979 89586
rect 86493 89528 86498 89584
rect 86554 89528 167918 89584
rect 167974 89528 167979 89584
rect 86493 89526 167979 89528
rect 86493 89523 86559 89526
rect 167913 89523 167979 89526
rect 112621 89450 112687 89453
rect 193949 89450 194015 89453
rect 112621 89448 194015 89450
rect 112621 89392 112626 89448
rect 112682 89392 193954 89448
rect 194010 89392 194015 89448
rect 112621 89390 194015 89392
rect 112621 89387 112687 89390
rect 193949 89387 194015 89390
rect 200757 89178 200823 89181
rect 224217 89178 224283 89181
rect 200757 89176 224283 89178
rect 200757 89120 200762 89176
rect 200818 89120 224222 89176
rect 224278 89120 224283 89176
rect 200757 89118 224283 89120
rect 200757 89115 200823 89118
rect 224217 89115 224283 89118
rect 185577 89042 185643 89045
rect 263133 89042 263199 89045
rect 185577 89040 263199 89042
rect 185577 88984 185582 89040
rect 185638 88984 263138 89040
rect 263194 88984 263199 89040
rect 185577 88982 263199 88984
rect 185577 88979 185643 88982
rect 263133 88979 263199 88982
rect 75269 88226 75335 88229
rect 187969 88226 188035 88229
rect 75269 88224 188035 88226
rect 75269 88168 75274 88224
rect 75330 88168 187974 88224
rect 188030 88168 188035 88224
rect 75269 88166 188035 88168
rect 75269 88163 75335 88166
rect 187969 88163 188035 88166
rect 108021 88090 108087 88093
rect 189809 88090 189875 88093
rect 108021 88088 189875 88090
rect 108021 88032 108026 88088
rect 108082 88032 189814 88088
rect 189870 88032 189875 88088
rect 108021 88030 189875 88032
rect 108021 88027 108087 88030
rect 189809 88027 189875 88030
rect 113357 87954 113423 87957
rect 169017 87954 169083 87957
rect 113357 87952 169083 87954
rect 113357 87896 113362 87952
rect 113418 87896 169022 87952
rect 169078 87896 169083 87952
rect 113357 87894 169083 87896
rect 113357 87891 113423 87894
rect 169017 87891 169083 87894
rect 196709 87546 196775 87549
rect 280153 87546 280219 87549
rect 196709 87544 280219 87546
rect 196709 87488 196714 87544
rect 196770 87488 280158 87544
rect 280214 87488 280219 87544
rect 196709 87486 280219 87488
rect 196709 87483 196775 87486
rect 280153 87483 280219 87486
rect 67265 86866 67331 86869
rect 214833 86866 214899 86869
rect 67265 86864 214899 86866
rect 67265 86808 67270 86864
rect 67326 86808 214838 86864
rect 214894 86808 214899 86864
rect 67265 86806 214899 86808
rect 67265 86803 67331 86806
rect 214833 86803 214899 86806
rect 91921 86730 91987 86733
rect 184473 86730 184539 86733
rect 91921 86728 184539 86730
rect 91921 86672 91926 86728
rect 91982 86672 184478 86728
rect 184534 86672 184539 86728
rect 91921 86670 184539 86672
rect 91921 86667 91987 86670
rect 184473 86667 184539 86670
rect 124765 86594 124831 86597
rect 184657 86594 184723 86597
rect 124765 86592 184723 86594
rect 124765 86536 124770 86592
rect 124826 86536 184662 86592
rect 184718 86536 184723 86592
rect 124765 86534 184723 86536
rect 124765 86531 124831 86534
rect 184657 86531 184723 86534
rect 204897 86186 204963 86189
rect 252093 86186 252159 86189
rect 204897 86184 252159 86186
rect 204897 86128 204902 86184
rect 204958 86128 252098 86184
rect 252154 86128 252159 86184
rect 204897 86126 252159 86128
rect 204897 86123 204963 86126
rect 252093 86123 252159 86126
rect 582465 86186 582531 86189
rect 583520 86186 584960 86276
rect 582465 86184 584960 86186
rect 582465 86128 582470 86184
rect 582526 86128 584960 86184
rect 582465 86126 584960 86128
rect 582465 86123 582531 86126
rect 583520 86036 584960 86126
rect 65977 85506 66043 85509
rect 213453 85506 213519 85509
rect 65977 85504 213519 85506
rect 65977 85448 65982 85504
rect 66038 85448 213458 85504
rect 213514 85448 213519 85504
rect 65977 85446 213519 85448
rect 65977 85443 66043 85446
rect 213453 85443 213519 85446
rect 101949 85370 102015 85373
rect 171777 85370 171843 85373
rect 101949 85368 171843 85370
rect 101949 85312 101954 85368
rect 102010 85312 171782 85368
rect 171838 85312 171843 85368
rect 101949 85310 171843 85312
rect 101949 85307 102015 85310
rect 171777 85307 171843 85310
rect 134517 85234 134583 85237
rect 164969 85234 165035 85237
rect 134517 85232 165035 85234
rect 134517 85176 134522 85232
rect 134578 85176 164974 85232
rect 165030 85176 165035 85232
rect 134517 85174 165035 85176
rect 134517 85171 134583 85174
rect 164969 85171 165035 85174
rect 202229 84826 202295 84829
rect 270493 84826 270559 84829
rect 202229 84824 270559 84826
rect -960 84690 480 84780
rect 202229 84768 202234 84824
rect 202290 84768 270498 84824
rect 270554 84768 270559 84824
rect 202229 84766 270559 84768
rect 202229 84763 202295 84766
rect 270493 84763 270559 84766
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 135897 84146 135963 84149
rect 203701 84146 203767 84149
rect 135897 84144 203767 84146
rect 135897 84088 135902 84144
rect 135958 84088 203706 84144
rect 203762 84088 203767 84144
rect 135897 84086 203767 84088
rect 135897 84083 135963 84086
rect 203701 84083 203767 84086
rect 115197 84010 115263 84013
rect 166390 84010 166396 84012
rect 115197 84008 166396 84010
rect 115197 83952 115202 84008
rect 115258 83952 166396 84008
rect 115197 83950 166396 83952
rect 115197 83947 115263 83950
rect 166390 83948 166396 83950
rect 166460 83948 166466 84012
rect 30281 83466 30347 83469
rect 260373 83466 260439 83469
rect 30281 83464 260439 83466
rect 30281 83408 30286 83464
rect 30342 83408 260378 83464
rect 260434 83408 260439 83464
rect 30281 83406 260439 83408
rect 30281 83403 30347 83406
rect 260373 83403 260439 83406
rect 88241 82786 88307 82789
rect 169109 82786 169175 82789
rect 88241 82784 169175 82786
rect 88241 82728 88246 82784
rect 88302 82728 169114 82784
rect 169170 82728 169175 82784
rect 88241 82726 169175 82728
rect 88241 82723 88307 82726
rect 169109 82723 169175 82726
rect 126881 82650 126947 82653
rect 171869 82650 171935 82653
rect 126881 82648 171935 82650
rect 126881 82592 126886 82648
rect 126942 82592 171874 82648
rect 171930 82592 171935 82648
rect 126881 82590 171935 82592
rect 126881 82587 126947 82590
rect 171869 82587 171935 82590
rect 175917 82242 175983 82245
rect 273253 82242 273319 82245
rect 175917 82240 273319 82242
rect 175917 82184 175922 82240
rect 175978 82184 273258 82240
rect 273314 82184 273319 82240
rect 175917 82182 273319 82184
rect 175917 82179 175983 82182
rect 273253 82179 273319 82182
rect 41229 82106 41295 82109
rect 263041 82106 263107 82109
rect 41229 82104 263107 82106
rect 41229 82048 41234 82104
rect 41290 82048 263046 82104
rect 263102 82048 263107 82104
rect 41229 82046 263107 82048
rect 41229 82043 41295 82046
rect 263041 82043 263107 82046
rect 108297 81426 108363 81429
rect 168966 81426 168972 81428
rect 108297 81424 168972 81426
rect 108297 81368 108302 81424
rect 108358 81368 168972 81424
rect 108297 81366 168972 81368
rect 108297 81363 108363 81366
rect 168966 81364 168972 81366
rect 169036 81364 169042 81428
rect 117037 80882 117103 80885
rect 264329 80882 264395 80885
rect 117037 80880 264395 80882
rect 117037 80824 117042 80880
rect 117098 80824 264334 80880
rect 264390 80824 264395 80880
rect 117037 80822 264395 80824
rect 117037 80819 117103 80822
rect 264329 80819 264395 80822
rect 12341 80746 12407 80749
rect 256141 80746 256207 80749
rect 12341 80744 256207 80746
rect 12341 80688 12346 80744
rect 12402 80688 256146 80744
rect 256202 80688 256207 80744
rect 12341 80686 256207 80688
rect 12341 80683 12407 80686
rect 256141 80683 256207 80686
rect 97901 80066 97967 80069
rect 185761 80066 185827 80069
rect 97901 80064 185827 80066
rect 97901 80008 97906 80064
rect 97962 80008 185766 80064
rect 185822 80008 185827 80064
rect 97901 80006 185827 80008
rect 97901 80003 97967 80006
rect 185761 80003 185827 80006
rect 5441 79522 5507 79525
rect 246481 79522 246547 79525
rect 5441 79520 246547 79522
rect 5441 79464 5446 79520
rect 5502 79464 246486 79520
rect 246542 79464 246547 79520
rect 5441 79462 246547 79464
rect 5441 79459 5507 79462
rect 246481 79459 246547 79462
rect 15837 79386 15903 79389
rect 265893 79386 265959 79389
rect 15837 79384 265959 79386
rect 15837 79328 15842 79384
rect 15898 79328 265898 79384
rect 265954 79328 265959 79384
rect 15837 79326 265959 79328
rect 15837 79323 15903 79326
rect 265893 79323 265959 79326
rect 89621 78570 89687 78573
rect 211889 78570 211955 78573
rect 89621 78568 211955 78570
rect 89621 78512 89626 78568
rect 89682 78512 211894 78568
rect 211950 78512 211955 78568
rect 89621 78510 211955 78512
rect 89621 78507 89687 78510
rect 211889 78507 211955 78510
rect 111057 78434 111123 78437
rect 177573 78434 177639 78437
rect 111057 78432 177639 78434
rect 111057 78376 111062 78432
rect 111118 78376 177578 78432
rect 177634 78376 177639 78432
rect 111057 78374 177639 78376
rect 111057 78371 111123 78374
rect 177573 78371 177639 78374
rect 13721 77890 13787 77893
rect 258901 77890 258967 77893
rect 13721 77888 258967 77890
rect 13721 77832 13726 77888
rect 13782 77832 258906 77888
rect 258962 77832 258967 77888
rect 13721 77830 258967 77832
rect 13721 77827 13787 77830
rect 258901 77827 258967 77830
rect 106181 76666 106247 76669
rect 257521 76666 257587 76669
rect 106181 76664 257587 76666
rect 106181 76608 106186 76664
rect 106242 76608 257526 76664
rect 257582 76608 257587 76664
rect 106181 76606 257587 76608
rect 106181 76603 106247 76606
rect 257521 76603 257587 76606
rect 43989 76530 44055 76533
rect 238109 76530 238175 76533
rect 43989 76528 238175 76530
rect 43989 76472 43994 76528
rect 44050 76472 238114 76528
rect 238170 76472 238175 76528
rect 43989 76470 238175 76472
rect 43989 76467 44055 76470
rect 238109 76467 238175 76470
rect 73061 75306 73127 75309
rect 241053 75306 241119 75309
rect 73061 75304 241119 75306
rect 73061 75248 73066 75304
rect 73122 75248 241058 75304
rect 241114 75248 241119 75304
rect 73061 75246 241119 75248
rect 73061 75243 73127 75246
rect 241053 75243 241119 75246
rect 19241 75170 19307 75173
rect 234153 75170 234219 75173
rect 19241 75168 234219 75170
rect 19241 75112 19246 75168
rect 19302 75112 234158 75168
rect 234214 75112 234219 75168
rect 19241 75110 234219 75112
rect 19241 75107 19307 75110
rect 234153 75107 234219 75110
rect 106917 74490 106983 74493
rect 171961 74490 172027 74493
rect 106917 74488 172027 74490
rect 106917 74432 106922 74488
rect 106978 74432 171966 74488
rect 172022 74432 172027 74488
rect 106917 74430 172027 74432
rect 106917 74427 106983 74430
rect 171961 74427 172027 74430
rect 71037 73946 71103 73949
rect 261753 73946 261819 73949
rect 71037 73944 261819 73946
rect 71037 73888 71042 73944
rect 71098 73888 261758 73944
rect 261814 73888 261819 73944
rect 71037 73886 261819 73888
rect 71037 73883 71103 73886
rect 261753 73883 261819 73886
rect 23381 73810 23447 73813
rect 249241 73810 249307 73813
rect 23381 73808 249307 73810
rect 23381 73752 23386 73808
rect 23442 73752 249246 73808
rect 249302 73752 249307 73808
rect 23381 73750 249307 73752
rect 23381 73747 23447 73750
rect 249241 73747 249307 73750
rect 583753 73266 583819 73269
rect 583710 73264 583819 73266
rect 583710 73208 583758 73264
rect 583814 73208 583819 73264
rect 583710 73203 583819 73208
rect 104157 73130 104223 73133
rect 191189 73130 191255 73133
rect 583710 73130 583770 73203
rect 104157 73128 191255 73130
rect 104157 73072 104162 73128
rect 104218 73072 191194 73128
rect 191250 73072 191255 73128
rect 104157 73070 191255 73072
rect 104157 73067 104223 73070
rect 191189 73067 191255 73070
rect 583342 73084 583770 73130
rect 583342 73070 584960 73084
rect 583342 72994 583402 73070
rect 583520 72994 584960 73070
rect 583342 72934 584960 72994
rect 583520 72844 584960 72934
rect 50889 72586 50955 72589
rect 262806 72586 262812 72588
rect 50889 72584 262812 72586
rect 50889 72528 50894 72584
rect 50950 72528 262812 72584
rect 50889 72526 262812 72528
rect 50889 72523 50955 72526
rect 262806 72524 262812 72526
rect 262876 72524 262882 72588
rect 41137 72450 41203 72453
rect 284293 72450 284359 72453
rect 41137 72448 284359 72450
rect 41137 72392 41142 72448
rect 41198 72392 284298 72448
rect 284354 72392 284359 72448
rect 41137 72390 284359 72392
rect 41137 72387 41203 72390
rect 284293 72387 284359 72390
rect -960 71634 480 71724
rect 3417 71634 3483 71637
rect -960 71632 3483 71634
rect -960 71576 3422 71632
rect 3478 71576 3483 71632
rect -960 71574 3483 71576
rect -960 71484 480 71574
rect 3417 71571 3483 71574
rect 104801 71226 104867 71229
rect 264421 71226 264487 71229
rect 104801 71224 264487 71226
rect 104801 71168 104806 71224
rect 104862 71168 264426 71224
rect 264482 71168 264487 71224
rect 104801 71166 264487 71168
rect 104801 71163 104867 71166
rect 264421 71163 264487 71166
rect 60641 71090 60707 71093
rect 248413 71090 248479 71093
rect 60641 71088 248479 71090
rect 60641 71032 60646 71088
rect 60702 71032 248418 71088
rect 248474 71032 248479 71088
rect 60641 71030 248479 71032
rect 60641 71027 60707 71030
rect 248413 71027 248479 71030
rect 56501 69730 56567 69733
rect 262213 69730 262279 69733
rect 56501 69728 262279 69730
rect 56501 69672 56506 69728
rect 56562 69672 262218 69728
rect 262274 69672 262279 69728
rect 56501 69670 262279 69672
rect 56501 69667 56567 69670
rect 262213 69667 262279 69670
rect 35801 69594 35867 69597
rect 242341 69594 242407 69597
rect 35801 69592 242407 69594
rect 35801 69536 35806 69592
rect 35862 69536 242346 69592
rect 242402 69536 242407 69592
rect 35801 69534 242407 69536
rect 35801 69531 35867 69534
rect 242341 69531 242407 69534
rect 64781 68370 64847 68373
rect 249057 68370 249123 68373
rect 64781 68368 249123 68370
rect 64781 68312 64786 68368
rect 64842 68312 249062 68368
rect 249118 68312 249123 68368
rect 64781 68310 249123 68312
rect 64781 68307 64847 68310
rect 249057 68307 249123 68310
rect 26141 68234 26207 68237
rect 256233 68234 256299 68237
rect 26141 68232 256299 68234
rect 26141 68176 26146 68232
rect 26202 68176 256238 68232
rect 256294 68176 256299 68232
rect 26141 68174 256299 68176
rect 26141 68171 26207 68174
rect 256233 68171 256299 68174
rect 160737 67146 160803 67149
rect 214741 67146 214807 67149
rect 160737 67144 214807 67146
rect 160737 67088 160742 67144
rect 160798 67088 214746 67144
rect 214802 67088 214807 67144
rect 160737 67086 214807 67088
rect 160737 67083 160803 67086
rect 214741 67083 214807 67086
rect 94957 67010 95023 67013
rect 250529 67010 250595 67013
rect 94957 67008 250595 67010
rect 94957 66952 94962 67008
rect 95018 66952 250534 67008
rect 250590 66952 250595 67008
rect 94957 66950 250595 66952
rect 94957 66947 95023 66950
rect 250529 66947 250595 66950
rect 15101 66874 15167 66877
rect 258574 66874 258580 66876
rect 15101 66872 258580 66874
rect 15101 66816 15106 66872
rect 15162 66816 258580 66872
rect 15101 66814 258580 66816
rect 15101 66811 15167 66814
rect 258574 66812 258580 66814
rect 258644 66812 258650 66876
rect 68921 65650 68987 65653
rect 247677 65650 247743 65653
rect 68921 65648 247743 65650
rect 68921 65592 68926 65648
rect 68982 65592 247682 65648
rect 247738 65592 247743 65648
rect 68921 65590 247743 65592
rect 68921 65587 68987 65590
rect 247677 65587 247743 65590
rect 63401 65514 63467 65517
rect 276013 65514 276079 65517
rect 63401 65512 276079 65514
rect 63401 65456 63406 65512
rect 63462 65456 276018 65512
rect 276074 65456 276079 65512
rect 63401 65454 276079 65456
rect 63401 65451 63467 65454
rect 276013 65451 276079 65454
rect 120073 64290 120139 64293
rect 225597 64290 225663 64293
rect 120073 64288 225663 64290
rect 120073 64232 120078 64288
rect 120134 64232 225602 64288
rect 225658 64232 225663 64288
rect 120073 64230 225663 64232
rect 120073 64227 120139 64230
rect 225597 64227 225663 64230
rect 75821 64154 75887 64157
rect 257337 64154 257403 64157
rect 75821 64152 257403 64154
rect 75821 64096 75826 64152
rect 75882 64096 257342 64152
rect 257398 64096 257403 64152
rect 75821 64094 257403 64096
rect 75821 64091 75887 64094
rect 257337 64091 257403 64094
rect 33041 62794 33107 62797
rect 253054 62794 253060 62796
rect 33041 62792 253060 62794
rect 33041 62736 33046 62792
rect 33102 62736 253060 62792
rect 33041 62734 253060 62736
rect 33041 62731 33107 62734
rect 253054 62732 253060 62734
rect 253124 62732 253130 62796
rect 87597 61434 87663 61437
rect 265617 61434 265683 61437
rect 87597 61432 265683 61434
rect 87597 61376 87602 61432
rect 87658 61376 265622 61432
rect 265678 61376 265683 61432
rect 87597 61374 265683 61376
rect 87597 61371 87663 61374
rect 265617 61371 265683 61374
rect 20529 59938 20595 59941
rect 246297 59938 246363 59941
rect 20529 59936 246363 59938
rect 20529 59880 20534 59936
rect 20590 59880 246302 59936
rect 246358 59880 246363 59936
rect 20529 59878 246363 59880
rect 20529 59875 20595 59878
rect 246297 59875 246363 59878
rect 580257 59666 580323 59669
rect 583520 59666 584960 59756
rect 580257 59664 584960 59666
rect 580257 59608 580262 59664
rect 580318 59608 584960 59664
rect 580257 59606 584960 59608
rect 580257 59603 580323 59606
rect 583520 59516 584960 59606
rect 32397 58714 32463 58717
rect 120073 58714 120139 58717
rect 32397 58712 120139 58714
rect -960 58578 480 58668
rect 32397 58656 32402 58712
rect 32458 58656 120078 58712
rect 120134 58656 120139 58712
rect 32397 58654 120139 58656
rect 32397 58651 32463 58654
rect 120073 58651 120139 58654
rect 3049 58578 3115 58581
rect -960 58576 3115 58578
rect -960 58520 3054 58576
rect 3110 58520 3115 58576
rect -960 58518 3115 58520
rect -960 58428 480 58518
rect 3049 58515 3115 58518
rect 89621 58578 89687 58581
rect 262949 58578 263015 58581
rect 89621 58576 263015 58578
rect 89621 58520 89626 58576
rect 89682 58520 262954 58576
rect 263010 58520 263015 58576
rect 89621 58518 263015 58520
rect 89621 58515 89687 58518
rect 262949 58515 263015 58518
rect 57830 57156 57836 57220
rect 57900 57218 57906 57220
rect 347037 57218 347103 57221
rect 57900 57216 347103 57218
rect 57900 57160 347042 57216
rect 347098 57160 347103 57216
rect 57900 57158 347103 57160
rect 57900 57156 57906 57158
rect 347037 57155 347103 57158
rect 17861 55858 17927 55861
rect 260046 55858 260052 55860
rect 17861 55856 260052 55858
rect 17861 55800 17866 55856
rect 17922 55800 260052 55856
rect 17861 55798 260052 55800
rect 17861 55795 17927 55798
rect 260046 55796 260052 55798
rect 260116 55796 260122 55860
rect 53649 54498 53715 54501
rect 261569 54498 261635 54501
rect 53649 54496 261635 54498
rect 53649 54440 53654 54496
rect 53710 54440 261574 54496
rect 261630 54440 261635 54496
rect 53649 54438 261635 54440
rect 53649 54435 53715 54438
rect 261569 54435 261635 54438
rect 57881 53138 57947 53141
rect 232589 53138 232655 53141
rect 57881 53136 232655 53138
rect 57881 53080 57886 53136
rect 57942 53080 232594 53136
rect 232650 53080 232655 53136
rect 57881 53078 232655 53080
rect 57881 53075 57947 53078
rect 232589 53075 232655 53078
rect 108941 51914 109007 51917
rect 247769 51914 247835 51917
rect 108941 51912 247835 51914
rect 108941 51856 108946 51912
rect 109002 51856 247774 51912
rect 247830 51856 247835 51912
rect 108941 51854 247835 51856
rect 108941 51851 109007 51854
rect 247769 51851 247835 51854
rect 10961 51778 11027 51781
rect 230974 51778 230980 51780
rect 10961 51776 230980 51778
rect 10961 51720 10966 51776
rect 11022 51720 230980 51776
rect 10961 51718 230980 51720
rect 10961 51715 11027 51718
rect 230974 51716 230980 51718
rect 231044 51716 231050 51780
rect 38561 50282 38627 50285
rect 238017 50282 238083 50285
rect 38561 50280 238083 50282
rect 38561 50224 38566 50280
rect 38622 50224 238022 50280
rect 238078 50224 238083 50280
rect 38561 50222 238083 50224
rect 38561 50219 38627 50222
rect 238017 50219 238083 50222
rect 37181 48922 37247 48925
rect 266854 48922 266860 48924
rect 37181 48920 266860 48922
rect 37181 48864 37186 48920
rect 37242 48864 266860 48920
rect 37181 48862 266860 48864
rect 37181 48859 37247 48862
rect 266854 48860 266860 48862
rect 266924 48860 266930 48924
rect 582833 46338 582899 46341
rect 583520 46338 584960 46428
rect 582833 46336 584960 46338
rect 582833 46280 582838 46336
rect 582894 46280 584960 46336
rect 582833 46278 584960 46280
rect 582833 46275 582899 46278
rect 180057 46202 180123 46205
rect 238017 46202 238083 46205
rect 180057 46200 238083 46202
rect 180057 46144 180062 46200
rect 180118 46144 238022 46200
rect 238078 46144 238083 46200
rect 583520 46188 584960 46278
rect 180057 46142 238083 46144
rect 180057 46139 180123 46142
rect 238017 46139 238083 46142
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 135253 43482 135319 43485
rect 169702 43482 169708 43484
rect 135253 43480 169708 43482
rect 135253 43424 135258 43480
rect 135314 43424 169708 43480
rect 135253 43422 169708 43424
rect 135253 43419 135319 43422
rect 169702 43420 169708 43422
rect 169772 43420 169778 43484
rect 180057 43482 180123 43485
rect 227069 43482 227135 43485
rect 180057 43480 227135 43482
rect 180057 43424 180062 43480
rect 180118 43424 227074 43480
rect 227130 43424 227135 43480
rect 180057 43422 227135 43424
rect 180057 43419 180123 43422
rect 227069 43419 227135 43422
rect 189717 42122 189783 42125
rect 240133 42122 240199 42125
rect 189717 42120 240199 42122
rect 189717 42064 189722 42120
rect 189778 42064 240138 42120
rect 240194 42064 240199 42120
rect 189717 42062 240199 42064
rect 189717 42059 189783 42062
rect 240133 42059 240199 42062
rect 70209 39402 70275 39405
rect 240726 39402 240732 39404
rect 70209 39400 240732 39402
rect 70209 39344 70214 39400
rect 70270 39344 240732 39400
rect 70209 39342 240732 39344
rect 70209 39339 70275 39342
rect 240726 39340 240732 39342
rect 240796 39340 240802 39404
rect 24761 39266 24827 39269
rect 264094 39266 264100 39268
rect 24761 39264 264100 39266
rect 24761 39208 24766 39264
rect 24822 39208 264100 39264
rect 24761 39206 264100 39208
rect 24761 39203 24827 39206
rect 264094 39204 264100 39206
rect 264164 39204 264170 39268
rect 180241 37906 180307 37909
rect 292573 37906 292639 37909
rect 180241 37904 292639 37906
rect 180241 37848 180246 37904
rect 180302 37848 292578 37904
rect 292634 37848 292639 37904
rect 180241 37846 292639 37848
rect 180241 37843 180307 37846
rect 292573 37843 292639 37846
rect 182817 35186 182883 35189
rect 258073 35186 258139 35189
rect 182817 35184 258139 35186
rect 182817 35128 182822 35184
rect 182878 35128 258078 35184
rect 258134 35128 258139 35184
rect 182817 35126 258139 35128
rect 182817 35123 182883 35126
rect 258073 35123 258139 35126
rect 582741 33146 582807 33149
rect 583520 33146 584960 33236
rect 582741 33144 584960 33146
rect 582741 33088 582746 33144
rect 582802 33088 584960 33144
rect 582741 33086 584960 33088
rect 582741 33083 582807 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 3141 32466 3207 32469
rect -960 32464 3207 32466
rect -960 32408 3146 32464
rect 3202 32408 3207 32464
rect -960 32406 3207 32408
rect -960 32316 480 32406
rect 3141 32403 3207 32406
rect 198181 30970 198247 30973
rect 263593 30970 263659 30973
rect 198181 30968 263659 30970
rect 198181 30912 198186 30968
rect 198242 30912 263598 30968
rect 263654 30912 263659 30968
rect 198181 30910 263659 30912
rect 198181 30907 198247 30910
rect 263593 30907 263659 30910
rect 192477 28250 192543 28253
rect 264973 28250 265039 28253
rect 192477 28248 265039 28250
rect 192477 28192 192482 28248
rect 192538 28192 264978 28248
rect 265034 28192 265039 28248
rect 192477 28190 265039 28192
rect 192477 28187 192543 28190
rect 264973 28187 265039 28190
rect 28901 26890 28967 26893
rect 267774 26890 267780 26892
rect 28901 26888 267780 26890
rect 28901 26832 28906 26888
rect 28962 26832 267780 26888
rect 28901 26830 267780 26832
rect 28901 26827 28967 26830
rect 267774 26828 267780 26830
rect 267844 26828 267850 26892
rect 3969 25530 4035 25533
rect 237966 25530 237972 25532
rect 3969 25528 237972 25530
rect 3969 25472 3974 25528
rect 4030 25472 237972 25528
rect 3969 25470 237972 25472
rect 3969 25467 4035 25470
rect 237966 25468 237972 25470
rect 238036 25468 238042 25532
rect 105 24170 171 24173
rect 227662 24170 227668 24172
rect 105 24168 227668 24170
rect 105 24112 110 24168
rect 166 24112 227668 24168
rect 105 24110 227668 24112
rect 105 24107 171 24110
rect 227662 24108 227668 24110
rect 227732 24108 227738 24172
rect 173014 22748 173020 22812
rect 173084 22810 173090 22812
rect 280797 22810 280863 22813
rect 173084 22808 280863 22810
rect 173084 22752 280802 22808
rect 280858 22752 280863 22808
rect 173084 22750 280863 22752
rect 173084 22748 173090 22750
rect 280797 22747 280863 22750
rect 59261 22674 59327 22677
rect 307845 22674 307911 22677
rect 59261 22672 307911 22674
rect 59261 22616 59266 22672
rect 59322 22616 307850 22672
rect 307906 22616 307911 22672
rect 59261 22614 307911 22616
rect 59261 22611 59327 22614
rect 307845 22611 307911 22614
rect 28809 21314 28875 21317
rect 262070 21314 262076 21316
rect 28809 21312 262076 21314
rect 28809 21256 28814 21312
rect 28870 21256 262076 21312
rect 28809 21254 262076 21256
rect 28809 21251 28875 21254
rect 262070 21252 262076 21254
rect 262140 21252 262146 21316
rect 583661 20362 583727 20365
rect 583526 20360 583727 20362
rect 583526 20304 583666 20360
rect 583722 20304 583727 20360
rect 583526 20302 583727 20304
rect 67766 19892 67772 19956
rect 67836 19954 67842 19956
rect 255313 19954 255379 19957
rect 583526 19954 583586 20302
rect 583661 20299 583727 20302
rect 67836 19952 255379 19954
rect 67836 19896 255318 19952
rect 255374 19896 255379 19952
rect 67836 19894 255379 19896
rect 67836 19892 67842 19894
rect 255313 19891 255379 19894
rect 583342 19908 583586 19954
rect 583342 19894 584960 19908
rect 583342 19818 583402 19894
rect 583520 19818 584960 19894
rect 583342 19758 584960 19818
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 55029 17234 55095 17237
rect 317413 17234 317479 17237
rect 55029 17232 317479 17234
rect 55029 17176 55034 17232
rect 55090 17176 317418 17232
rect 317474 17176 317479 17232
rect 55029 17174 317479 17176
rect 55029 17171 55095 17174
rect 317413 17171 317479 17174
rect 45277 15874 45343 15877
rect 168414 15874 168420 15876
rect 45277 15872 168420 15874
rect 45277 15816 45282 15872
rect 45338 15816 168420 15872
rect 45277 15814 168420 15816
rect 45277 15811 45343 15814
rect 168414 15812 168420 15814
rect 168484 15812 168490 15876
rect 195094 14452 195100 14516
rect 195164 14514 195170 14516
rect 268377 14514 268443 14517
rect 195164 14512 268443 14514
rect 195164 14456 268382 14512
rect 268438 14456 268443 14512
rect 195164 14454 268443 14456
rect 195164 14452 195170 14454
rect 268377 14451 268443 14454
rect 132953 13018 133019 13021
rect 166942 13018 166948 13020
rect 132953 13016 166948 13018
rect 132953 12960 132958 13016
rect 133014 12960 166948 13016
rect 132953 12958 166948 12960
rect 132953 12955 133019 12958
rect 166942 12956 166948 12958
rect 167012 12956 167018 13020
rect 188286 12956 188292 13020
rect 188356 13018 188362 13020
rect 261753 13018 261819 13021
rect 188356 13016 261819 13018
rect 188356 12960 261758 13016
rect 261814 12960 261819 13016
rect 188356 12958 261819 12960
rect 188356 12956 188362 12958
rect 261753 12955 261819 12958
rect 66110 11596 66116 11660
rect 66180 11658 66186 11660
rect 251173 11658 251239 11661
rect 66180 11656 251239 11658
rect 66180 11600 251178 11656
rect 251234 11600 251239 11656
rect 66180 11598 251239 11600
rect 66180 11596 66186 11598
rect 251173 11595 251239 11598
rect 193857 10298 193923 10301
rect 259453 10298 259519 10301
rect 193857 10296 259519 10298
rect 193857 10240 193862 10296
rect 193918 10240 259458 10296
rect 259514 10240 259519 10296
rect 193857 10238 259519 10240
rect 193857 10235 193923 10238
rect 259453 10235 259519 10238
rect 60825 8938 60891 8941
rect 206277 8938 206343 8941
rect 60825 8936 206343 8938
rect 60825 8880 60830 8936
rect 60886 8880 206282 8936
rect 206338 8880 206343 8936
rect 60825 8878 206343 8880
rect 60825 8875 60891 8878
rect 206277 8875 206343 8878
rect 41873 7714 41939 7717
rect 223614 7714 223620 7716
rect 41873 7712 223620 7714
rect 41873 7656 41878 7712
rect 41934 7656 223620 7712
rect 41873 7654 223620 7656
rect 41873 7651 41939 7654
rect 223614 7652 223620 7654
rect 223684 7652 223690 7716
rect 66713 7578 66779 7581
rect 250294 7578 250300 7580
rect 66713 7576 250300 7578
rect 66713 7520 66718 7576
rect 66774 7520 250300 7576
rect 66713 7518 250300 7520
rect 66713 7515 66779 7518
rect 250294 7516 250300 7518
rect 250364 7516 250370 7580
rect 13 6762 79 6765
rect 13 6760 122 6762
rect 13 6704 18 6760
rect 74 6704 122 6760
rect 13 6699 122 6704
rect 62 6626 122 6699
rect 582649 6626 582715 6629
rect 583520 6626 584960 6716
rect 62 6580 674 6626
rect -960 6566 674 6580
rect -960 6490 480 6566
rect 614 6490 674 6566
rect 582649 6624 584960 6626
rect 582649 6568 582654 6624
rect 582710 6568 584960 6624
rect 582649 6566 584960 6568
rect 582649 6563 582715 6566
rect -960 6430 674 6490
rect 583520 6476 584960 6566
rect -960 6340 480 6430
rect 73797 4858 73863 4861
rect 236637 4858 236703 4861
rect 73797 4856 236703 4858
rect 73797 4800 73802 4856
rect 73858 4800 236642 4856
rect 236698 4800 236703 4856
rect 73797 4798 236703 4800
rect 73797 4795 73863 4798
rect 236637 4795 236703 4798
rect 302734 4796 302740 4860
rect 302804 4858 302810 4860
rect 313825 4858 313891 4861
rect 302804 4856 313891 4858
rect 302804 4800 313830 4856
rect 313886 4800 313891 4856
rect 302804 4798 313891 4800
rect 302804 4796 302810 4798
rect 313825 4795 313891 4798
rect 295926 3980 295932 4044
rect 295996 4042 296002 4044
rect 298461 4042 298527 4045
rect 295996 4040 298527 4042
rect 295996 3984 298466 4040
rect 298522 3984 298527 4040
rect 295996 3982 298527 3984
rect 295996 3980 296002 3982
rect 298461 3979 298527 3982
rect 294873 3906 294939 3909
rect 298134 3906 298140 3908
rect 294873 3904 298140 3906
rect 294873 3848 294878 3904
rect 294934 3848 298140 3904
rect 294873 3846 298140 3848
rect 294873 3843 294939 3846
rect 298134 3844 298140 3846
rect 298204 3844 298210 3908
rect 246389 3634 246455 3637
rect 238710 3632 246455 3634
rect 238710 3576 246394 3632
rect 246450 3576 246455 3632
rect 238710 3574 246455 3576
rect 85665 3498 85731 3501
rect 124857 3498 124923 3501
rect 85665 3496 124923 3498
rect 85665 3440 85670 3496
rect 85726 3440 124862 3496
rect 124918 3440 124923 3496
rect 85665 3438 124923 3440
rect 85665 3435 85731 3438
rect 124857 3435 124923 3438
rect 125869 3498 125935 3501
rect 191097 3498 191163 3501
rect 125869 3496 191163 3498
rect 125869 3440 125874 3496
rect 125930 3440 191102 3496
rect 191158 3440 191163 3496
rect 125869 3438 191163 3440
rect 125869 3435 125935 3438
rect 191097 3435 191163 3438
rect 196617 3498 196683 3501
rect 238710 3498 238770 3574
rect 246389 3571 246455 3574
rect 251766 3572 251772 3636
rect 251836 3634 251842 3636
rect 251836 3574 252570 3634
rect 251836 3572 251842 3574
rect 196617 3496 238770 3498
rect 196617 3440 196622 3496
rect 196678 3440 238770 3496
rect 196617 3438 238770 3440
rect 196617 3435 196683 3438
rect 246246 3436 246252 3500
rect 246316 3498 246322 3500
rect 247585 3498 247651 3501
rect 246316 3496 247651 3498
rect 246316 3440 247590 3496
rect 247646 3440 247651 3496
rect 246316 3438 247651 3440
rect 246316 3436 246322 3438
rect 247585 3435 247651 3438
rect 249006 3436 249012 3500
rect 249076 3498 249082 3500
rect 252369 3498 252435 3501
rect 249076 3496 252435 3498
rect 249076 3440 252374 3496
rect 252430 3440 252435 3496
rect 249076 3438 252435 3440
rect 252510 3498 252570 3574
rect 255814 3572 255820 3636
rect 255884 3634 255890 3636
rect 266537 3634 266603 3637
rect 255884 3632 266603 3634
rect 255884 3576 266542 3632
rect 266598 3576 266603 3632
rect 255884 3574 266603 3576
rect 255884 3572 255890 3574
rect 266537 3571 266603 3574
rect 351637 3634 351703 3637
rect 358813 3634 358879 3637
rect 351637 3632 358879 3634
rect 351637 3576 351642 3632
rect 351698 3576 358818 3632
rect 358874 3576 358879 3632
rect 351637 3574 358879 3576
rect 351637 3571 351703 3574
rect 358813 3571 358879 3574
rect 274817 3498 274883 3501
rect 252510 3496 274883 3498
rect 252510 3440 274822 3496
rect 274878 3440 274883 3496
rect 252510 3438 274883 3440
rect 249076 3436 249082 3438
rect 252369 3435 252435 3438
rect 274817 3435 274883 3438
rect 285806 3436 285812 3500
rect 285876 3498 285882 3500
rect 286593 3498 286659 3501
rect 285876 3496 286659 3498
rect 285876 3440 286598 3496
rect 286654 3440 286659 3496
rect 285876 3438 286659 3440
rect 285876 3436 285882 3438
rect 286593 3435 286659 3438
rect 287094 3436 287100 3500
rect 287164 3498 287170 3500
rect 287789 3498 287855 3501
rect 287164 3496 287855 3498
rect 287164 3440 287794 3496
rect 287850 3440 287855 3496
rect 287164 3438 287855 3440
rect 287164 3436 287170 3438
rect 287789 3435 287855 3438
rect 288382 3436 288388 3500
rect 288452 3498 288458 3500
rect 288985 3498 289051 3501
rect 288452 3496 289051 3498
rect 288452 3440 288990 3496
rect 289046 3440 289051 3496
rect 288452 3438 289051 3440
rect 288452 3436 288458 3438
rect 288985 3435 289051 3438
rect 291142 3436 291148 3500
rect 291212 3498 291218 3500
rect 291377 3498 291443 3501
rect 291212 3496 291443 3498
rect 291212 3440 291382 3496
rect 291438 3440 291443 3496
rect 291212 3438 291443 3440
rect 291212 3436 291218 3438
rect 291377 3435 291443 3438
rect 299606 3436 299612 3500
rect 299676 3498 299682 3500
rect 300761 3498 300827 3501
rect 299676 3496 300827 3498
rect 299676 3440 300766 3496
rect 300822 3440 300827 3496
rect 299676 3438 300827 3440
rect 299676 3436 299682 3438
rect 300761 3435 300827 3438
rect 304901 3498 304967 3501
rect 305545 3498 305611 3501
rect 304901 3496 305611 3498
rect 304901 3440 304906 3496
rect 304962 3440 305550 3496
rect 305606 3440 305611 3496
rect 304901 3438 305611 3440
rect 304901 3435 304967 3438
rect 305545 3435 305611 3438
rect 348049 3498 348115 3501
rect 357433 3498 357499 3501
rect 348049 3496 357499 3498
rect 348049 3440 348054 3496
rect 348110 3440 357438 3496
rect 357494 3440 357499 3496
rect 348049 3438 357499 3440
rect 348049 3435 348115 3438
rect 357433 3435 357499 3438
rect 15929 3362 15995 3365
rect 200757 3362 200823 3365
rect 15929 3360 200823 3362
rect 15929 3304 15934 3360
rect 15990 3304 200762 3360
rect 200818 3304 200823 3360
rect 15929 3302 200823 3304
rect 15929 3299 15995 3302
rect 200757 3299 200823 3302
rect 213177 3362 213243 3365
rect 276013 3362 276079 3365
rect 213177 3360 276079 3362
rect 213177 3304 213182 3360
rect 213238 3304 276018 3360
rect 276074 3304 276079 3360
rect 213177 3302 276079 3304
rect 213177 3299 213243 3302
rect 276013 3299 276079 3302
rect 344553 3362 344619 3365
rect 356053 3362 356119 3365
rect 344553 3360 356119 3362
rect 344553 3304 344558 3360
rect 344614 3304 356058 3360
rect 356114 3304 356119 3360
rect 344553 3302 356119 3304
rect 344553 3299 344619 3302
rect 356053 3299 356119 3302
rect 186814 2076 186820 2140
rect 186884 2138 186890 2140
rect 239305 2138 239371 2141
rect 186884 2136 239371 2138
rect 186884 2080 239310 2136
rect 239366 2080 239371 2136
rect 186884 2078 239371 2080
rect 186884 2076 186890 2078
rect 239305 2075 239371 2078
rect 82077 2002 82143 2005
rect 195237 2002 195303 2005
rect 82077 2000 195303 2002
rect 82077 1944 82082 2000
rect 82138 1944 195242 2000
rect 195298 1944 195303 2000
rect 82077 1942 195303 1944
rect 82077 1939 82143 1942
rect 195237 1939 195303 1942
<< via3 >>
rect 69612 702476 69676 702540
rect 76052 699484 76116 699548
rect 84332 591908 84396 591972
rect 84332 590820 84396 590884
rect 88196 590684 88260 590748
rect 93900 590004 93964 590068
rect 84332 588704 84396 588708
rect 84332 588648 84382 588704
rect 84382 588648 84396 588704
rect 84332 588644 84396 588648
rect 87828 588704 87892 588708
rect 87828 588648 87878 588704
rect 87878 588648 87892 588704
rect 87828 588644 87892 588648
rect 88932 588432 88996 588436
rect 88932 588376 88946 588432
rect 88946 588376 88996 588432
rect 88932 588372 88996 588376
rect 169708 586468 169772 586532
rect 88196 585516 88260 585580
rect 88932 582932 88996 582996
rect 69428 582252 69492 582316
rect 122604 581572 122668 581636
rect 119476 580212 119540 580276
rect 67772 578308 67836 578372
rect 111012 553420 111076 553484
rect 66668 550836 66732 550900
rect 99972 550700 100036 550764
rect 76052 538052 76116 538116
rect 68140 535468 68204 535532
rect 69612 535528 69676 535532
rect 69612 535472 69662 535528
rect 69662 535472 69676 535528
rect 69612 535468 69676 535472
rect 71820 535468 71884 535532
rect 102180 512620 102244 512684
rect 67772 467740 67836 467804
rect 107700 467060 107764 467124
rect 106412 464340 106476 464404
rect 111748 463524 111812 463588
rect 89668 462844 89732 462908
rect 98132 461484 98196 461548
rect 115980 461484 116044 461548
rect 88196 460124 88260 460188
rect 109172 458220 109236 458284
rect 104940 458084 105004 458148
rect 96660 457404 96724 457468
rect 100708 456044 100772 456108
rect 92796 454684 92860 454748
rect 91140 453188 91204 453252
rect 160140 451284 160204 451348
rect 132540 449924 132604 449988
rect 120028 447884 120092 447948
rect 95188 447748 95252 447812
rect 122972 447748 123036 447812
rect 92612 445708 92676 445772
rect 93900 445708 93964 445772
rect 96476 445708 96540 445772
rect 102364 445708 102428 445772
rect 111564 445708 111628 445772
rect 118556 445708 118620 445772
rect 68876 444756 68940 444820
rect 114324 444756 114388 444820
rect 109540 444680 109604 444684
rect 109540 444624 109554 444680
rect 109554 444624 109604 444680
rect 109540 444620 109604 444624
rect 143580 444620 143644 444684
rect 122604 435780 122668 435844
rect 120028 431428 120092 431492
rect 122604 430884 122668 430948
rect 122972 426260 123036 426324
rect 69244 419324 69308 419388
rect 66668 411300 66732 411364
rect 146892 406268 146956 406332
rect 122972 394708 123036 394772
rect 122788 393212 122852 393276
rect 66116 392532 66180 392596
rect 72372 391172 72436 391236
rect 92796 390960 92860 390964
rect 92796 390904 92846 390960
rect 92846 390904 92860 390960
rect 92796 390900 92860 390904
rect 102180 390960 102244 390964
rect 102180 390904 102194 390960
rect 102194 390904 102244 390960
rect 102180 390900 102244 390904
rect 111012 390900 111076 390964
rect 69612 390356 69676 390420
rect 71820 390416 71884 390420
rect 71820 390360 71870 390416
rect 71870 390360 71884 390416
rect 71820 390356 71884 390360
rect 89668 390356 89732 390420
rect 91140 390356 91204 390420
rect 96660 390356 96724 390420
rect 98132 390356 98196 390420
rect 100708 390416 100772 390420
rect 100708 390360 100722 390416
rect 100722 390360 100772 390416
rect 100708 390356 100772 390360
rect 104940 390356 105004 390420
rect 106412 390356 106476 390420
rect 107700 390356 107764 390420
rect 109172 390356 109236 390420
rect 115980 390416 116044 390420
rect 115980 390360 115994 390416
rect 115994 390360 116044 390416
rect 115980 390356 116044 390360
rect 120028 390356 120092 390420
rect 67772 388996 67836 389060
rect 68140 388996 68204 389060
rect 95188 388996 95252 389060
rect 111748 389056 111812 389060
rect 111748 389000 111798 389056
rect 111798 389000 111812 389056
rect 111748 388996 111812 389000
rect 99972 388860 100036 388924
rect 166948 377300 167012 377364
rect 68876 375940 68940 376004
rect 244228 375396 244292 375460
rect 70164 370500 70228 370564
rect 96476 369608 96540 369612
rect 96476 369552 96490 369608
rect 96490 369552 96540 369608
rect 96476 369548 96540 369552
rect 114324 368324 114388 368388
rect 69796 367644 69860 367708
rect 208900 367100 208964 367164
rect 218652 365740 218716 365804
rect 184060 364380 184124 364444
rect 138060 362204 138124 362268
rect 147444 361796 147508 361860
rect 122604 361660 122668 361724
rect 123340 360224 123404 360228
rect 123340 360168 123354 360224
rect 123354 360168 123404 360224
rect 123340 360164 123404 360168
rect 248460 360164 248524 360228
rect 252508 358804 252572 358868
rect 109540 358668 109604 358732
rect 151860 356628 151924 356692
rect 111564 356084 111628 356148
rect 232452 354860 232516 354924
rect 92612 353288 92676 353292
rect 92612 353232 92662 353288
rect 92662 353232 92676 353288
rect 92612 353228 92676 353232
rect 69612 351052 69676 351116
rect 102364 351052 102428 351116
rect 155172 351052 155236 351116
rect 178540 350644 178604 350708
rect 233740 350508 233804 350572
rect 136036 349692 136100 349756
rect 118556 349148 118620 349212
rect 70164 347788 70228 347852
rect 223620 347788 223684 347852
rect 66668 347652 66732 347716
rect 156460 346972 156524 347036
rect 66668 346700 66732 346764
rect 115060 346564 115124 346628
rect 203012 346624 203076 346628
rect 203012 346568 203062 346624
rect 203062 346568 203076 346624
rect 203012 346564 203076 346568
rect 67772 346292 67836 346356
rect 67956 345748 68020 345812
rect 186820 345204 186884 345268
rect 228220 340988 228284 341052
rect 291148 339492 291212 339556
rect 159220 335684 159284 335748
rect 212580 334324 212644 334388
rect 295932 334052 295996 334116
rect 115060 333236 115124 333300
rect 93900 332420 93964 332484
rect 84700 330244 84764 330308
rect 145420 330244 145484 330308
rect 137140 328612 137204 328676
rect 67404 328340 67468 328404
rect 84700 327524 84764 327588
rect 86724 327524 86788 327588
rect 154252 327660 154316 327724
rect 207980 327660 208044 327724
rect 154988 327388 155052 327452
rect 83964 327176 84028 327180
rect 83964 327120 83978 327176
rect 83978 327120 84028 327176
rect 83964 327116 84028 327120
rect 150388 327116 150452 327180
rect 154436 327116 154500 327180
rect 155172 324396 155236 324460
rect 154252 323580 154316 323644
rect 155172 323444 155236 323508
rect 154988 322220 155052 322284
rect 65932 320240 65996 320244
rect 159220 320724 159284 320788
rect 65932 320184 65982 320240
rect 65982 320184 65996 320240
rect 65932 320180 65996 320184
rect 238524 318276 238588 318340
rect 66668 316372 66732 316436
rect 69428 315828 69492 315892
rect 66116 314196 66180 314260
rect 154436 313924 154500 313988
rect 195100 313244 195164 313308
rect 302740 309164 302804 309228
rect 67404 307940 67468 308004
rect 246252 304132 246316 304196
rect 57836 303724 57900 303788
rect 188292 301004 188356 301068
rect 244044 299644 244108 299708
rect 214052 297468 214116 297532
rect 69428 295428 69492 295492
rect 160140 295292 160204 295356
rect 197860 292572 197924 292636
rect 199332 291484 199396 291548
rect 156460 291076 156524 291140
rect 249748 288628 249812 288692
rect 285628 288492 285692 288556
rect 284340 287540 284404 287604
rect 173020 287132 173084 287196
rect 159220 286316 159284 286380
rect 195468 286316 195532 286380
rect 210740 285772 210804 285836
rect 223620 285636 223684 285700
rect 236500 285636 236564 285700
rect 198780 284548 198844 284612
rect 200620 284548 200684 284612
rect 237420 284548 237484 284612
rect 66116 283732 66180 283796
rect 154252 283460 154316 283524
rect 222700 284004 222764 284068
rect 226932 284004 226996 284068
rect 205404 283928 205468 283932
rect 205404 283872 205418 283928
rect 205418 283872 205468 283928
rect 205404 283868 205468 283872
rect 212396 283868 212460 283932
rect 214420 283928 214484 283932
rect 214420 283872 214470 283928
rect 214470 283872 214484 283928
rect 214420 283868 214484 283872
rect 215892 283928 215956 283932
rect 215892 283872 215942 283928
rect 215942 283872 215956 283928
rect 215892 283868 215956 283872
rect 216628 283868 216692 283932
rect 221228 283928 221292 283932
rect 221228 283872 221278 283928
rect 221278 283872 221292 283928
rect 221228 283868 221292 283872
rect 224724 283928 224788 283932
rect 224724 283872 224738 283928
rect 224738 283872 224788 283928
rect 224724 283868 224788 283872
rect 226196 283868 226260 283932
rect 230244 283868 230308 283932
rect 231716 283868 231780 283932
rect 236500 283868 236564 283932
rect 240364 283868 240428 283932
rect 244412 282372 244476 282436
rect 184060 280740 184124 280804
rect 196572 280740 196636 280804
rect 67956 279380 68020 279444
rect 199332 279380 199396 279444
rect 251220 278896 251284 278900
rect 251220 278840 251270 278896
rect 251270 278840 251284 278896
rect 251220 278836 251284 278840
rect 197860 277204 197924 277268
rect 67956 276116 68020 276180
rect 244228 275572 244292 275636
rect 246252 273260 246316 273324
rect 274588 272172 274652 272236
rect 244228 270540 244292 270604
rect 161980 269316 162044 269380
rect 244044 269044 244108 269108
rect 67404 266868 67468 266932
rect 166212 265508 166276 265572
rect 198780 265508 198844 265572
rect 155356 264148 155420 264212
rect 198780 259388 198844 259452
rect 69428 258708 69492 258772
rect 168972 258028 169036 258092
rect 193812 254356 193876 254420
rect 66668 251908 66732 251972
rect 244044 250548 244108 250612
rect 67772 248916 67836 248980
rect 245700 247284 245764 247348
rect 198780 247012 198844 247076
rect 199884 247012 199948 247076
rect 195468 245924 195532 245988
rect 154436 243884 154500 243948
rect 195284 243748 195348 243812
rect 69428 243340 69492 243404
rect 154804 243204 154868 243268
rect 248460 242932 248524 242996
rect 67404 242796 67468 242860
rect 136036 242040 136100 242044
rect 136036 241984 136050 242040
rect 136050 241984 136100 242040
rect 136036 241980 136100 241984
rect 138060 241980 138124 242044
rect 147444 241980 147508 242044
rect 151860 241980 151924 242044
rect 191604 241632 191668 241636
rect 191604 241576 191654 241632
rect 191654 241576 191668 241632
rect 191604 241572 191668 241576
rect 69612 240756 69676 240820
rect 154436 240348 154500 240412
rect 245884 240212 245948 240276
rect 200252 240076 200316 240140
rect 200436 240076 200500 240140
rect 218652 240076 218716 240140
rect 228220 240076 228284 240140
rect 233740 240076 233804 240140
rect 238524 240076 238588 240140
rect 200252 239668 200316 239732
rect 207980 239396 208044 239460
rect 238892 238776 238956 238780
rect 238892 238720 238942 238776
rect 238942 238720 238956 238776
rect 238892 238716 238956 238720
rect 203012 238580 203076 238644
rect 212580 238580 212644 238644
rect 214052 238580 214116 238644
rect 232452 238580 232516 238644
rect 242020 237492 242084 237556
rect 137140 237280 137204 237284
rect 137140 237224 137154 237280
rect 137154 237224 137204 237280
rect 137140 237220 137204 237224
rect 155356 237220 155420 237284
rect 208900 237220 208964 237284
rect 252508 235860 252572 235924
rect 159220 235724 159284 235788
rect 72372 235588 72436 235652
rect 195284 235588 195348 235652
rect 196572 235588 196636 235652
rect 69796 234228 69860 234292
rect 240364 233956 240428 234020
rect 132540 233004 132604 233068
rect 143580 231100 143644 231164
rect 216628 230420 216692 230484
rect 154068 230284 154132 230348
rect 245700 230284 245764 230348
rect 67956 228924 68020 228988
rect 84700 227564 84764 227628
rect 245884 227564 245948 227628
rect 86724 227428 86788 227492
rect 215892 226400 215956 226404
rect 215892 226344 215942 226400
rect 215942 226344 215956 226400
rect 215892 226340 215956 226344
rect 223620 225932 223684 225996
rect 230244 225116 230308 225180
rect 244228 224768 244292 224772
rect 244228 224712 244278 224768
rect 244278 224712 244292 224768
rect 244228 224708 244292 224712
rect 150388 224164 150452 224228
rect 251220 223076 251284 223140
rect 216628 222804 216692 222868
rect 193812 220764 193876 220828
rect 280292 219404 280356 219468
rect 231900 216744 231964 216748
rect 231900 216688 231914 216744
rect 231914 216688 231964 216744
rect 231900 216684 231964 216688
rect 299612 214508 299676 214572
rect 191604 211108 191668 211172
rect 214420 211168 214484 211172
rect 214420 211112 214470 211168
rect 214470 211112 214484 211168
rect 214420 211108 214484 211112
rect 210740 207844 210804 207908
rect 154620 207572 154684 207636
rect 298140 206212 298204 206276
rect 244044 205124 244108 205188
rect 66668 204852 66732 204916
rect 83964 203492 84028 203556
rect 251772 203492 251836 203556
rect 166212 201316 166276 201380
rect 288388 200772 288452 200836
rect 252508 199548 252572 199612
rect 240364 199412 240428 199476
rect 222700 198188 222764 198252
rect 224724 196692 224788 196756
rect 169524 194380 169588 194444
rect 65932 193972 65996 194036
rect 283788 193972 283852 194036
rect 287100 193836 287164 193900
rect 280476 192612 280540 192676
rect 255820 192476 255884 192540
rect 249012 191116 249076 191180
rect 161980 189620 162044 189684
rect 221228 188532 221292 188596
rect 242940 188396 243004 188460
rect 240732 186356 240796 186420
rect 246252 185676 246316 185740
rect 291332 185676 291396 185740
rect 168972 185540 169036 185604
rect 145420 184180 145484 184244
rect 288572 184180 288636 184244
rect 237604 183092 237668 183156
rect 226932 182956 226996 183020
rect 284524 182956 284588 183020
rect 285812 182820 285876 182884
rect 233188 182004 233252 182068
rect 230612 181460 230676 181524
rect 281580 181460 281644 181524
rect 229876 180644 229940 180708
rect 274588 179012 274652 179076
rect 278820 178604 278884 178668
rect 231716 178332 231780 178396
rect 113220 178196 113284 178260
rect 166212 178060 166276 178124
rect 97028 177924 97092 177988
rect 98316 177516 98380 177580
rect 100708 177576 100772 177580
rect 100708 177520 100758 177576
rect 100758 177520 100772 177576
rect 100708 177516 100772 177520
rect 105676 177516 105740 177580
rect 108068 177516 108132 177580
rect 115796 177576 115860 177580
rect 115796 177520 115846 177576
rect 115846 177520 115860 177576
rect 115796 177516 115860 177520
rect 119476 177576 119540 177580
rect 119476 177520 119526 177576
rect 119526 177520 119540 177576
rect 119476 177516 119540 177520
rect 121868 177516 121932 177580
rect 123156 177516 123220 177580
rect 125732 177516 125796 177580
rect 127020 177516 127084 177580
rect 129412 177516 129476 177580
rect 132356 177576 132420 177580
rect 132356 177520 132406 177576
rect 132406 177520 132420 177576
rect 132356 177516 132420 177520
rect 133092 177576 133156 177580
rect 133092 177520 133142 177576
rect 133142 177520 133156 177576
rect 133092 177516 133156 177520
rect 134380 177516 134444 177580
rect 148180 177576 148244 177580
rect 148180 177520 148230 177576
rect 148230 177520 148244 177576
rect 148180 177516 148244 177520
rect 230428 177380 230492 177444
rect 287284 177380 287348 177444
rect 104572 177244 104636 177308
rect 106964 177108 107028 177172
rect 109540 176972 109604 177036
rect 112116 176972 112180 177036
rect 279372 176972 279436 177036
rect 101996 176836 102060 176900
rect 229140 176896 229204 176900
rect 229140 176840 229190 176896
rect 229190 176840 229204 176896
rect 229140 176836 229204 176840
rect 116900 176760 116964 176764
rect 116900 176704 116950 176760
rect 116950 176704 116964 176760
rect 116900 176700 116964 176704
rect 120764 176700 120828 176764
rect 124444 176760 124508 176764
rect 124444 176704 124494 176760
rect 124494 176704 124508 176760
rect 124444 176700 124508 176704
rect 136036 176760 136100 176764
rect 136036 176704 136086 176760
rect 136086 176704 136100 176760
rect 136036 176700 136100 176704
rect 158852 176700 158916 176764
rect 226196 176564 226260 176628
rect 230612 176564 230676 176628
rect 99420 176428 99484 176492
rect 103284 176428 103348 176492
rect 128124 176428 128188 176492
rect 118372 175884 118436 175948
rect 223620 175944 223684 175948
rect 223620 175888 223670 175944
rect 223670 175888 223684 175944
rect 223620 175884 223684 175888
rect 130700 175672 130764 175676
rect 130700 175616 130750 175672
rect 130750 175616 130764 175672
rect 130700 175612 130764 175616
rect 232084 175884 232148 175948
rect 234660 175748 234724 175812
rect 114324 175476 114388 175540
rect 110644 175340 110708 175404
rect 229876 173844 229940 173908
rect 279372 173708 279436 173772
rect 232084 170852 232148 170916
rect 281580 170852 281644 170916
rect 237420 167996 237484 168060
rect 284524 167860 284588 167924
rect 279372 167588 279436 167652
rect 240364 166908 240428 166972
rect 236500 165140 236564 165204
rect 244228 160652 244292 160716
rect 233740 159020 233804 159084
rect 232636 157932 232700 157996
rect 231900 157388 231964 157452
rect 291332 156028 291396 156092
rect 166212 154532 166276 154596
rect 238892 153716 238956 153780
rect 230980 152356 231044 152420
rect 244780 151812 244844 151876
rect 249748 151812 249812 151876
rect 233004 151132 233068 151196
rect 242020 151132 242084 151196
rect 229140 149636 229204 149700
rect 287284 149092 287348 149156
rect 242020 148004 242084 148068
rect 230428 145284 230492 145348
rect 240732 144604 240796 144668
rect 250484 143924 250548 143988
rect 169524 142700 169588 142764
rect 231164 142700 231228 142764
rect 233004 142428 233068 142492
rect 232636 142020 232700 142084
rect 232452 141068 232516 141132
rect 252508 140116 252572 140180
rect 237972 139708 238036 139772
rect 233188 139164 233252 139228
rect 237604 138756 237668 138820
rect 238156 138348 238220 138412
rect 234660 137804 234724 137868
rect 242940 136308 243004 136372
rect 283788 135084 283852 135148
rect 260052 134540 260116 134604
rect 178540 133044 178604 133108
rect 166212 132772 166276 132836
rect 230980 131548 231044 131612
rect 262812 131004 262876 131068
rect 266860 129236 266924 129300
rect 253060 128692 253124 128756
rect 267780 128420 267844 128484
rect 264100 127876 264164 127940
rect 258580 127060 258644 127124
rect 280108 126788 280172 126852
rect 230980 126516 231044 126580
rect 231164 123524 231228 123588
rect 280292 120668 280356 120732
rect 250300 119172 250364 119236
rect 240732 119036 240796 119100
rect 233740 118356 233804 118420
rect 262076 114548 262140 114612
rect 230244 112100 230308 112164
rect 284340 111556 284404 111620
rect 250484 111012 250548 111076
rect 285628 106932 285692 106996
rect 242020 106116 242084 106180
rect 288572 104892 288636 104956
rect 166396 103804 166460 103868
rect 260052 102716 260116 102780
rect 168972 101356 169036 101420
rect 262996 100404 263060 100468
rect 260052 99724 260116 99788
rect 263180 99180 263244 99244
rect 238156 98772 238220 98836
rect 262996 98772 263060 98836
rect 232452 97956 232516 98020
rect 268516 97548 268580 97612
rect 168420 96596 168484 96660
rect 229140 96596 229204 96660
rect 244780 96460 244844 96524
rect 263180 96324 263244 96388
rect 223620 95976 223684 95980
rect 223620 95920 223670 95976
rect 223670 95920 223684 95976
rect 223620 95916 223684 95920
rect 230244 95236 230308 95300
rect 205404 95100 205468 95164
rect 212396 94964 212460 95028
rect 106478 94828 106542 94892
rect 106780 94828 106844 94892
rect 151308 94828 151372 94892
rect 151766 94828 151830 94892
rect 268516 94828 268580 94892
rect 106228 94692 106292 94756
rect 106614 94692 106678 94756
rect 110150 94752 110214 94756
rect 110150 94696 110198 94752
rect 110198 94696 110214 94752
rect 110150 94692 110214 94696
rect 125382 94752 125446 94756
rect 125382 94696 125414 94752
rect 125414 94696 125446 94752
rect 125382 94692 125446 94696
rect 166212 94420 166276 94484
rect 98500 93876 98564 93940
rect 131988 93740 132052 93804
rect 111932 93604 111996 93668
rect 200620 93604 200684 93668
rect 108068 93528 108132 93532
rect 108068 93472 108118 93528
rect 108118 93472 108132 93528
rect 108068 93468 108132 93472
rect 121684 93528 121748 93532
rect 121684 93472 121734 93528
rect 121734 93472 121748 93528
rect 121684 93468 121748 93472
rect 123156 93468 123220 93532
rect 99972 92440 100036 92444
rect 99972 92384 100022 92440
rect 100022 92384 100036 92440
rect 99972 92380 100036 92384
rect 105676 92440 105740 92444
rect 105676 92384 105726 92440
rect 105726 92384 105740 92440
rect 105676 92380 105740 92384
rect 111196 92380 111260 92444
rect 113220 92380 113284 92444
rect 115428 92440 115492 92444
rect 115428 92384 115478 92440
rect 115478 92384 115492 92440
rect 115428 92380 115492 92384
rect 118004 92440 118068 92444
rect 118004 92384 118054 92440
rect 118054 92384 118068 92440
rect 118004 92380 118068 92384
rect 136036 92440 136100 92444
rect 136036 92384 136086 92440
rect 136086 92384 136100 92440
rect 136036 92380 136100 92384
rect 152044 92440 152108 92444
rect 152044 92384 152094 92440
rect 152094 92384 152108 92440
rect 152044 92380 152108 92384
rect 125732 92244 125796 92308
rect 127572 92108 127636 92172
rect 106228 91972 106292 92036
rect 85804 91700 85868 91764
rect 104204 91700 104268 91764
rect 112300 91700 112364 91764
rect 114876 91700 114940 91764
rect 120580 91700 120644 91764
rect 100892 91564 100956 91628
rect 122788 91428 122852 91492
rect 151492 91488 151556 91492
rect 151492 91432 151542 91488
rect 151542 91432 151556 91488
rect 151492 91428 151556 91432
rect 93900 91292 93964 91356
rect 96660 91292 96724 91356
rect 101996 91352 102060 91356
rect 101996 91296 102010 91352
rect 102010 91296 102060 91352
rect 101996 91292 102060 91296
rect 109172 91292 109236 91356
rect 116716 91292 116780 91356
rect 119660 91352 119724 91356
rect 119660 91296 119710 91352
rect 119710 91296 119724 91352
rect 119660 91292 119724 91296
rect 151308 91292 151372 91356
rect 74764 91156 74828 91220
rect 84332 91156 84396 91220
rect 86724 91216 86788 91220
rect 86724 91160 86774 91216
rect 86774 91160 86788 91216
rect 86724 91156 86788 91160
rect 88012 91156 88076 91220
rect 88932 91156 88996 91220
rect 90220 91156 90284 91220
rect 91324 91156 91388 91220
rect 92612 91156 92676 91220
rect 95004 91216 95068 91220
rect 95004 91160 95054 91216
rect 95054 91160 95068 91216
rect 95004 91156 95068 91160
rect 96292 91156 96356 91220
rect 97212 91156 97276 91220
rect 98132 91156 98196 91220
rect 99052 91156 99116 91220
rect 100524 91216 100588 91220
rect 100524 91160 100574 91216
rect 100574 91160 100588 91216
rect 100524 91156 100588 91160
rect 101812 91156 101876 91220
rect 102732 91156 102796 91220
rect 104572 91156 104636 91220
rect 105492 91216 105556 91220
rect 105492 91160 105542 91216
rect 105542 91160 105556 91216
rect 105492 91156 105556 91160
rect 106780 91156 106844 91220
rect 107700 91156 107764 91220
rect 109540 91156 109604 91220
rect 110644 91156 110708 91220
rect 113220 91156 113284 91220
rect 114324 91216 114388 91220
rect 114324 91160 114338 91216
rect 114338 91160 114388 91216
rect 114324 91156 114388 91160
rect 115796 91156 115860 91220
rect 117084 91156 117148 91220
rect 118188 91156 118252 91220
rect 119292 91156 119356 91220
rect 120212 91156 120276 91220
rect 122052 91156 122116 91220
rect 124076 91216 124140 91220
rect 124076 91160 124126 91216
rect 124126 91160 124140 91216
rect 124076 91156 124140 91160
rect 124444 91156 124508 91220
rect 126468 91216 126532 91220
rect 126468 91160 126518 91216
rect 126518 91160 126532 91216
rect 126468 91156 126532 91160
rect 126652 91156 126716 91220
rect 129412 91156 129476 91220
rect 130700 91156 130764 91220
rect 133092 91156 133156 91220
rect 134380 91156 134444 91220
rect 151676 91216 151740 91220
rect 151676 91160 151690 91216
rect 151690 91160 151740 91216
rect 151676 91156 151740 91160
rect 102548 90884 102612 90948
rect 166396 83948 166460 84012
rect 168972 81364 169036 81428
rect 262812 72524 262876 72588
rect 258580 66812 258644 66876
rect 253060 62732 253124 62796
rect 57836 57156 57900 57220
rect 260052 55796 260116 55860
rect 230980 51716 231044 51780
rect 266860 48860 266924 48924
rect 169708 43420 169772 43484
rect 240732 39340 240796 39404
rect 264100 39204 264164 39268
rect 267780 26828 267844 26892
rect 237972 25468 238036 25532
rect 227668 24108 227732 24172
rect 173020 22748 173084 22812
rect 262076 21252 262140 21316
rect 67772 19892 67836 19956
rect 168420 15812 168484 15876
rect 195100 14452 195164 14516
rect 166948 12956 167012 13020
rect 188292 12956 188356 13020
rect 66116 11596 66180 11660
rect 223620 7652 223684 7716
rect 250300 7516 250364 7580
rect 302740 4796 302804 4860
rect 295932 3980 295996 4044
rect 298140 3844 298204 3908
rect 251772 3572 251836 3636
rect 246252 3436 246316 3500
rect 249012 3436 249076 3500
rect 255820 3572 255884 3636
rect 285812 3436 285876 3500
rect 287100 3436 287164 3500
rect 288388 3436 288452 3500
rect 291148 3436 291212 3500
rect 299612 3436 299676 3500
rect 186820 2076 186884 2140
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 457174 60134 492618
rect 59514 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 60134 457174
rect 59514 456854 60134 456938
rect 59514 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 60134 456854
rect 59514 421174 60134 456618
rect 59514 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 60134 421174
rect 59514 420854 60134 420938
rect 59514 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 60134 420854
rect 59514 385174 60134 420618
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 57835 303788 57901 303789
rect 57835 303724 57836 303788
rect 57900 303724 57901 303788
rect 57835 303723 57901 303724
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 57838 57221 57898 303723
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 205174 60134 240618
rect 59514 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 60134 205174
rect 59514 204854 60134 204938
rect 59514 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 60134 204854
rect 59514 169174 60134 204618
rect 59514 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 60134 169174
rect 59514 168854 60134 168938
rect 59514 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 60134 168854
rect 59514 133174 60134 168618
rect 59514 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 60134 133174
rect 59514 132854 60134 132938
rect 59514 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 60134 132854
rect 59514 97174 60134 132618
rect 59514 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 60134 97174
rect 59514 96854 60134 96938
rect 59514 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 60134 96854
rect 59514 61174 60134 96618
rect 59514 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 60134 61174
rect 59514 60854 60134 60938
rect 59514 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 60134 60854
rect 55794 57134 56414 57218
rect 57835 57220 57901 57221
rect 57835 57156 57836 57220
rect 57900 57156 57901 57220
rect 57835 57155 57901 57156
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 60618
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 69611 702540 69677 702541
rect 69611 702476 69612 702540
rect 69676 702476 69677 702540
rect 69611 702475 69677 702476
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 591166 67574 608058
rect 69614 586530 69674 702475
rect 73794 687454 74414 704282
rect 76051 699548 76117 699549
rect 76051 699484 76052 699548
rect 76116 699484 76117 699548
rect 76051 699483 76117 699484
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 591166 74414 614898
rect 69430 586470 69674 586530
rect 69430 582317 69490 586470
rect 69427 582316 69493 582317
rect 69427 582252 69428 582316
rect 69492 582252 69493 582316
rect 69427 582251 69493 582252
rect 72679 579454 72999 579486
rect 72679 579218 72721 579454
rect 72957 579218 72999 579454
rect 72679 579134 72999 579218
rect 72679 578898 72721 579134
rect 72957 578898 72999 579134
rect 72679 578866 72999 578898
rect 67771 578372 67837 578373
rect 67771 578308 67772 578372
rect 67836 578308 67837 578372
rect 67771 578307 67837 578308
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 66667 550900 66733 550901
rect 66667 550836 66668 550900
rect 66732 550836 66733 550900
rect 66667 550835 66733 550836
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 460894 63854 496338
rect 63234 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 63854 460894
rect 63234 460574 63854 460658
rect 63234 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 63854 460574
rect 63234 424894 63854 460338
rect 63234 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 63854 424894
rect 63234 424574 63854 424658
rect 63234 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 63854 424574
rect 63234 388894 63854 424338
rect 66670 411365 66730 550835
rect 66954 536614 67574 537166
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 464614 67574 500058
rect 67774 467805 67834 578307
rect 75644 561454 75964 561486
rect 75644 561218 75686 561454
rect 75922 561218 75964 561454
rect 75644 561134 75964 561218
rect 75644 560898 75686 561134
rect 75922 560898 75964 561134
rect 75644 560866 75964 560898
rect 72679 543454 72999 543486
rect 72679 543218 72721 543454
rect 72957 543218 72999 543454
rect 72679 543134 72999 543218
rect 72679 542898 72721 543134
rect 72957 542898 72999 543134
rect 72679 542866 72999 542898
rect 76054 538117 76114 699483
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 591166 78134 618618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 591166 81854 622338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84331 591972 84397 591973
rect 84331 591908 84332 591972
rect 84396 591908 84397 591972
rect 84331 591907 84397 591908
rect 84334 590885 84394 591907
rect 84954 591166 85574 626058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 84331 590884 84397 590885
rect 84331 590820 84332 590884
rect 84396 590820 84397 590884
rect 84331 590819 84397 590820
rect 84334 588709 84394 590819
rect 88195 590748 88261 590749
rect 88195 590684 88196 590748
rect 88260 590684 88261 590748
rect 88195 590683 88261 590684
rect 84331 588708 84397 588709
rect 84331 588644 84332 588708
rect 84396 588644 84397 588708
rect 84331 588643 84397 588644
rect 87827 588708 87893 588709
rect 87827 588644 87828 588708
rect 87892 588644 87893 588708
rect 87827 588643 87893 588644
rect 87830 582390 87890 588643
rect 88198 585581 88258 590683
rect 88931 588436 88997 588437
rect 88931 588372 88932 588436
rect 88996 588372 88997 588436
rect 88931 588371 88997 588372
rect 88195 585580 88261 585581
rect 88195 585516 88196 585580
rect 88260 585516 88261 585580
rect 88195 585515 88261 585516
rect 88934 582997 88994 588371
rect 88931 582996 88997 582997
rect 88931 582932 88932 582996
rect 88996 582932 88997 582996
rect 88931 582931 88997 582932
rect 87830 582330 88258 582390
rect 78609 579454 78929 579486
rect 78609 579218 78651 579454
rect 78887 579218 78929 579454
rect 78609 579134 78929 579218
rect 78609 578898 78651 579134
rect 78887 578898 78929 579134
rect 78609 578866 78929 578898
rect 84540 579454 84860 579486
rect 84540 579218 84582 579454
rect 84818 579218 84860 579454
rect 84540 579134 84860 579218
rect 84540 578898 84582 579134
rect 84818 578898 84860 579134
rect 84540 578866 84860 578898
rect 81575 561454 81895 561486
rect 81575 561218 81617 561454
rect 81853 561218 81895 561454
rect 81575 561134 81895 561218
rect 81575 560898 81617 561134
rect 81853 560898 81895 561134
rect 81575 560866 81895 560898
rect 78609 543454 78929 543486
rect 78609 543218 78651 543454
rect 78887 543218 78929 543454
rect 78609 543134 78929 543218
rect 78609 542898 78651 543134
rect 78887 542898 78929 543134
rect 78609 542866 78929 542898
rect 84540 543454 84860 543486
rect 84540 543218 84582 543454
rect 84818 543218 84860 543454
rect 84540 543134 84860 543218
rect 84540 542898 84582 543134
rect 84818 542898 84860 543134
rect 84540 542866 84860 542898
rect 76051 538116 76117 538117
rect 76051 538052 76052 538116
rect 76116 538052 76117 538116
rect 76051 538051 76117 538052
rect 68139 535532 68205 535533
rect 68139 535468 68140 535532
rect 68204 535468 68205 535532
rect 68139 535467 68205 535468
rect 69611 535532 69677 535533
rect 69611 535468 69612 535532
rect 69676 535468 69677 535532
rect 69611 535467 69677 535468
rect 71819 535532 71885 535533
rect 71819 535468 71820 535532
rect 71884 535468 71885 535532
rect 71819 535467 71885 535468
rect 67771 467804 67837 467805
rect 67771 467740 67772 467804
rect 67836 467740 67837 467804
rect 67771 467739 67837 467740
rect 66954 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 67574 464614
rect 66954 464294 67574 464378
rect 66954 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 67574 464294
rect 66954 446407 67574 464058
rect 66667 411364 66733 411365
rect 66667 411300 66668 411364
rect 66732 411300 66733 411364
rect 66667 411299 66733 411300
rect 66115 392596 66181 392597
rect 66115 392532 66116 392596
rect 66180 392532 66181 392596
rect 66115 392531 66181 392532
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 65931 320244 65997 320245
rect 65931 320180 65932 320244
rect 65996 320180 65997 320244
rect 65931 320179 65997 320180
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 208894 63854 244338
rect 63234 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 63854 208894
rect 63234 208574 63854 208658
rect 63234 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 63854 208574
rect 63234 172894 63854 208338
rect 65934 194037 65994 320179
rect 66118 314261 66178 392531
rect 68142 389061 68202 535467
rect 68875 444820 68941 444821
rect 68875 444756 68876 444820
rect 68940 444756 68941 444820
rect 68875 444755 68941 444756
rect 67771 389060 67837 389061
rect 67771 388996 67772 389060
rect 67836 388996 67837 389060
rect 67771 388995 67837 388996
rect 68139 389060 68205 389061
rect 68139 388996 68140 389060
rect 68204 388996 68205 389060
rect 68139 388995 68205 388996
rect 66954 356614 67574 388356
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66667 347716 66733 347717
rect 66667 347652 66668 347716
rect 66732 347652 66733 347716
rect 66667 347651 66733 347652
rect 66670 346765 66730 347651
rect 66667 346764 66733 346765
rect 66667 346700 66668 346764
rect 66732 346700 66733 346764
rect 66667 346699 66733 346700
rect 66670 316437 66730 346699
rect 66954 329592 67574 356058
rect 67774 346357 67834 388995
rect 68878 376005 68938 444755
rect 69614 425070 69674 535467
rect 69062 425010 69674 425070
rect 69062 417890 69122 425010
rect 69243 419388 69309 419389
rect 69243 419324 69244 419388
rect 69308 419386 69309 419388
rect 69308 419326 69858 419386
rect 69308 419324 69309 419326
rect 69243 419323 69309 419324
rect 69062 417830 69674 417890
rect 69614 390421 69674 417830
rect 69611 390420 69677 390421
rect 69611 390356 69612 390420
rect 69676 390356 69677 390420
rect 69611 390355 69677 390356
rect 68875 376004 68941 376005
rect 68875 375940 68876 376004
rect 68940 375940 68941 376004
rect 68875 375939 68941 375940
rect 69798 367709 69858 419326
rect 71822 390421 71882 535467
rect 73794 507454 74414 537166
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 471454 74414 506898
rect 73794 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 74414 471454
rect 73794 471134 74414 471218
rect 73794 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 74414 471134
rect 73794 446407 74414 470898
rect 77514 511174 78134 537166
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 475174 78134 510618
rect 77514 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 78134 475174
rect 77514 474854 78134 474938
rect 77514 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 78134 474854
rect 77514 446407 78134 474618
rect 81234 514894 81854 537166
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 478894 81854 514338
rect 81234 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 81854 478894
rect 81234 478574 81854 478658
rect 81234 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 81854 478574
rect 81234 446407 81854 478338
rect 84954 518614 85574 537166
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 482614 85574 518058
rect 84954 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 85574 482614
rect 84954 482294 85574 482378
rect 84954 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 85574 482294
rect 84954 446407 85574 482058
rect 88198 460189 88258 582330
rect 91794 561454 92414 596898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 93899 590068 93965 590069
rect 93899 590004 93900 590068
rect 93964 590004 93965 590068
rect 93899 590003 93965 590004
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 89667 462908 89733 462909
rect 89667 462844 89668 462908
rect 89732 462844 89733 462908
rect 89667 462843 89733 462844
rect 88195 460188 88261 460189
rect 88195 460124 88196 460188
rect 88260 460124 88261 460188
rect 88195 460123 88261 460124
rect 72978 435454 73298 435486
rect 72978 435218 73020 435454
rect 73256 435218 73298 435454
rect 72978 435134 73298 435218
rect 72978 434898 73020 435134
rect 73256 434898 73298 435134
rect 72978 434866 73298 434898
rect 88338 417454 88658 417486
rect 88338 417218 88380 417454
rect 88616 417218 88658 417454
rect 88338 417134 88658 417218
rect 88338 416898 88380 417134
rect 88616 416898 88658 417134
rect 88338 416866 88658 416898
rect 72978 399454 73298 399486
rect 72978 399218 73020 399454
rect 73256 399218 73298 399454
rect 72978 399134 73298 399218
rect 72978 398898 73020 399134
rect 73256 398898 73298 399134
rect 72978 398866 73298 398898
rect 72371 391236 72437 391237
rect 72371 391172 72372 391236
rect 72436 391172 72437 391236
rect 72371 391171 72437 391172
rect 71819 390420 71885 390421
rect 71819 390356 71820 390420
rect 71884 390356 71885 390420
rect 71819 390355 71885 390356
rect 70163 370564 70229 370565
rect 70163 370500 70164 370564
rect 70228 370500 70229 370564
rect 70163 370499 70229 370500
rect 69795 367708 69861 367709
rect 69795 367644 69796 367708
rect 69860 367644 69861 367708
rect 69795 367643 69861 367644
rect 69611 351116 69677 351117
rect 69611 351052 69612 351116
rect 69676 351052 69677 351116
rect 69611 351051 69677 351052
rect 67771 346356 67837 346357
rect 67771 346292 67772 346356
rect 67836 346292 67837 346356
rect 67771 346291 67837 346292
rect 67955 345812 68021 345813
rect 67955 345748 67956 345812
rect 68020 345748 68021 345812
rect 67955 345747 68021 345748
rect 67403 328404 67469 328405
rect 67403 328340 67404 328404
rect 67468 328340 67469 328404
rect 67403 328339 67469 328340
rect 66667 316436 66733 316437
rect 66667 316372 66668 316436
rect 66732 316372 66733 316436
rect 66667 316371 66733 316372
rect 66115 314260 66181 314261
rect 66115 314196 66116 314260
rect 66180 314196 66181 314260
rect 66115 314195 66181 314196
rect 67406 308005 67466 328339
rect 67403 308004 67469 308005
rect 67403 307940 67404 308004
rect 67468 307940 67469 308004
rect 67403 307939 67469 307940
rect 66115 283796 66181 283797
rect 66115 283732 66116 283796
rect 66180 283732 66181 283796
rect 66115 283731 66181 283732
rect 65931 194036 65997 194037
rect 65931 193972 65932 194036
rect 65996 193972 65997 194036
rect 65931 193971 65997 193972
rect 63234 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 63854 172894
rect 63234 172574 63854 172658
rect 63234 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 63854 172574
rect 63234 136894 63854 172338
rect 63234 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 63854 136894
rect 63234 136574 63854 136658
rect 63234 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 63854 136574
rect 63234 100894 63854 136338
rect 63234 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 63854 100894
rect 63234 100574 63854 100658
rect 63234 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 63854 100574
rect 63234 64894 63854 100338
rect 63234 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 63854 64894
rect 63234 64574 63854 64658
rect 63234 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 63854 64574
rect 63234 28894 63854 64338
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 66118 11661 66178 283731
rect 67958 279445 68018 345747
rect 69614 321570 69674 351051
rect 70166 347853 70226 370499
rect 70163 347852 70229 347853
rect 70163 347788 70164 347852
rect 70228 347788 70229 347852
rect 70163 347787 70229 347788
rect 70166 335370 70226 347787
rect 69246 321510 69674 321570
rect 69798 335310 70226 335370
rect 69246 311910 69306 321510
rect 69798 317250 69858 335310
rect 69430 317190 69858 317250
rect 69430 315893 69490 317190
rect 69427 315892 69493 315893
rect 69427 315828 69428 315892
rect 69492 315828 69493 315892
rect 69427 315827 69493 315828
rect 69246 311850 69674 311910
rect 69614 296730 69674 311850
rect 69430 296670 69674 296730
rect 69430 295493 69490 296670
rect 69427 295492 69493 295493
rect 69427 295428 69428 295492
rect 69492 295428 69493 295492
rect 69427 295427 69493 295428
rect 67955 279444 68021 279445
rect 67955 279380 67956 279444
rect 68020 279380 68021 279444
rect 67955 279379 68021 279380
rect 67955 276180 68021 276181
rect 67955 276116 67956 276180
rect 68020 276116 68021 276180
rect 67955 276115 68021 276116
rect 67403 266932 67469 266933
rect 67403 266868 67404 266932
rect 67468 266868 67469 266932
rect 67403 266867 67469 266868
rect 66667 251972 66733 251973
rect 66667 251908 66668 251972
rect 66732 251908 66733 251972
rect 66667 251907 66733 251908
rect 66670 204917 66730 251907
rect 67406 242861 67466 266867
rect 67771 248980 67837 248981
rect 67771 248916 67772 248980
rect 67836 248916 67837 248980
rect 67771 248915 67837 248916
rect 67403 242860 67469 242861
rect 67403 242796 67404 242860
rect 67468 242796 67469 242860
rect 67403 242795 67469 242796
rect 66954 212614 67574 239592
rect 66954 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 67574 212614
rect 66954 212294 67574 212378
rect 66954 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 67574 212294
rect 66667 204916 66733 204917
rect 66667 204852 66668 204916
rect 66732 204852 66733 204916
rect 66667 204851 66733 204852
rect 66954 176600 67574 212058
rect 66954 68614 67574 93100
rect 66954 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 67574 68614
rect 66954 68294 67574 68378
rect 66954 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 67574 68294
rect 66954 32614 67574 68058
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 66115 11660 66181 11661
rect 66115 11596 66116 11660
rect 66180 11596 66181 11660
rect 66115 11595 66181 11596
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 67774 19957 67834 248915
rect 67958 228989 68018 276115
rect 69427 258772 69493 258773
rect 69427 258708 69428 258772
rect 69492 258708 69493 258772
rect 69427 258707 69493 258708
rect 69430 258090 69490 258707
rect 69430 258030 69674 258090
rect 69427 243404 69493 243405
rect 69427 243340 69428 243404
rect 69492 243340 69493 243404
rect 69427 243339 69493 243340
rect 69430 238770 69490 243339
rect 69614 240821 69674 258030
rect 69611 240820 69677 240821
rect 69611 240756 69612 240820
rect 69676 240756 69677 240820
rect 69611 240755 69677 240756
rect 69430 238710 69858 238770
rect 69798 234293 69858 238710
rect 72374 235653 72434 391171
rect 89670 390421 89730 462843
rect 91794 453454 92414 488898
rect 92795 454748 92861 454749
rect 92795 454684 92796 454748
rect 92860 454684 92861 454748
rect 92795 454683 92861 454684
rect 91139 453252 91205 453253
rect 91139 453188 91140 453252
rect 91204 453188 91205 453252
rect 91139 453187 91205 453188
rect 91794 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 92414 453454
rect 91142 390421 91202 453187
rect 91794 453134 92414 453218
rect 91794 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 92414 453134
rect 91794 446407 92414 452898
rect 92611 445772 92677 445773
rect 92611 445708 92612 445772
rect 92676 445708 92677 445772
rect 92611 445707 92677 445708
rect 89667 390420 89733 390421
rect 89667 390356 89668 390420
rect 89732 390356 89733 390420
rect 89667 390355 89733 390356
rect 91139 390420 91205 390421
rect 91139 390356 91140 390420
rect 91204 390356 91205 390420
rect 91139 390355 91205 390356
rect 73794 363454 74414 388356
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 329592 74414 362898
rect 77514 367174 78134 388356
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 329592 78134 330618
rect 81234 370894 81854 388356
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 329592 81854 334338
rect 84954 374614 85574 388356
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84699 330308 84765 330309
rect 84699 330244 84700 330308
rect 84764 330244 84765 330308
rect 84699 330243 84765 330244
rect 84702 327589 84762 330243
rect 84954 329592 85574 338058
rect 91794 381454 92414 388356
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 92614 353293 92674 445707
rect 92798 390965 92858 454683
rect 93902 445773 93962 590003
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 95514 457174 96134 492618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 99971 550764 100037 550765
rect 99971 550700 99972 550764
rect 100036 550700 100037 550764
rect 99971 550699 100037 550700
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 98131 461548 98197 461549
rect 98131 461484 98132 461548
rect 98196 461484 98197 461548
rect 98131 461483 98197 461484
rect 96659 457468 96725 457469
rect 96659 457404 96660 457468
rect 96724 457404 96725 457468
rect 96659 457403 96725 457404
rect 95514 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 96134 457174
rect 95514 456854 96134 456938
rect 95514 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 96134 456854
rect 95187 447812 95253 447813
rect 95187 447748 95188 447812
rect 95252 447748 95253 447812
rect 95187 447747 95253 447748
rect 93899 445772 93965 445773
rect 93899 445708 93900 445772
rect 93964 445708 93965 445772
rect 93899 445707 93965 445708
rect 92795 390964 92861 390965
rect 92795 390900 92796 390964
rect 92860 390900 92861 390964
rect 92795 390899 92861 390900
rect 92611 353292 92677 353293
rect 92611 353228 92612 353292
rect 92676 353228 92677 353292
rect 92611 353227 92677 353228
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 329592 92414 344898
rect 93902 332485 93962 445707
rect 95190 389061 95250 447747
rect 95514 446407 96134 456618
rect 96475 445772 96541 445773
rect 96475 445708 96476 445772
rect 96540 445708 96541 445772
rect 96475 445707 96541 445708
rect 95187 389060 95253 389061
rect 95187 388996 95188 389060
rect 95252 388996 95253 389060
rect 95187 388995 95253 388996
rect 95514 385174 96134 388356
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 96478 369613 96538 445707
rect 96662 390421 96722 457403
rect 98134 390421 98194 461483
rect 99234 460894 99854 496338
rect 99234 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 99854 460894
rect 99234 460574 99854 460658
rect 99234 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 99854 460574
rect 99234 446407 99854 460338
rect 96659 390420 96725 390421
rect 96659 390356 96660 390420
rect 96724 390356 96725 390420
rect 96659 390355 96725 390356
rect 98131 390420 98197 390421
rect 98131 390356 98132 390420
rect 98196 390356 98197 390420
rect 98131 390355 98197 390356
rect 99974 388925 100034 550699
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102179 512684 102245 512685
rect 102179 512620 102180 512684
rect 102244 512620 102245 512684
rect 102179 512619 102245 512620
rect 100707 456108 100773 456109
rect 100707 456044 100708 456108
rect 100772 456044 100773 456108
rect 100707 456043 100773 456044
rect 100710 390421 100770 456043
rect 102182 390965 102242 512619
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 102954 464614 103574 500058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 111011 553484 111077 553485
rect 111011 553420 111012 553484
rect 111076 553420 111077 553484
rect 111011 553419 111077 553420
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 471454 110414 506898
rect 109794 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 110414 471454
rect 109794 471134 110414 471218
rect 109794 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 110414 471134
rect 107699 467124 107765 467125
rect 107699 467060 107700 467124
rect 107764 467060 107765 467124
rect 107699 467059 107765 467060
rect 102954 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 103574 464614
rect 102954 464294 103574 464378
rect 106411 464404 106477 464405
rect 106411 464340 106412 464404
rect 106476 464340 106477 464404
rect 106411 464339 106477 464340
rect 102954 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 103574 464294
rect 102954 446407 103574 464058
rect 104939 458148 105005 458149
rect 104939 458084 104940 458148
rect 105004 458084 105005 458148
rect 104939 458083 105005 458084
rect 102363 445772 102429 445773
rect 102363 445708 102364 445772
rect 102428 445708 102429 445772
rect 102363 445707 102429 445708
rect 102179 390964 102245 390965
rect 102179 390900 102180 390964
rect 102244 390900 102245 390964
rect 102179 390899 102245 390900
rect 100707 390420 100773 390421
rect 100707 390356 100708 390420
rect 100772 390356 100773 390420
rect 100707 390355 100773 390356
rect 99971 388924 100037 388925
rect 99971 388860 99972 388924
rect 100036 388860 100037 388924
rect 99971 388859 100037 388860
rect 96475 369612 96541 369613
rect 96475 369548 96476 369612
rect 96540 369548 96541 369612
rect 96475 369547 96541 369548
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 93899 332484 93965 332485
rect 93899 332420 93900 332484
rect 93964 332420 93965 332484
rect 93899 332419 93965 332420
rect 95514 329592 96134 348618
rect 99234 352894 99854 388356
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 329592 99854 352338
rect 102366 351117 102426 445707
rect 103698 435454 104018 435486
rect 103698 435218 103740 435454
rect 103976 435218 104018 435454
rect 103698 435134 104018 435218
rect 103698 434898 103740 435134
rect 103976 434898 104018 435134
rect 103698 434866 104018 434898
rect 103698 399454 104018 399486
rect 103698 399218 103740 399454
rect 103976 399218 104018 399454
rect 103698 399134 104018 399218
rect 103698 398898 103740 399134
rect 103976 398898 104018 399134
rect 103698 398866 104018 398898
rect 104942 390421 105002 458083
rect 106414 390421 106474 464339
rect 107702 390421 107762 467059
rect 109171 458284 109237 458285
rect 109171 458220 109172 458284
rect 109236 458220 109237 458284
rect 109171 458219 109237 458220
rect 109174 390421 109234 458219
rect 109794 446407 110414 470898
rect 109539 444684 109605 444685
rect 109539 444620 109540 444684
rect 109604 444620 109605 444684
rect 109539 444619 109605 444620
rect 104939 390420 105005 390421
rect 104939 390356 104940 390420
rect 105004 390356 105005 390420
rect 104939 390355 105005 390356
rect 106411 390420 106477 390421
rect 106411 390356 106412 390420
rect 106476 390356 106477 390420
rect 106411 390355 106477 390356
rect 107699 390420 107765 390421
rect 107699 390356 107700 390420
rect 107764 390356 107765 390420
rect 107699 390355 107765 390356
rect 109171 390420 109237 390421
rect 109171 390356 109172 390420
rect 109236 390356 109237 390420
rect 109171 390355 109237 390356
rect 102954 356614 103574 388356
rect 109542 358733 109602 444619
rect 111014 390965 111074 553419
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 113514 475174 114134 510618
rect 113514 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 114134 475174
rect 113514 474854 114134 474938
rect 113514 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 114134 474854
rect 111747 463588 111813 463589
rect 111747 463524 111748 463588
rect 111812 463524 111813 463588
rect 111747 463523 111813 463524
rect 111563 445772 111629 445773
rect 111563 445708 111564 445772
rect 111628 445708 111629 445772
rect 111563 445707 111629 445708
rect 111011 390964 111077 390965
rect 111011 390900 111012 390964
rect 111076 390900 111077 390964
rect 111011 390899 111077 390900
rect 109794 363454 110414 388356
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109539 358732 109605 358733
rect 109539 358668 109540 358732
rect 109604 358668 109605 358732
rect 109539 358667 109605 358668
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102363 351116 102429 351117
rect 102363 351052 102364 351116
rect 102428 351052 102429 351116
rect 102363 351051 102429 351052
rect 102954 329592 103574 356058
rect 109794 329592 110414 362898
rect 111566 356149 111626 445707
rect 111750 389061 111810 463523
rect 113514 446407 114134 474618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 119475 580276 119541 580277
rect 119475 580212 119476 580276
rect 119540 580212 119541 580276
rect 119475 580211 119541 580212
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 478894 117854 514338
rect 117234 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 117854 478894
rect 117234 478574 117854 478658
rect 117234 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 117854 478574
rect 115979 461548 116045 461549
rect 115979 461484 115980 461548
rect 116044 461484 116045 461548
rect 115979 461483 116045 461484
rect 114323 444820 114389 444821
rect 114323 444756 114324 444820
rect 114388 444756 114389 444820
rect 114323 444755 114389 444756
rect 111747 389060 111813 389061
rect 111747 388996 111748 389060
rect 111812 388996 111813 389060
rect 111747 388995 111813 388996
rect 113514 367174 114134 388356
rect 114326 368389 114386 444755
rect 115982 390421 116042 461483
rect 117234 446407 117854 478338
rect 118555 445772 118621 445773
rect 118555 445708 118556 445772
rect 118620 445708 118621 445772
rect 118555 445707 118621 445708
rect 115979 390420 116045 390421
rect 115979 390356 115980 390420
rect 116044 390356 116045 390420
rect 115979 390355 116045 390356
rect 117234 370894 117854 388356
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 114323 368388 114389 368389
rect 114323 368324 114324 368388
rect 114388 368324 114389 368388
rect 114323 368323 114389 368324
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 111563 356148 111629 356149
rect 111563 356084 111564 356148
rect 111628 356084 111629 356148
rect 111563 356083 111629 356084
rect 113514 331174 114134 366618
rect 115059 346628 115125 346629
rect 115059 346564 115060 346628
rect 115124 346564 115125 346628
rect 115059 346563 115125 346564
rect 115062 333301 115122 346563
rect 117234 334894 117854 370338
rect 118558 349213 118618 445707
rect 119478 441630 119538 580211
rect 120954 554614 121574 590058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 122603 581636 122669 581637
rect 122603 581572 122604 581636
rect 122668 581572 122669 581636
rect 122603 581571 122669 581572
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 120954 482614 121574 518058
rect 120954 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 121574 482614
rect 120954 482294 121574 482378
rect 120954 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 121574 482294
rect 120027 447948 120093 447949
rect 120027 447884 120028 447948
rect 120092 447884 120093 447948
rect 120027 447883 120093 447884
rect 120030 441630 120090 447883
rect 120954 446407 121574 482058
rect 119478 441570 119906 441630
rect 120030 441570 120458 441630
rect 119846 431490 119906 441570
rect 120027 431492 120093 431493
rect 120027 431490 120028 431492
rect 119846 431430 120028 431490
rect 120027 431428 120028 431430
rect 120092 431428 120093 431492
rect 120027 431427 120093 431428
rect 119058 417454 119378 417486
rect 119058 417218 119100 417454
rect 119336 417218 119378 417454
rect 119058 417134 119378 417218
rect 119058 416898 119100 417134
rect 119336 416898 119378 417134
rect 119058 416866 119378 416898
rect 120398 412650 120458 441570
rect 122606 435845 122666 581571
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 127794 453454 128414 488898
rect 127794 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 128414 453454
rect 127794 453134 128414 453218
rect 127794 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 128414 453134
rect 122971 447812 123037 447813
rect 122971 447748 122972 447812
rect 123036 447748 123037 447812
rect 122971 447747 123037 447748
rect 122603 435844 122669 435845
rect 122603 435780 122604 435844
rect 122668 435780 122669 435844
rect 122603 435779 122669 435780
rect 122603 430948 122669 430949
rect 122603 430884 122604 430948
rect 122668 430884 122669 430948
rect 122603 430883 122669 430884
rect 120030 412590 120458 412650
rect 120030 390421 120090 412590
rect 120027 390420 120093 390421
rect 120027 390356 120028 390420
rect 120092 390356 120093 390420
rect 120027 390355 120093 390356
rect 120954 374614 121574 388356
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 118555 349212 118621 349213
rect 118555 349148 118556 349212
rect 118620 349148 118621 349212
rect 118555 349147 118621 349148
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 115059 333300 115125 333301
rect 115059 333236 115060 333300
rect 115124 333236 115125 333300
rect 115059 333235 115125 333236
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 329592 114134 330618
rect 117234 329592 117854 334338
rect 120954 338614 121574 374058
rect 122606 361725 122666 430883
rect 122974 426325 123034 447747
rect 122971 426324 123037 426325
rect 122971 426260 122972 426324
rect 123036 426260 123037 426324
rect 122971 426259 123037 426260
rect 122974 422310 123034 426259
rect 122974 422250 123402 422310
rect 122971 394772 123037 394773
rect 122971 394708 122972 394772
rect 123036 394708 123037 394772
rect 122971 394707 123037 394708
rect 122974 393330 123034 394707
rect 122790 393277 123034 393330
rect 122787 393276 123034 393277
rect 122787 393212 122788 393276
rect 122852 393270 123034 393276
rect 122852 393212 122853 393270
rect 122787 393211 122853 393212
rect 122603 361724 122669 361725
rect 122603 361660 122604 361724
rect 122668 361660 122669 361724
rect 122603 361659 122669 361660
rect 123342 360229 123402 422250
rect 127794 417454 128414 452898
rect 127794 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 128414 417454
rect 127794 417134 128414 417218
rect 127794 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 128414 417134
rect 127794 381454 128414 416898
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 123339 360228 123405 360229
rect 123339 360164 123340 360228
rect 123404 360164 123405 360228
rect 123339 360163 123405 360164
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 329592 121574 338058
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 329592 128414 344898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 131514 457174 132134 492618
rect 131514 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 132134 457174
rect 131514 456854 132134 456938
rect 131514 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 132134 456854
rect 131514 421174 132134 456618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 460894 135854 496338
rect 135234 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 135854 460894
rect 135234 460574 135854 460658
rect 135234 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 135854 460574
rect 132539 449988 132605 449989
rect 132539 449924 132540 449988
rect 132604 449924 132605 449988
rect 132539 449923 132605 449924
rect 131514 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 132134 421174
rect 131514 420854 132134 420938
rect 131514 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 132134 420854
rect 131514 385174 132134 420618
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 329592 132134 348618
rect 84699 327588 84765 327589
rect 84699 327524 84700 327588
rect 84764 327524 84765 327588
rect 84699 327523 84765 327524
rect 86723 327588 86789 327589
rect 86723 327524 86724 327588
rect 86788 327524 86789 327588
rect 86723 327523 86789 327524
rect 83963 327180 84029 327181
rect 83963 327116 83964 327180
rect 84028 327116 84029 327180
rect 83963 327115 84029 327116
rect 72978 291454 73298 291486
rect 72978 291218 73020 291454
rect 73256 291218 73298 291454
rect 72978 291134 73298 291218
rect 72978 290898 73020 291134
rect 73256 290898 73298 291134
rect 72978 290866 73298 290898
rect 72978 255454 73298 255486
rect 72978 255218 73020 255454
rect 73256 255218 73298 255454
rect 72978 255134 73298 255218
rect 72978 254898 73020 255134
rect 73256 254898 73298 255134
rect 72978 254866 73298 254898
rect 72371 235652 72437 235653
rect 72371 235588 72372 235652
rect 72436 235588 72437 235652
rect 72371 235587 72437 235588
rect 69795 234292 69861 234293
rect 69795 234228 69796 234292
rect 69860 234228 69861 234292
rect 69795 234227 69861 234228
rect 67955 228988 68021 228989
rect 67955 228924 67956 228988
rect 68020 228924 68021 228988
rect 67955 228923 68021 228924
rect 73794 219454 74414 239592
rect 73794 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 74414 219454
rect 73794 219134 74414 219218
rect 73794 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 74414 219134
rect 73794 183454 74414 218898
rect 73794 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 74414 183454
rect 73794 183134 74414 183218
rect 73794 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 74414 183134
rect 73794 176600 74414 182898
rect 77514 223174 78134 239592
rect 77514 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 78134 223174
rect 77514 222854 78134 222938
rect 77514 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 78134 222854
rect 77514 187174 78134 222618
rect 77514 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 78134 187174
rect 77514 186854 78134 186938
rect 77514 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 78134 186854
rect 77514 176600 78134 186618
rect 81234 226894 81854 239592
rect 81234 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 81854 226894
rect 81234 226574 81854 226658
rect 81234 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 81854 226574
rect 81234 190894 81854 226338
rect 83966 203557 84026 327115
rect 84702 227629 84762 327523
rect 84954 230614 85574 239592
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84699 227628 84765 227629
rect 84699 227564 84700 227628
rect 84764 227564 84765 227628
rect 84699 227563 84765 227564
rect 83963 203556 84029 203557
rect 83963 203492 83964 203556
rect 84028 203492 84029 203556
rect 83963 203491 84029 203492
rect 81234 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 81854 190894
rect 81234 190574 81854 190658
rect 81234 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 81854 190574
rect 81234 176600 81854 190338
rect 84954 194614 85574 230058
rect 86726 227493 86786 327523
rect 88338 309454 88658 309486
rect 88338 309218 88380 309454
rect 88616 309218 88658 309454
rect 88338 309134 88658 309218
rect 88338 308898 88380 309134
rect 88616 308898 88658 309134
rect 88338 308866 88658 308898
rect 119058 309454 119378 309486
rect 119058 309218 119100 309454
rect 119336 309218 119378 309454
rect 119058 309134 119378 309218
rect 119058 308898 119100 309134
rect 119336 308898 119378 309134
rect 119058 308866 119378 308898
rect 103698 291454 104018 291486
rect 103698 291218 103740 291454
rect 103976 291218 104018 291454
rect 103698 291134 104018 291218
rect 103698 290898 103740 291134
rect 103976 290898 104018 291134
rect 103698 290866 104018 290898
rect 88338 273454 88658 273486
rect 88338 273218 88380 273454
rect 88616 273218 88658 273454
rect 88338 273134 88658 273218
rect 88338 272898 88380 273134
rect 88616 272898 88658 273134
rect 88338 272866 88658 272898
rect 119058 273454 119378 273486
rect 119058 273218 119100 273454
rect 119336 273218 119378 273454
rect 119058 273134 119378 273218
rect 119058 272898 119100 273134
rect 119336 272898 119378 273134
rect 119058 272866 119378 272898
rect 103698 255454 104018 255486
rect 103698 255218 103740 255454
rect 103976 255218 104018 255454
rect 103698 255134 104018 255218
rect 103698 254898 103740 255134
rect 103976 254898 104018 255134
rect 103698 254866 104018 254898
rect 91794 237454 92414 239592
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 86723 227492 86789 227493
rect 86723 227428 86724 227492
rect 86788 227428 86789 227492
rect 86723 227427 86789 227428
rect 84954 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 85574 194614
rect 84954 194294 85574 194378
rect 84954 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 85574 194294
rect 84954 176600 85574 194058
rect 91794 201454 92414 236898
rect 91794 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 92414 201454
rect 91794 201134 92414 201218
rect 91794 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 92414 201134
rect 91794 176600 92414 200898
rect 95514 205174 96134 239592
rect 95514 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 96134 205174
rect 95514 204854 96134 204938
rect 95514 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 96134 204854
rect 95514 176600 96134 204618
rect 99234 208894 99854 239592
rect 99234 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 99854 208894
rect 99234 208574 99854 208658
rect 99234 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 99854 208574
rect 97027 177988 97093 177989
rect 97027 177924 97028 177988
rect 97092 177924 97093 177988
rect 97027 177923 97093 177924
rect 97030 175130 97090 177923
rect 98315 177580 98381 177581
rect 98315 177516 98316 177580
rect 98380 177516 98381 177580
rect 98315 177515 98381 177516
rect 96960 175070 97090 175130
rect 98318 175130 98378 177515
rect 99234 176600 99854 208338
rect 102954 212614 103574 239592
rect 102954 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 103574 212614
rect 102954 212294 103574 212378
rect 102954 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 103574 212294
rect 100707 177580 100773 177581
rect 100707 177516 100708 177580
rect 100772 177516 100773 177580
rect 100707 177515 100773 177516
rect 99419 176492 99485 176493
rect 99419 176428 99420 176492
rect 99484 176428 99485 176492
rect 99419 176427 99485 176428
rect 99422 175130 99482 176427
rect 98318 175070 98380 175130
rect 96960 174494 97020 175070
rect 98320 174494 98380 175070
rect 99408 175070 99482 175130
rect 100710 175130 100770 177515
rect 101995 176900 102061 176901
rect 101995 176836 101996 176900
rect 102060 176836 102061 176900
rect 101995 176835 102061 176836
rect 101998 175130 102058 176835
rect 102954 176600 103574 212058
rect 109794 219454 110414 239592
rect 109794 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 110414 219454
rect 109794 219134 110414 219218
rect 109794 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 110414 219134
rect 109794 183454 110414 218898
rect 109794 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 110414 183454
rect 109794 183134 110414 183218
rect 109794 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 110414 183134
rect 105675 177580 105741 177581
rect 105675 177516 105676 177580
rect 105740 177516 105741 177580
rect 105675 177515 105741 177516
rect 108067 177580 108133 177581
rect 108067 177516 108068 177580
rect 108132 177516 108133 177580
rect 108067 177515 108133 177516
rect 104571 177308 104637 177309
rect 104571 177244 104572 177308
rect 104636 177244 104637 177308
rect 104571 177243 104637 177244
rect 103283 176492 103349 176493
rect 103283 176428 103284 176492
rect 103348 176428 103349 176492
rect 103283 176427 103349 176428
rect 100710 175070 100828 175130
rect 99408 174494 99468 175070
rect 100768 174494 100828 175070
rect 101992 175070 102058 175130
rect 103286 175130 103346 176427
rect 104574 175130 104634 177243
rect 105678 175130 105738 177515
rect 106963 177172 107029 177173
rect 106963 177108 106964 177172
rect 107028 177108 107029 177172
rect 106963 177107 107029 177108
rect 103286 175070 103412 175130
rect 104574 175070 104636 175130
rect 101992 174494 102052 175070
rect 103352 174494 103412 175070
rect 104576 174494 104636 175070
rect 105664 175070 105738 175130
rect 106966 175130 107026 177107
rect 108070 175130 108130 177515
rect 109539 177036 109605 177037
rect 109539 176972 109540 177036
rect 109604 176972 109605 177036
rect 109539 176971 109605 176972
rect 109542 175130 109602 176971
rect 109794 176600 110414 182898
rect 113514 223174 114134 239592
rect 113514 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 114134 223174
rect 113514 222854 114134 222938
rect 113514 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 114134 222854
rect 113514 187174 114134 222618
rect 113514 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 114134 187174
rect 113514 186854 114134 186938
rect 113514 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 114134 186854
rect 113219 178260 113285 178261
rect 113219 178196 113220 178260
rect 113284 178196 113285 178260
rect 113219 178195 113285 178196
rect 112115 177036 112181 177037
rect 112115 176972 112116 177036
rect 112180 176972 112181 177036
rect 112115 176971 112181 176972
rect 110643 175404 110709 175405
rect 110643 175340 110644 175404
rect 110708 175340 110709 175404
rect 110643 175339 110709 175340
rect 106966 175070 107084 175130
rect 108070 175070 108172 175130
rect 105664 174494 105724 175070
rect 107024 174494 107084 175070
rect 108112 174494 108172 175070
rect 109472 175070 109602 175130
rect 110646 175130 110706 175339
rect 112118 175130 112178 176971
rect 113222 175130 113282 178195
rect 113514 176600 114134 186618
rect 117234 226894 117854 239592
rect 117234 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 117854 226894
rect 117234 226574 117854 226658
rect 117234 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 117854 226574
rect 117234 190894 117854 226338
rect 117234 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 117854 190894
rect 117234 190574 117854 190658
rect 117234 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 117854 190574
rect 115795 177580 115861 177581
rect 115795 177516 115796 177580
rect 115860 177516 115861 177580
rect 115795 177515 115861 177516
rect 114323 175540 114389 175541
rect 114323 175476 114324 175540
rect 114388 175476 114389 175540
rect 114323 175475 114389 175476
rect 110646 175070 110756 175130
rect 109472 174494 109532 175070
rect 110696 174494 110756 175070
rect 112056 175070 112178 175130
rect 113144 175070 113282 175130
rect 114326 175130 114386 175475
rect 115798 175130 115858 177515
rect 116899 176764 116965 176765
rect 116899 176700 116900 176764
rect 116964 176700 116965 176764
rect 116899 176699 116965 176700
rect 114326 175070 114428 175130
rect 112056 174494 112116 175070
rect 113144 174494 113204 175070
rect 114368 174494 114428 175070
rect 115728 175070 115858 175130
rect 116902 175130 116962 176699
rect 117234 176600 117854 190338
rect 120954 230614 121574 239592
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 194614 121574 230058
rect 120954 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 121574 194614
rect 120954 194294 121574 194378
rect 120954 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 121574 194294
rect 119475 177580 119541 177581
rect 119475 177516 119476 177580
rect 119540 177516 119541 177580
rect 119475 177515 119541 177516
rect 118371 175948 118437 175949
rect 118371 175884 118372 175948
rect 118436 175884 118437 175948
rect 118371 175883 118437 175884
rect 118374 175130 118434 175883
rect 119478 175130 119538 177515
rect 120763 176764 120829 176765
rect 120763 176700 120764 176764
rect 120828 176700 120829 176764
rect 120763 176699 120829 176700
rect 120766 175130 120826 176699
rect 120954 176600 121574 194058
rect 127794 237454 128414 239592
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 201454 128414 236898
rect 127794 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 128414 201454
rect 127794 201134 128414 201218
rect 127794 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 128414 201134
rect 121867 177580 121933 177581
rect 121867 177516 121868 177580
rect 121932 177516 121933 177580
rect 121867 177515 121933 177516
rect 123155 177580 123221 177581
rect 123155 177516 123156 177580
rect 123220 177516 123221 177580
rect 123155 177515 123221 177516
rect 125731 177580 125797 177581
rect 125731 177516 125732 177580
rect 125796 177516 125797 177580
rect 125731 177515 125797 177516
rect 127019 177580 127085 177581
rect 127019 177516 127020 177580
rect 127084 177516 127085 177580
rect 127019 177515 127085 177516
rect 121870 175130 121930 177515
rect 123158 175130 123218 177515
rect 124443 176764 124509 176765
rect 124443 176700 124444 176764
rect 124508 176700 124509 176764
rect 124443 176699 124509 176700
rect 124446 175130 124506 176699
rect 125734 175130 125794 177515
rect 127022 175130 127082 177515
rect 127794 176600 128414 200898
rect 131514 205174 132134 239592
rect 132542 233069 132602 449923
rect 135234 424894 135854 460338
rect 135234 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 135854 424894
rect 135234 424574 135854 424658
rect 135234 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 135854 424574
rect 135234 388894 135854 424338
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138954 464614 139574 500058
rect 138954 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 139574 464614
rect 138954 464294 139574 464378
rect 138954 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 139574 464294
rect 138954 428614 139574 464058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145794 471454 146414 506898
rect 145794 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 146414 471454
rect 145794 471134 146414 471218
rect 145794 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 146414 471134
rect 143579 444684 143645 444685
rect 143579 444620 143580 444684
rect 143644 444620 143645 444684
rect 143579 444619 143645 444620
rect 138954 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 139574 428614
rect 138954 428294 139574 428378
rect 138954 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 139574 428294
rect 138954 392614 139574 428058
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138059 362268 138125 362269
rect 138059 362204 138060 362268
rect 138124 362204 138125 362268
rect 138059 362203 138125 362204
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 329592 135854 352338
rect 136035 349756 136101 349757
rect 136035 349692 136036 349756
rect 136100 349692 136101 349756
rect 136035 349691 136101 349692
rect 134418 291454 134738 291486
rect 134418 291218 134460 291454
rect 134696 291218 134738 291454
rect 134418 291134 134738 291218
rect 134418 290898 134460 291134
rect 134696 290898 134738 291134
rect 134418 290866 134738 290898
rect 134418 255454 134738 255486
rect 134418 255218 134460 255454
rect 134696 255218 134738 255454
rect 134418 255134 134738 255218
rect 134418 254898 134460 255134
rect 134696 254898 134738 255134
rect 134418 254866 134738 254898
rect 136038 242045 136098 349691
rect 137139 328676 137205 328677
rect 137139 328612 137140 328676
rect 137204 328612 137205 328676
rect 137139 328611 137205 328612
rect 136035 242044 136101 242045
rect 136035 241980 136036 242044
rect 136100 241980 136101 242044
rect 136035 241979 136101 241980
rect 132539 233068 132605 233069
rect 132539 233004 132540 233068
rect 132604 233004 132605 233068
rect 132539 233003 132605 233004
rect 131514 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 132134 205174
rect 131514 204854 132134 204938
rect 131514 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 132134 204854
rect 129411 177580 129477 177581
rect 129411 177516 129412 177580
rect 129476 177516 129477 177580
rect 129411 177515 129477 177516
rect 128123 176492 128189 176493
rect 128123 176428 128124 176492
rect 128188 176428 128189 176492
rect 128123 176427 128189 176428
rect 128126 175130 128186 176427
rect 116902 175070 117012 175130
rect 115728 174494 115788 175070
rect 116952 174494 117012 175070
rect 118312 175070 118434 175130
rect 119400 175070 119538 175130
rect 120760 175070 120826 175130
rect 121848 175070 121930 175130
rect 123072 175070 123218 175130
rect 124432 175070 124506 175130
rect 125656 175070 125794 175130
rect 127016 175070 127082 175130
rect 128104 175070 128186 175130
rect 129414 175130 129474 177515
rect 131514 176600 132134 204618
rect 135234 208894 135854 239592
rect 137142 237285 137202 328611
rect 138062 242045 138122 362203
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 329592 139574 356058
rect 138059 242044 138125 242045
rect 138059 241980 138060 242044
rect 138124 241980 138125 242044
rect 138059 241979 138125 241980
rect 137139 237284 137205 237285
rect 137139 237220 137140 237284
rect 137204 237220 137205 237284
rect 137139 237219 137205 237220
rect 135234 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 135854 208894
rect 135234 208574 135854 208658
rect 135234 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 135854 208574
rect 132355 177580 132421 177581
rect 132355 177516 132356 177580
rect 132420 177516 132421 177580
rect 132355 177515 132421 177516
rect 133091 177580 133157 177581
rect 133091 177516 133092 177580
rect 133156 177516 133157 177580
rect 133091 177515 133157 177516
rect 134379 177580 134445 177581
rect 134379 177516 134380 177580
rect 134444 177516 134445 177580
rect 134379 177515 134445 177516
rect 130699 175676 130765 175677
rect 130699 175612 130700 175676
rect 130764 175612 130765 175676
rect 130699 175611 130765 175612
rect 130702 175130 130762 175611
rect 132358 175130 132418 177515
rect 129414 175070 129524 175130
rect 118312 174494 118372 175070
rect 119400 174494 119460 175070
rect 120760 174494 120820 175070
rect 121848 174494 121908 175070
rect 123072 174494 123132 175070
rect 124432 174494 124492 175070
rect 125656 174494 125716 175070
rect 127016 174494 127076 175070
rect 128104 174494 128164 175070
rect 129464 174494 129524 175070
rect 130688 175070 130762 175130
rect 132048 175070 132418 175130
rect 133094 175130 133154 177515
rect 134382 175130 134442 177515
rect 135234 176600 135854 208338
rect 138954 212614 139574 239592
rect 143582 231165 143642 444619
rect 145794 435454 146414 470898
rect 145794 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 146414 435454
rect 145794 435134 146414 435218
rect 145794 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 146414 435134
rect 145794 399454 146414 434898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 475174 150134 510618
rect 149514 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 150134 475174
rect 149514 474854 150134 474938
rect 149514 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 150134 474854
rect 149514 439174 150134 474618
rect 149514 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 150134 439174
rect 149514 438854 150134 438938
rect 149514 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 150134 438854
rect 146891 406332 146957 406333
rect 146891 406268 146892 406332
rect 146956 406268 146957 406332
rect 146891 406267 146957 406268
rect 145794 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 146414 399454
rect 145794 399134 146414 399218
rect 145794 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 146414 399134
rect 145794 363454 146414 398898
rect 146894 364350 146954 406267
rect 149514 403174 150134 438618
rect 149514 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 150134 403174
rect 149514 402854 150134 402938
rect 149514 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 150134 402854
rect 149514 367174 150134 402618
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 146894 364290 147506 364350
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145419 330308 145485 330309
rect 145419 330244 145420 330308
rect 145484 330244 145485 330308
rect 145419 330243 145485 330244
rect 143579 231164 143645 231165
rect 143579 231100 143580 231164
rect 143644 231100 143645 231164
rect 143579 231099 143645 231100
rect 138954 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 139574 212614
rect 138954 212294 139574 212378
rect 138954 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 139574 212294
rect 136035 176764 136101 176765
rect 136035 176700 136036 176764
rect 136100 176700 136101 176764
rect 136035 176699 136101 176700
rect 136038 175130 136098 176699
rect 138954 176600 139574 212058
rect 145422 184245 145482 330243
rect 145794 329592 146414 362898
rect 147446 361861 147506 364290
rect 147443 361860 147509 361861
rect 147443 361796 147444 361860
rect 147508 361796 147509 361860
rect 147443 361795 147509 361796
rect 147446 242045 147506 361795
rect 149514 331174 150134 366618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 153234 478894 153854 514338
rect 153234 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 153854 478894
rect 153234 478574 153854 478658
rect 153234 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 153854 478574
rect 153234 442894 153854 478338
rect 153234 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 153854 442894
rect 153234 442574 153854 442658
rect 153234 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 153854 442574
rect 153234 406894 153854 442338
rect 153234 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 153854 406894
rect 153234 406574 153854 406658
rect 153234 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 153854 406574
rect 153234 370894 153854 406338
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 151859 356692 151925 356693
rect 151859 356628 151860 356692
rect 151924 356628 151925 356692
rect 151859 356627 151925 356628
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 329592 150134 330618
rect 150387 327180 150453 327181
rect 150387 327116 150388 327180
rect 150452 327116 150453 327180
rect 150387 327115 150453 327116
rect 149778 309454 150098 309486
rect 149778 309218 149820 309454
rect 150056 309218 150098 309454
rect 149778 309134 150098 309218
rect 149778 308898 149820 309134
rect 150056 308898 150098 309134
rect 149778 308866 150098 308898
rect 149778 273454 150098 273486
rect 149778 273218 149820 273454
rect 150056 273218 150098 273454
rect 149778 273134 150098 273218
rect 149778 272898 149820 273134
rect 150056 272898 150098 273134
rect 149778 272866 150098 272898
rect 147443 242044 147509 242045
rect 147443 241980 147444 242044
rect 147508 241980 147509 242044
rect 147443 241979 147509 241980
rect 145794 219454 146414 239592
rect 145794 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 146414 219454
rect 145794 219134 146414 219218
rect 145794 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 146414 219134
rect 145419 184244 145485 184245
rect 145419 184180 145420 184244
rect 145484 184180 145485 184244
rect 145419 184179 145485 184180
rect 145794 183454 146414 218898
rect 145794 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 146414 183454
rect 145794 183134 146414 183218
rect 145794 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 146414 183134
rect 145794 176600 146414 182898
rect 149514 223174 150134 239592
rect 150390 224229 150450 327115
rect 151862 242045 151922 356627
rect 153234 334894 153854 370338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 482614 157574 518058
rect 156954 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 157574 482614
rect 156954 482294 157574 482378
rect 156954 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 157574 482294
rect 156954 446614 157574 482058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 163794 453454 164414 488898
rect 163794 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 164414 453454
rect 163794 453134 164414 453218
rect 163794 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 164414 453134
rect 160139 451348 160205 451349
rect 160139 451284 160140 451348
rect 160204 451284 160205 451348
rect 160139 451283 160205 451284
rect 156954 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 157574 446614
rect 156954 446294 157574 446378
rect 156954 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 157574 446294
rect 156954 410614 157574 446058
rect 156954 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 157574 410614
rect 156954 410294 157574 410378
rect 156954 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 157574 410294
rect 156954 374614 157574 410058
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 155171 351116 155237 351117
rect 155171 351052 155172 351116
rect 155236 351052 155237 351116
rect 155171 351051 155237 351052
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 329592 153854 334338
rect 154251 327724 154317 327725
rect 154251 327660 154252 327724
rect 154316 327660 154317 327724
rect 154251 327659 154317 327660
rect 154254 323645 154314 327659
rect 154987 327452 155053 327453
rect 154987 327388 154988 327452
rect 155052 327388 155053 327452
rect 154987 327387 155053 327388
rect 154435 327180 154501 327181
rect 154435 327116 154436 327180
rect 154500 327116 154501 327180
rect 154435 327115 154501 327116
rect 154251 323644 154317 323645
rect 154251 323580 154252 323644
rect 154316 323580 154317 323644
rect 154251 323579 154317 323580
rect 154438 313989 154498 327115
rect 154990 322285 155050 327387
rect 155174 324461 155234 351051
rect 156459 347036 156525 347037
rect 156459 346972 156460 347036
rect 156524 346972 156525 347036
rect 156459 346971 156525 346972
rect 155171 324460 155237 324461
rect 155171 324396 155172 324460
rect 155236 324396 155237 324460
rect 155171 324395 155237 324396
rect 155174 323509 155234 324395
rect 155171 323508 155237 323509
rect 155171 323444 155172 323508
rect 155236 323444 155237 323508
rect 155171 323443 155237 323444
rect 154987 322284 155053 322285
rect 154987 322220 154988 322284
rect 155052 322220 155053 322284
rect 154987 322219 155053 322220
rect 154435 313988 154501 313989
rect 154435 313924 154436 313988
rect 154500 313924 154501 313988
rect 154435 313923 154501 313924
rect 156462 291141 156522 346971
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 159219 335748 159285 335749
rect 159219 335684 159220 335748
rect 159284 335684 159285 335748
rect 159219 335683 159285 335684
rect 159222 320789 159282 335683
rect 159219 320788 159285 320789
rect 159219 320724 159220 320788
rect 159284 320724 159285 320788
rect 159219 320723 159285 320724
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156459 291140 156525 291141
rect 156459 291076 156460 291140
rect 156524 291076 156525 291140
rect 156459 291075 156525 291076
rect 154251 283524 154317 283525
rect 154251 283460 154252 283524
rect 154316 283460 154317 283524
rect 154251 283459 154317 283460
rect 154254 277410 154314 283459
rect 154070 277350 154314 277410
rect 151859 242044 151925 242045
rect 151859 241980 151860 242044
rect 151924 241980 151925 242044
rect 151859 241979 151925 241980
rect 153234 226894 153854 239592
rect 154070 230349 154130 277350
rect 156954 266614 157574 302058
rect 160142 295357 160202 451283
rect 163794 417454 164414 452898
rect 163794 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 164414 417454
rect 163794 417134 164414 417218
rect 163794 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 164414 417134
rect 163794 381454 164414 416898
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 169707 586532 169773 586533
rect 169707 586468 169708 586532
rect 169772 586468 169773 586532
rect 169707 586467 169773 586468
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 457174 168134 492618
rect 167514 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 168134 457174
rect 167514 456854 168134 456938
rect 167514 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 168134 456854
rect 167514 421174 168134 456618
rect 167514 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 168134 421174
rect 167514 420854 168134 420938
rect 167514 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 168134 420854
rect 167514 385174 168134 420618
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 166947 377364 167013 377365
rect 166947 377300 166948 377364
rect 167012 377300 167013 377364
rect 166947 377299 167013 377300
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 160139 295356 160205 295357
rect 160139 295292 160140 295356
rect 160204 295292 160205 295356
rect 160139 295291 160205 295292
rect 159219 286380 159285 286381
rect 159219 286316 159220 286380
rect 159284 286316 159285 286380
rect 159219 286315 159285 286316
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 155355 264212 155421 264213
rect 155355 264148 155356 264212
rect 155420 264148 155421 264212
rect 155355 264147 155421 264148
rect 154435 243948 154501 243949
rect 154435 243884 154436 243948
rect 154500 243884 154501 243948
rect 154435 243883 154501 243884
rect 154438 240413 154498 243883
rect 154803 243268 154869 243269
rect 154803 243204 154804 243268
rect 154868 243204 154869 243268
rect 154803 243203 154869 243204
rect 154435 240412 154501 240413
rect 154435 240348 154436 240412
rect 154500 240348 154501 240412
rect 154435 240347 154501 240348
rect 154806 238770 154866 243203
rect 154622 238710 154866 238770
rect 154067 230348 154133 230349
rect 154067 230284 154068 230348
rect 154132 230284 154133 230348
rect 154067 230283 154133 230284
rect 153234 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 153854 226894
rect 153234 226574 153854 226658
rect 153234 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 153854 226574
rect 150387 224228 150453 224229
rect 150387 224164 150388 224228
rect 150452 224164 150453 224228
rect 150387 224163 150453 224164
rect 149514 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 150134 223174
rect 149514 222854 150134 222938
rect 149514 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 150134 222854
rect 149514 187174 150134 222618
rect 149514 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 150134 187174
rect 149514 186854 150134 186938
rect 149514 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 150134 186854
rect 148179 177580 148245 177581
rect 148179 177516 148180 177580
rect 148244 177516 148245 177580
rect 148179 177515 148245 177516
rect 133094 175070 133196 175130
rect 130688 174494 130748 175070
rect 132048 174494 132108 175070
rect 133136 174494 133196 175070
rect 134360 175070 134442 175130
rect 135720 175070 136098 175130
rect 148182 175130 148242 177515
rect 149514 176600 150134 186618
rect 153234 190894 153854 226338
rect 154622 207637 154682 238710
rect 155358 237285 155418 264147
rect 155355 237284 155421 237285
rect 155355 237220 155356 237284
rect 155420 237220 155421 237284
rect 155355 237219 155421 237220
rect 156954 230614 157574 266058
rect 159222 235789 159282 286315
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 161979 269380 162045 269381
rect 161979 269316 161980 269380
rect 162044 269316 162045 269380
rect 161979 269315 162045 269316
rect 159219 235788 159285 235789
rect 159219 235724 159220 235788
rect 159284 235724 159285 235788
rect 159219 235723 159285 235724
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 154619 207636 154685 207637
rect 154619 207572 154620 207636
rect 154684 207572 154685 207636
rect 154619 207571 154685 207572
rect 153234 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 153854 190894
rect 153234 190574 153854 190658
rect 153234 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 153854 190574
rect 153234 176600 153854 190338
rect 156954 194614 157574 230058
rect 156954 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 157574 194614
rect 156954 194294 157574 194378
rect 156954 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 157574 194294
rect 156954 176600 157574 194058
rect 161982 189685 162042 269315
rect 163794 237454 164414 272898
rect 166211 265572 166277 265573
rect 166211 265508 166212 265572
rect 166276 265508 166277 265572
rect 166211 265507 166277 265508
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 201454 164414 236898
rect 163794 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 164414 201454
rect 166214 201381 166274 265507
rect 166211 201380 166277 201381
rect 166211 201316 166212 201380
rect 166276 201316 166277 201380
rect 166211 201315 166277 201316
rect 163794 201134 164414 201218
rect 163794 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 164414 201134
rect 161979 189684 162045 189685
rect 161979 189620 161980 189684
rect 162044 189620 162045 189684
rect 161979 189619 162045 189620
rect 158851 176764 158917 176765
rect 158851 176700 158852 176764
rect 158916 176700 158917 176764
rect 158851 176699 158917 176700
rect 158854 175130 158914 176699
rect 163794 176600 164414 200898
rect 166211 178124 166277 178125
rect 166211 178060 166212 178124
rect 166276 178060 166277 178124
rect 166211 178059 166277 178060
rect 148182 175070 148292 175130
rect 134360 174494 134420 175070
rect 135720 174494 135780 175070
rect 148232 174494 148292 175070
rect 158840 175070 158914 175130
rect 158840 174494 158900 175070
rect 69072 165454 69420 165486
rect 69072 165218 69128 165454
rect 69364 165218 69420 165454
rect 69072 165134 69420 165218
rect 69072 164898 69128 165134
rect 69364 164898 69420 165134
rect 69072 164866 69420 164898
rect 164136 165454 164484 165486
rect 164136 165218 164192 165454
rect 164428 165218 164484 165454
rect 164136 165134 164484 165218
rect 164136 164898 164192 165134
rect 164428 164898 164484 165134
rect 164136 164866 164484 164898
rect 166214 154597 166274 178059
rect 166211 154596 166277 154597
rect 166211 154532 166212 154596
rect 166276 154532 166277 154596
rect 166211 154531 166277 154532
rect 69752 147454 70100 147486
rect 69752 147218 69808 147454
rect 70044 147218 70100 147454
rect 69752 147134 70100 147218
rect 69752 146898 69808 147134
rect 70044 146898 70100 147134
rect 69752 146866 70100 146898
rect 163456 147454 163804 147486
rect 163456 147218 163512 147454
rect 163748 147218 163804 147454
rect 163456 147134 163804 147218
rect 163456 146898 163512 147134
rect 163748 146898 163804 147134
rect 163456 146866 163804 146898
rect 166211 132836 166277 132837
rect 166211 132772 166212 132836
rect 166276 132772 166277 132836
rect 166211 132771 166277 132772
rect 69072 129454 69420 129486
rect 69072 129218 69128 129454
rect 69364 129218 69420 129454
rect 69072 129134 69420 129218
rect 69072 128898 69128 129134
rect 69364 128898 69420 129134
rect 69072 128866 69420 128898
rect 164136 129454 164484 129486
rect 164136 129218 164192 129454
rect 164428 129218 164484 129454
rect 164136 129134 164484 129218
rect 164136 128898 164192 129134
rect 164428 128898 164484 129134
rect 164136 128866 164484 128898
rect 69752 111454 70100 111486
rect 69752 111218 69808 111454
rect 70044 111218 70100 111454
rect 69752 111134 70100 111218
rect 69752 110898 69808 111134
rect 70044 110898 70100 111134
rect 69752 110866 70100 110898
rect 163456 111454 163804 111486
rect 163456 111218 163512 111454
rect 163748 111218 163804 111454
rect 163456 111134 163804 111218
rect 163456 110898 163512 111134
rect 163748 110898 163804 111134
rect 163456 110866 163804 110898
rect 74656 94890 74716 95200
rect 84312 94890 84372 95200
rect 85536 94890 85596 95200
rect 86624 94890 86684 95200
rect 87984 94890 88044 95200
rect 88936 94890 88996 95200
rect 74656 94830 74826 94890
rect 84312 94830 84394 94890
rect 85536 94830 85866 94890
rect 86624 94830 86786 94890
rect 87984 94830 88074 94890
rect 73794 75454 74414 93100
rect 74766 91221 74826 94830
rect 74763 91220 74829 91221
rect 74763 91156 74764 91220
rect 74828 91156 74829 91220
rect 74763 91155 74829 91156
rect 73794 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 74414 75454
rect 73794 75134 74414 75218
rect 73794 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 74414 75134
rect 73794 39454 74414 74898
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 67771 19956 67837 19957
rect 67771 19892 67772 19956
rect 67836 19892 67837 19956
rect 67771 19891 67837 19892
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 79174 78134 93100
rect 77514 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 78134 79174
rect 77514 78854 78134 78938
rect 77514 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 78134 78854
rect 77514 43174 78134 78618
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 82894 81854 93100
rect 84334 91221 84394 94830
rect 84331 91220 84397 91221
rect 84331 91156 84332 91220
rect 84396 91156 84397 91220
rect 84331 91155 84397 91156
rect 81234 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 81854 82894
rect 81234 82574 81854 82658
rect 81234 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 81854 82574
rect 81234 46894 81854 82338
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 86614 85574 93100
rect 85806 91765 85866 94830
rect 85803 91764 85869 91765
rect 85803 91700 85804 91764
rect 85868 91700 85869 91764
rect 85803 91699 85869 91700
rect 86726 91221 86786 94830
rect 88014 91221 88074 94830
rect 88934 94830 88996 94890
rect 90160 94890 90220 95200
rect 91384 94890 91444 95200
rect 90160 94830 90282 94890
rect 88934 91221 88994 94830
rect 90222 91221 90282 94830
rect 91326 94830 91444 94890
rect 92472 94890 92532 95200
rect 93832 94890 93892 95200
rect 94920 94890 94980 95200
rect 96008 94890 96068 95200
rect 96688 94890 96748 95200
rect 92472 94830 92674 94890
rect 93832 94830 93962 94890
rect 94920 94830 95066 94890
rect 96008 94830 96354 94890
rect 91326 91221 91386 94830
rect 86723 91220 86789 91221
rect 86723 91156 86724 91220
rect 86788 91156 86789 91220
rect 86723 91155 86789 91156
rect 88011 91220 88077 91221
rect 88011 91156 88012 91220
rect 88076 91156 88077 91220
rect 88011 91155 88077 91156
rect 88931 91220 88997 91221
rect 88931 91156 88932 91220
rect 88996 91156 88997 91220
rect 88931 91155 88997 91156
rect 90219 91220 90285 91221
rect 90219 91156 90220 91220
rect 90284 91156 90285 91220
rect 90219 91155 90285 91156
rect 91323 91220 91389 91221
rect 91323 91156 91324 91220
rect 91388 91156 91389 91220
rect 91323 91155 91389 91156
rect 84954 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 85574 86614
rect 84954 86294 85574 86378
rect 84954 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 85574 86294
rect 84954 50614 85574 86058
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 93100
rect 92614 91221 92674 94830
rect 93902 91357 93962 94830
rect 93899 91356 93965 91357
rect 93899 91292 93900 91356
rect 93964 91292 93965 91356
rect 93899 91291 93965 91292
rect 95006 91221 95066 94830
rect 92611 91220 92677 91221
rect 92611 91156 92612 91220
rect 92676 91156 92677 91220
rect 92611 91155 92677 91156
rect 95003 91220 95069 91221
rect 95003 91156 95004 91220
rect 95068 91156 95069 91220
rect 95003 91155 95069 91156
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 61174 96134 93100
rect 96294 91221 96354 94830
rect 96662 94830 96748 94890
rect 97096 94890 97156 95200
rect 98048 94890 98108 95200
rect 98456 94890 98516 95200
rect 99136 94890 99196 95200
rect 97096 94830 97274 94890
rect 98048 94830 98194 94890
rect 98456 94830 98562 94890
rect 96662 91357 96722 94830
rect 96659 91356 96725 91357
rect 96659 91292 96660 91356
rect 96724 91292 96725 91356
rect 96659 91291 96725 91292
rect 97214 91221 97274 94830
rect 98134 91221 98194 94830
rect 98502 93941 98562 94830
rect 99054 94830 99196 94890
rect 99544 94890 99604 95200
rect 100632 94890 100692 95200
rect 99544 94830 100034 94890
rect 98499 93940 98565 93941
rect 98499 93876 98500 93940
rect 98564 93876 98565 93940
rect 98499 93875 98565 93876
rect 99054 91221 99114 94830
rect 96291 91220 96357 91221
rect 96291 91156 96292 91220
rect 96356 91156 96357 91220
rect 96291 91155 96357 91156
rect 97211 91220 97277 91221
rect 97211 91156 97212 91220
rect 97276 91156 97277 91220
rect 97211 91155 97277 91156
rect 98131 91220 98197 91221
rect 98131 91156 98132 91220
rect 98196 91156 98197 91220
rect 98131 91155 98197 91156
rect 99051 91220 99117 91221
rect 99051 91156 99052 91220
rect 99116 91156 99117 91220
rect 99051 91155 99117 91156
rect 95514 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 96134 61174
rect 95514 60854 96134 60938
rect 95514 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 96134 60854
rect 95514 25174 96134 60618
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 64894 99854 93100
rect 99974 92445 100034 94830
rect 100526 94830 100692 94890
rect 100768 94890 100828 95200
rect 101856 94890 101916 95200
rect 100768 94830 100954 94890
rect 99971 92444 100037 92445
rect 99971 92380 99972 92444
rect 100036 92380 100037 92444
rect 99971 92379 100037 92380
rect 100526 91221 100586 94830
rect 100894 91629 100954 94830
rect 101814 94830 101916 94890
rect 101992 94890 102052 95200
rect 102944 94890 103004 95200
rect 103216 94890 103276 95200
rect 104304 94890 104364 95200
rect 101992 94830 102058 94890
rect 100891 91628 100957 91629
rect 100891 91564 100892 91628
rect 100956 91564 100957 91628
rect 100891 91563 100957 91564
rect 101814 91221 101874 94830
rect 101998 91357 102058 94830
rect 102550 94830 103004 94890
rect 103102 94830 103276 94890
rect 104206 94830 104364 94890
rect 104440 94890 104500 95200
rect 105392 94890 105452 95200
rect 105664 94890 105724 95200
rect 106480 94893 106540 95200
rect 106477 94892 106543 94893
rect 104440 94830 104634 94890
rect 105392 94830 105554 94890
rect 105664 94830 105738 94890
rect 101995 91356 102061 91357
rect 101995 91292 101996 91356
rect 102060 91292 102061 91356
rect 101995 91291 102061 91292
rect 100523 91220 100589 91221
rect 100523 91156 100524 91220
rect 100588 91156 100589 91220
rect 100523 91155 100589 91156
rect 101811 91220 101877 91221
rect 101811 91156 101812 91220
rect 101876 91156 101877 91220
rect 101811 91155 101877 91156
rect 102550 90949 102610 94830
rect 103102 93870 103162 94830
rect 102734 93810 103162 93870
rect 102734 91221 102794 93810
rect 102731 91220 102797 91221
rect 102731 91156 102732 91220
rect 102796 91156 102797 91220
rect 102731 91155 102797 91156
rect 102547 90948 102613 90949
rect 102547 90884 102548 90948
rect 102612 90884 102613 90948
rect 102547 90883 102613 90884
rect 99234 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 99854 64894
rect 99234 64574 99854 64658
rect 99234 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 99854 64574
rect 99234 28894 99854 64338
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 68614 103574 93100
rect 104206 91765 104266 94830
rect 104203 91764 104269 91765
rect 104203 91700 104204 91764
rect 104268 91700 104269 91764
rect 104203 91699 104269 91700
rect 104574 91221 104634 94830
rect 105494 91221 105554 94830
rect 105678 92445 105738 94830
rect 106477 94828 106478 94892
rect 106542 94828 106543 94892
rect 106477 94827 106543 94828
rect 106616 94757 106676 95200
rect 106779 94892 106845 94893
rect 106779 94828 106780 94892
rect 106844 94828 106845 94892
rect 107704 94890 107764 95200
rect 108112 94890 108172 95200
rect 106779 94827 106845 94828
rect 107702 94830 107764 94890
rect 108070 94830 108172 94890
rect 109064 94890 109124 95200
rect 109472 94890 109532 95200
rect 109064 94830 109234 94890
rect 109472 94830 109602 94890
rect 106227 94756 106293 94757
rect 106227 94692 106228 94756
rect 106292 94692 106293 94756
rect 106227 94691 106293 94692
rect 106613 94756 106679 94757
rect 106613 94692 106614 94756
rect 106678 94692 106679 94756
rect 106613 94691 106679 94692
rect 105675 92444 105741 92445
rect 105675 92380 105676 92444
rect 105740 92380 105741 92444
rect 105675 92379 105741 92380
rect 106230 92037 106290 94691
rect 106227 92036 106293 92037
rect 106227 91972 106228 92036
rect 106292 91972 106293 92036
rect 106227 91971 106293 91972
rect 106782 91221 106842 94827
rect 107702 91221 107762 94830
rect 108070 93533 108130 94830
rect 108067 93532 108133 93533
rect 108067 93468 108068 93532
rect 108132 93468 108133 93532
rect 108067 93467 108133 93468
rect 109174 91357 109234 94830
rect 109171 91356 109237 91357
rect 109171 91292 109172 91356
rect 109236 91292 109237 91356
rect 109171 91291 109237 91292
rect 109542 91221 109602 94830
rect 110152 94757 110212 95200
rect 110696 94890 110756 95200
rect 111240 94890 111300 95200
rect 110646 94830 110756 94890
rect 111198 94830 111300 94890
rect 111920 94890 111980 95200
rect 112328 94890 112388 95200
rect 113144 94890 113204 95200
rect 113688 94890 113748 95200
rect 114368 94890 114428 95200
rect 111920 94830 111994 94890
rect 110149 94756 110215 94757
rect 110149 94692 110150 94756
rect 110214 94692 110215 94756
rect 110149 94691 110215 94692
rect 104571 91220 104637 91221
rect 104571 91156 104572 91220
rect 104636 91156 104637 91220
rect 104571 91155 104637 91156
rect 105491 91220 105557 91221
rect 105491 91156 105492 91220
rect 105556 91156 105557 91220
rect 105491 91155 105557 91156
rect 106779 91220 106845 91221
rect 106779 91156 106780 91220
rect 106844 91156 106845 91220
rect 106779 91155 106845 91156
rect 107699 91220 107765 91221
rect 107699 91156 107700 91220
rect 107764 91156 107765 91220
rect 107699 91155 107765 91156
rect 109539 91220 109605 91221
rect 109539 91156 109540 91220
rect 109604 91156 109605 91220
rect 109539 91155 109605 91156
rect 102954 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 103574 68614
rect 102954 68294 103574 68378
rect 102954 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 103574 68294
rect 102954 32614 103574 68058
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 75454 110414 93100
rect 110646 91221 110706 94830
rect 111198 92445 111258 94830
rect 111934 93669 111994 94830
rect 112302 94830 112388 94890
rect 113038 94830 113204 94890
rect 113406 94830 113748 94890
rect 114326 94830 114428 94890
rect 114776 94890 114836 95200
rect 115456 94890 115516 95200
rect 115864 94890 115924 95200
rect 114776 94830 114938 94890
rect 111931 93668 111997 93669
rect 111931 93604 111932 93668
rect 111996 93604 111997 93668
rect 111931 93603 111997 93604
rect 111195 92444 111261 92445
rect 111195 92380 111196 92444
rect 111260 92380 111261 92444
rect 111195 92379 111261 92380
rect 112302 91765 112362 94830
rect 113038 92170 113098 94830
rect 113406 93870 113466 94830
rect 113222 93810 113466 93870
rect 113222 92445 113282 93810
rect 113219 92444 113285 92445
rect 113219 92380 113220 92444
rect 113284 92380 113285 92444
rect 113219 92379 113285 92380
rect 113038 92110 113282 92170
rect 112299 91764 112365 91765
rect 112299 91700 112300 91764
rect 112364 91700 112365 91764
rect 112299 91699 112365 91700
rect 113222 91221 113282 92110
rect 110643 91220 110709 91221
rect 110643 91156 110644 91220
rect 110708 91156 110709 91220
rect 110643 91155 110709 91156
rect 113219 91220 113285 91221
rect 113219 91156 113220 91220
rect 113284 91156 113285 91220
rect 113219 91155 113285 91156
rect 109794 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 110414 75454
rect 109794 75134 110414 75218
rect 109794 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 110414 75134
rect 109794 39454 110414 74898
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 79174 114134 93100
rect 114326 91221 114386 94830
rect 114878 91765 114938 94830
rect 115430 94830 115516 94890
rect 115798 94830 115924 94890
rect 116680 94890 116740 95200
rect 117088 94890 117148 95200
rect 116680 94830 116778 94890
rect 115430 92445 115490 94830
rect 115427 92444 115493 92445
rect 115427 92380 115428 92444
rect 115492 92380 115493 92444
rect 115427 92379 115493 92380
rect 114875 91764 114941 91765
rect 114875 91700 114876 91764
rect 114940 91700 114941 91764
rect 114875 91699 114941 91700
rect 115798 91221 115858 94830
rect 116718 91357 116778 94830
rect 117086 94830 117148 94890
rect 117904 94890 117964 95200
rect 118176 94890 118236 95200
rect 119400 94890 119460 95200
rect 117904 94830 118066 94890
rect 118176 94830 118250 94890
rect 116715 91356 116781 91357
rect 116715 91292 116716 91356
rect 116780 91292 116781 91356
rect 116715 91291 116781 91292
rect 117086 91221 117146 94830
rect 114323 91220 114389 91221
rect 114323 91156 114324 91220
rect 114388 91156 114389 91220
rect 114323 91155 114389 91156
rect 115795 91220 115861 91221
rect 115795 91156 115796 91220
rect 115860 91156 115861 91220
rect 115795 91155 115861 91156
rect 117083 91220 117149 91221
rect 117083 91156 117084 91220
rect 117148 91156 117149 91220
rect 117083 91155 117149 91156
rect 113514 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 114134 79174
rect 113514 78854 114134 78938
rect 113514 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 114134 78854
rect 113514 43174 114134 78618
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 82894 117854 93100
rect 118006 92445 118066 94830
rect 118003 92444 118069 92445
rect 118003 92380 118004 92444
rect 118068 92380 118069 92444
rect 118003 92379 118069 92380
rect 118190 91221 118250 94830
rect 119294 94830 119460 94890
rect 119536 94890 119596 95200
rect 120216 94890 120276 95200
rect 120624 94890 120684 95200
rect 121712 94890 121772 95200
rect 119536 94830 119722 94890
rect 119294 91221 119354 94830
rect 119662 91357 119722 94830
rect 120214 94830 120276 94890
rect 120582 94830 120684 94890
rect 121686 94830 121772 94890
rect 121984 94890 122044 95200
rect 122800 94890 122860 95200
rect 123208 94890 123268 95200
rect 121984 94830 122114 94890
rect 122800 94830 123034 94890
rect 119659 91356 119725 91357
rect 119659 91292 119660 91356
rect 119724 91292 119725 91356
rect 119659 91291 119725 91292
rect 120214 91221 120274 94830
rect 120582 91765 120642 94830
rect 121686 93533 121746 94830
rect 121683 93532 121749 93533
rect 121683 93468 121684 93532
rect 121748 93468 121749 93532
rect 121683 93467 121749 93468
rect 120579 91764 120645 91765
rect 120579 91700 120580 91764
rect 120644 91700 120645 91764
rect 120579 91699 120645 91700
rect 118187 91220 118253 91221
rect 118187 91156 118188 91220
rect 118252 91156 118253 91220
rect 118187 91155 118253 91156
rect 119291 91220 119357 91221
rect 119291 91156 119292 91220
rect 119356 91156 119357 91220
rect 119291 91155 119357 91156
rect 120211 91220 120277 91221
rect 120211 91156 120212 91220
rect 120276 91156 120277 91220
rect 120211 91155 120277 91156
rect 117234 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 117854 82894
rect 117234 82574 117854 82658
rect 117234 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 117854 82574
rect 117234 46894 117854 82338
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 86614 121574 93100
rect 122054 91221 122114 94830
rect 122974 93870 123034 94830
rect 122606 93810 123034 93870
rect 123158 94830 123268 94890
rect 124024 94890 124084 95200
rect 124432 94890 124492 95200
rect 124024 94830 124138 94890
rect 124432 94830 124506 94890
rect 122606 91490 122666 93810
rect 123158 93533 123218 94830
rect 123155 93532 123221 93533
rect 123155 93468 123156 93532
rect 123220 93468 123221 93532
rect 123155 93467 123221 93468
rect 122787 91492 122853 91493
rect 122787 91490 122788 91492
rect 122606 91430 122788 91490
rect 122787 91428 122788 91430
rect 122852 91428 122853 91492
rect 122787 91427 122853 91428
rect 124078 91221 124138 94830
rect 124446 91221 124506 94830
rect 125384 94757 125444 95200
rect 125656 94890 125716 95200
rect 126472 94890 126532 95200
rect 125656 94830 125794 94890
rect 125381 94756 125447 94757
rect 125381 94692 125382 94756
rect 125446 94692 125447 94756
rect 125381 94691 125447 94692
rect 125734 92309 125794 94830
rect 126470 94830 126532 94890
rect 126608 94890 126668 95200
rect 128104 94890 128164 95200
rect 126608 94830 126714 94890
rect 125731 92308 125797 92309
rect 125731 92244 125732 92308
rect 125796 92244 125797 92308
rect 125731 92243 125797 92244
rect 126470 91221 126530 94830
rect 126654 91221 126714 94830
rect 127574 94830 128164 94890
rect 129328 94890 129388 95200
rect 130688 94890 130748 95200
rect 131912 94890 131972 95200
rect 133136 94890 133196 95200
rect 129328 94830 129474 94890
rect 130688 94830 130762 94890
rect 131912 94830 132050 94890
rect 127574 92173 127634 94830
rect 127571 92172 127637 92173
rect 127571 92108 127572 92172
rect 127636 92108 127637 92172
rect 127571 92107 127637 92108
rect 122051 91220 122117 91221
rect 122051 91156 122052 91220
rect 122116 91156 122117 91220
rect 122051 91155 122117 91156
rect 124075 91220 124141 91221
rect 124075 91156 124076 91220
rect 124140 91156 124141 91220
rect 124075 91155 124141 91156
rect 124443 91220 124509 91221
rect 124443 91156 124444 91220
rect 124508 91156 124509 91220
rect 124443 91155 124509 91156
rect 126467 91220 126533 91221
rect 126467 91156 126468 91220
rect 126532 91156 126533 91220
rect 126467 91155 126533 91156
rect 126651 91220 126717 91221
rect 126651 91156 126652 91220
rect 126716 91156 126717 91220
rect 126651 91155 126717 91156
rect 120954 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 121574 86614
rect 120954 86294 121574 86378
rect 120954 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 121574 86294
rect 120954 50614 121574 86058
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 93100
rect 129414 91221 129474 94830
rect 130702 91221 130762 94830
rect 131990 93805 132050 94830
rect 133094 94830 133196 94890
rect 134360 94890 134420 95200
rect 135584 94890 135644 95200
rect 151307 94892 151373 94893
rect 134360 94830 134442 94890
rect 135584 94830 136098 94890
rect 131987 93804 132053 93805
rect 131987 93740 131988 93804
rect 132052 93740 132053 93804
rect 131987 93739 132053 93740
rect 129411 91220 129477 91221
rect 129411 91156 129412 91220
rect 129476 91156 129477 91220
rect 129411 91155 129477 91156
rect 130699 91220 130765 91221
rect 130699 91156 130700 91220
rect 130764 91156 130765 91220
rect 130699 91155 130765 91156
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 61174 132134 93100
rect 133094 91221 133154 94830
rect 134382 91221 134442 94830
rect 133091 91220 133157 91221
rect 133091 91156 133092 91220
rect 133156 91156 133157 91220
rect 133091 91155 133157 91156
rect 134379 91220 134445 91221
rect 134379 91156 134380 91220
rect 134444 91156 134445 91220
rect 134379 91155 134445 91156
rect 131514 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 132134 61174
rect 131514 60854 132134 60938
rect 131514 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 132134 60854
rect 131514 25174 132134 60618
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 64894 135854 93100
rect 136038 92445 136098 94830
rect 151307 94828 151308 94892
rect 151372 94828 151373 94892
rect 151307 94827 151373 94828
rect 136035 92444 136101 92445
rect 136035 92380 136036 92444
rect 136100 92380 136101 92444
rect 136035 92379 136101 92380
rect 135234 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 135854 64894
rect 135234 64574 135854 64658
rect 135234 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 135854 64574
rect 135234 28894 135854 64338
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 68614 139574 93100
rect 138954 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 139574 68614
rect 138954 68294 139574 68378
rect 138954 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 139574 68294
rect 138954 32614 139574 68058
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 75454 146414 93100
rect 145794 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 146414 75454
rect 145794 75134 146414 75218
rect 145794 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 146414 75134
rect 145794 39454 146414 74898
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 79174 150134 93100
rect 151310 91357 151370 94827
rect 151496 94754 151556 95200
rect 151494 94694 151556 94754
rect 151632 94754 151692 95200
rect 151768 94893 151828 95200
rect 151765 94892 151831 94893
rect 151765 94828 151766 94892
rect 151830 94828 151831 94892
rect 151765 94827 151831 94828
rect 151904 94754 151964 95200
rect 151632 94694 151738 94754
rect 151904 94694 152106 94754
rect 151494 91493 151554 94694
rect 151491 91492 151557 91493
rect 151491 91428 151492 91492
rect 151556 91428 151557 91492
rect 151491 91427 151557 91428
rect 151307 91356 151373 91357
rect 151307 91292 151308 91356
rect 151372 91292 151373 91356
rect 151307 91291 151373 91292
rect 151678 91221 151738 94694
rect 152046 92445 152106 94694
rect 166214 94485 166274 132771
rect 166395 103868 166461 103869
rect 166395 103804 166396 103868
rect 166460 103804 166461 103868
rect 166395 103803 166461 103804
rect 166211 94484 166277 94485
rect 166211 94420 166212 94484
rect 166276 94420 166277 94484
rect 166211 94419 166277 94420
rect 152043 92444 152109 92445
rect 152043 92380 152044 92444
rect 152108 92380 152109 92444
rect 152043 92379 152109 92380
rect 151675 91220 151741 91221
rect 151675 91156 151676 91220
rect 151740 91156 151741 91220
rect 151675 91155 151741 91156
rect 149514 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 150134 79174
rect 149514 78854 150134 78938
rect 149514 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 150134 78854
rect 149514 43174 150134 78618
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 82894 153854 93100
rect 153234 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 153854 82894
rect 153234 82574 153854 82658
rect 153234 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 153854 82574
rect 153234 46894 153854 82338
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 86614 157574 93100
rect 156954 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 157574 86614
rect 156954 86294 157574 86378
rect 156954 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 157574 86294
rect 156954 50614 157574 86058
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 93100
rect 166398 84013 166458 103803
rect 166395 84012 166461 84013
rect 166395 83948 166396 84012
rect 166460 83948 166461 84012
rect 166395 83947 166461 83948
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 166950 13021 167010 377299
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 168971 258092 169037 258093
rect 168971 258028 168972 258092
rect 169036 258028 169037 258092
rect 168971 258027 169037 258028
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 205174 168134 240618
rect 167514 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 168134 205174
rect 167514 204854 168134 204938
rect 167514 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 168134 204854
rect 167514 169174 168134 204618
rect 168974 185605 169034 258027
rect 169523 194444 169589 194445
rect 169523 194380 169524 194444
rect 169588 194380 169589 194444
rect 169523 194379 169589 194380
rect 168971 185604 169037 185605
rect 168971 185540 168972 185604
rect 169036 185540 169037 185604
rect 168971 185539 169037 185540
rect 167514 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 168134 169174
rect 167514 168854 168134 168938
rect 167514 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 168134 168854
rect 167514 133174 168134 168618
rect 169526 142765 169586 194379
rect 169523 142764 169589 142765
rect 169523 142700 169524 142764
rect 169588 142700 169589 142764
rect 169523 142699 169589 142700
rect 167514 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 168134 133174
rect 167514 132854 168134 132938
rect 167514 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 168134 132854
rect 167514 97174 168134 132618
rect 168971 101420 169037 101421
rect 168971 101356 168972 101420
rect 169036 101356 169037 101420
rect 168971 101355 169037 101356
rect 167514 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 168134 97174
rect 167514 96854 168134 96938
rect 167514 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 168134 96854
rect 167514 61174 168134 96618
rect 168419 96660 168485 96661
rect 168419 96596 168420 96660
rect 168484 96596 168485 96660
rect 168419 96595 168485 96596
rect 167514 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 168134 61174
rect 167514 60854 168134 60938
rect 167514 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 168134 60854
rect 167514 25174 168134 60618
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 166947 13020 167013 13021
rect 166947 12956 166948 13020
rect 167012 12956 167013 13020
rect 166947 12955 167013 12956
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 -3226 168134 24618
rect 168422 15877 168482 96595
rect 168974 81429 169034 101355
rect 168971 81428 169037 81429
rect 168971 81364 168972 81428
rect 169036 81364 169037 81428
rect 168971 81363 169037 81364
rect 169710 43485 169770 586467
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 460894 171854 496338
rect 171234 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 171854 460894
rect 171234 460574 171854 460658
rect 171234 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 171854 460574
rect 171234 424894 171854 460338
rect 171234 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 171854 424894
rect 171234 424574 171854 424658
rect 171234 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 171854 424574
rect 171234 388894 171854 424338
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 464614 175574 500058
rect 174954 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 175574 464614
rect 174954 464294 175574 464378
rect 174954 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 175574 464294
rect 174954 428614 175574 464058
rect 174954 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 175574 428614
rect 174954 428294 175574 428378
rect 174954 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 175574 428294
rect 174954 392614 175574 428058
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 471454 182414 506898
rect 181794 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 182414 471454
rect 181794 471134 182414 471218
rect 181794 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 182414 471134
rect 181794 435454 182414 470898
rect 181794 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 182414 435454
rect 181794 435134 182414 435218
rect 181794 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 182414 435134
rect 181794 399454 182414 434898
rect 181794 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 182414 399454
rect 181794 399134 182414 399218
rect 181794 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 182414 399134
rect 181794 363454 182414 398898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 475174 186134 510618
rect 185514 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 186134 475174
rect 185514 474854 186134 474938
rect 185514 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 186134 474854
rect 185514 439174 186134 474618
rect 185514 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 186134 439174
rect 185514 438854 186134 438938
rect 185514 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 186134 438854
rect 185514 403174 186134 438618
rect 185514 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 186134 403174
rect 185514 402854 186134 402938
rect 185514 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 186134 402854
rect 185514 367174 186134 402618
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 184059 364444 184125 364445
rect 184059 364380 184060 364444
rect 184124 364380 184125 364444
rect 184059 364379 184125 364380
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 178539 350708 178605 350709
rect 178539 350644 178540 350708
rect 178604 350644 178605 350708
rect 178539 350643 178605 350644
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 173019 287196 173085 287197
rect 173019 287132 173020 287196
rect 173084 287132 173085 287196
rect 173019 287131 173085 287132
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 208894 171854 244338
rect 171234 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 171854 208894
rect 171234 208574 171854 208658
rect 171234 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 171854 208574
rect 171234 172894 171854 208338
rect 171234 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 171854 172894
rect 171234 172574 171854 172658
rect 171234 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 171854 172574
rect 171234 136894 171854 172338
rect 171234 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 171854 136894
rect 171234 136574 171854 136658
rect 171234 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 171854 136574
rect 171234 100894 171854 136338
rect 171234 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 171854 100894
rect 171234 100574 171854 100658
rect 171234 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 171854 100574
rect 171234 64894 171854 100338
rect 171234 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 171854 64894
rect 171234 64574 171854 64658
rect 171234 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 171854 64574
rect 169707 43484 169773 43485
rect 169707 43420 169708 43484
rect 169772 43420 169773 43484
rect 169707 43419 169773 43420
rect 171234 28894 171854 64338
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 168419 15876 168485 15877
rect 168419 15812 168420 15876
rect 168484 15812 168485 15876
rect 168419 15811 168485 15812
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 -5146 171854 28338
rect 173022 22813 173082 287131
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 212614 175574 248058
rect 174954 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 175574 212614
rect 174954 212294 175574 212378
rect 174954 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 175574 212294
rect 174954 176614 175574 212058
rect 174954 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 175574 176614
rect 174954 176294 175574 176378
rect 174954 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 175574 176294
rect 174954 140614 175574 176058
rect 174954 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 175574 140614
rect 174954 140294 175574 140378
rect 174954 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 175574 140294
rect 174954 104614 175574 140058
rect 178542 133109 178602 350643
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 184062 280805 184122 364379
rect 185514 331174 186134 366618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 478894 189854 514338
rect 189234 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 189854 478894
rect 189234 478574 189854 478658
rect 189234 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 189854 478574
rect 189234 442894 189854 478338
rect 189234 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 189854 442894
rect 189234 442574 189854 442658
rect 189234 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 189854 442574
rect 189234 406894 189854 442338
rect 189234 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 189854 406894
rect 189234 406574 189854 406658
rect 189234 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 189854 406574
rect 189234 370894 189854 406338
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 186819 345268 186885 345269
rect 186819 345204 186820 345268
rect 186884 345204 186885 345268
rect 186819 345203 186885 345204
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 184059 280804 184125 280805
rect 184059 280740 184060 280804
rect 184124 280740 184125 280804
rect 184059 280739 184125 280740
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 219454 182414 254898
rect 181794 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 182414 219454
rect 181794 219134 182414 219218
rect 181794 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 182414 219134
rect 181794 183454 182414 218898
rect 181794 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 182414 183454
rect 181794 183134 182414 183218
rect 181794 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 182414 183134
rect 181794 147454 182414 182898
rect 181794 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 182414 147454
rect 181794 147134 182414 147218
rect 181794 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 182414 147134
rect 178539 133108 178605 133109
rect 178539 133044 178540 133108
rect 178604 133044 178605 133108
rect 178539 133043 178605 133044
rect 174954 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 175574 104614
rect 174954 104294 175574 104378
rect 174954 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 175574 104294
rect 174954 68614 175574 104058
rect 174954 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 175574 68614
rect 174954 68294 175574 68378
rect 174954 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 175574 68294
rect 174954 32614 175574 68058
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 173019 22812 173085 22813
rect 173019 22748 173020 22812
rect 173084 22748 173085 22812
rect 173019 22747 173085 22748
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 111454 182414 146898
rect 181794 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 182414 111454
rect 181794 111134 182414 111218
rect 181794 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 182414 111134
rect 181794 75454 182414 110898
rect 181794 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 182414 75454
rect 181794 75134 182414 75218
rect 181794 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 182414 75134
rect 181794 39454 182414 74898
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 223174 186134 258618
rect 185514 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 186134 223174
rect 185514 222854 186134 222938
rect 185514 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 186134 222854
rect 185514 187174 186134 222618
rect 185514 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 186134 187174
rect 185514 186854 186134 186938
rect 185514 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 186134 186854
rect 185514 151174 186134 186618
rect 185514 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 186134 151174
rect 185514 150854 186134 150938
rect 185514 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 186134 150854
rect 185514 115174 186134 150618
rect 185514 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 186134 115174
rect 185514 114854 186134 114938
rect 185514 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 186134 114854
rect 185514 79174 186134 114618
rect 185514 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 186134 79174
rect 185514 78854 186134 78938
rect 185514 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 186134 78854
rect 185514 43174 186134 78618
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 186822 2141 186882 345203
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 188291 301068 188357 301069
rect 188291 301004 188292 301068
rect 188356 301004 188357 301068
rect 188291 301003 188357 301004
rect 188294 13021 188354 301003
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 226894 189854 262338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 482614 193574 518058
rect 192954 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 193574 482614
rect 192954 482294 193574 482378
rect 192954 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 193574 482294
rect 192954 446614 193574 482058
rect 192954 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 193574 446614
rect 192954 446294 193574 446378
rect 192954 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 193574 446294
rect 192954 410614 193574 446058
rect 192954 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 193574 410614
rect 192954 410294 193574 410378
rect 192954 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 193574 410294
rect 192954 374614 193574 410058
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203011 346628 203077 346629
rect 203011 346564 203012 346628
rect 203076 346564 203077 346628
rect 203011 346563 203077 346564
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 195099 313308 195165 313309
rect 195099 313244 195100 313308
rect 195164 313244 195165 313308
rect 195099 313243 195165 313244
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 191603 241636 191669 241637
rect 191603 241572 191604 241636
rect 191668 241572 191669 241636
rect 191603 241571 191669 241572
rect 189234 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 189854 226894
rect 189234 226574 189854 226658
rect 189234 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 189854 226574
rect 189234 190894 189854 226338
rect 191606 211173 191666 241571
rect 192954 230614 193574 266058
rect 193811 254420 193877 254421
rect 193811 254356 193812 254420
rect 193876 254356 193877 254420
rect 193811 254355 193877 254356
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 191603 211172 191669 211173
rect 191603 211108 191604 211172
rect 191668 211108 191669 211172
rect 191603 211107 191669 211108
rect 189234 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 189854 190894
rect 189234 190574 189854 190658
rect 189234 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 189854 190574
rect 189234 154894 189854 190338
rect 189234 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 189854 154894
rect 189234 154574 189854 154658
rect 189234 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 189854 154574
rect 189234 118894 189854 154338
rect 189234 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 189854 118894
rect 189234 118574 189854 118658
rect 189234 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 189854 118574
rect 189234 82894 189854 118338
rect 189234 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 189854 82894
rect 189234 82574 189854 82658
rect 189234 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 189854 82574
rect 189234 46894 189854 82338
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 188291 13020 188357 13021
rect 188291 12956 188292 13020
rect 188356 12956 188357 13020
rect 188291 12955 188357 12956
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 186819 2140 186885 2141
rect 186819 2076 186820 2140
rect 186884 2076 186885 2140
rect 186819 2075 186885 2076
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 194614 193574 230058
rect 193814 220829 193874 254355
rect 193811 220828 193877 220829
rect 193811 220764 193812 220828
rect 193876 220764 193877 220828
rect 193811 220763 193877 220764
rect 192954 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 193574 194614
rect 192954 194294 193574 194378
rect 192954 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 193574 194294
rect 192954 158614 193574 194058
rect 192954 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 193574 158614
rect 192954 158294 193574 158378
rect 192954 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 193574 158294
rect 192954 122614 193574 158058
rect 192954 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 193574 122614
rect 192954 122294 193574 122378
rect 192954 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 193574 122294
rect 192954 86614 193574 122058
rect 192954 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 193574 86614
rect 192954 86294 193574 86378
rect 192954 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 193574 86294
rect 192954 50614 193574 86058
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 195102 14517 195162 313243
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 197859 292636 197925 292637
rect 197859 292572 197860 292636
rect 197924 292572 197925 292636
rect 197859 292571 197925 292572
rect 195467 286380 195533 286381
rect 195467 286316 195468 286380
rect 195532 286316 195533 286380
rect 195467 286315 195533 286316
rect 195470 245989 195530 286315
rect 196571 280804 196637 280805
rect 196571 280740 196572 280804
rect 196636 280740 196637 280804
rect 196571 280739 196637 280740
rect 195467 245988 195533 245989
rect 195467 245924 195468 245988
rect 195532 245924 195533 245988
rect 195467 245923 195533 245924
rect 195283 243812 195349 243813
rect 195283 243748 195284 243812
rect 195348 243748 195349 243812
rect 195283 243747 195349 243748
rect 195286 235653 195346 243747
rect 196574 235653 196634 280739
rect 197862 277269 197922 292571
rect 199331 291548 199397 291549
rect 199331 291484 199332 291548
rect 199396 291484 199397 291548
rect 199331 291483 199397 291484
rect 198779 284612 198845 284613
rect 198779 284548 198780 284612
rect 198844 284548 198845 284612
rect 198779 284547 198845 284548
rect 197859 277268 197925 277269
rect 197859 277204 197860 277268
rect 197924 277204 197925 277268
rect 197859 277203 197925 277204
rect 198782 265573 198842 284547
rect 199334 279445 199394 291483
rect 199794 286182 200414 308898
rect 200619 284612 200685 284613
rect 200619 284548 200620 284612
rect 200684 284548 200685 284612
rect 200619 284547 200685 284548
rect 199331 279444 199397 279445
rect 199331 279380 199332 279444
rect 199396 279380 199397 279444
rect 199331 279379 199397 279380
rect 198779 265572 198845 265573
rect 198779 265508 198780 265572
rect 198844 265508 198845 265572
rect 198779 265507 198845 265508
rect 198779 259452 198845 259453
rect 198779 259388 198780 259452
rect 198844 259388 198845 259452
rect 198779 259387 198845 259388
rect 198782 247077 198842 259387
rect 198779 247076 198845 247077
rect 198779 247012 198780 247076
rect 198844 247012 198845 247076
rect 198779 247011 198845 247012
rect 199883 247076 199949 247077
rect 199883 247012 199884 247076
rect 199948 247012 199949 247076
rect 199883 247011 199949 247012
rect 199886 240410 199946 247011
rect 199886 240350 200498 240410
rect 200438 240141 200498 240350
rect 200251 240140 200317 240141
rect 200251 240076 200252 240140
rect 200316 240076 200317 240140
rect 200251 240075 200317 240076
rect 200435 240140 200501 240141
rect 200435 240076 200436 240140
rect 200500 240076 200501 240140
rect 200435 240075 200501 240076
rect 200254 239733 200314 240075
rect 200251 239732 200317 239733
rect 200251 239668 200252 239732
rect 200316 239668 200317 239732
rect 200251 239667 200317 239668
rect 199794 237454 200414 238182
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 195283 235652 195349 235653
rect 195283 235588 195284 235652
rect 195348 235588 195349 235652
rect 195283 235587 195349 235588
rect 196571 235652 196637 235653
rect 196571 235588 196572 235652
rect 196636 235588 196637 235652
rect 196571 235587 196637 235588
rect 199794 201454 200414 236898
rect 199794 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 200414 201454
rect 199794 201134 200414 201218
rect 199794 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 200414 201134
rect 199794 165454 200414 200898
rect 199794 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 200414 165454
rect 199794 165134 200414 165218
rect 199794 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 200414 165134
rect 199794 129454 200414 164898
rect 199794 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 200414 129454
rect 199794 129134 200414 129218
rect 199794 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 200414 129134
rect 199794 93454 200414 128898
rect 200622 93669 200682 284547
rect 203014 238645 203074 346563
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 286182 204134 312618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 208899 367164 208965 367165
rect 208899 367100 208900 367164
rect 208964 367100 208965 367164
rect 208899 367099 208965 367100
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207979 327724 208045 327725
rect 207979 327660 207980 327724
rect 208044 327660 208045 327724
rect 207979 327659 208045 327660
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 286182 207854 316338
rect 205403 283932 205469 283933
rect 205403 283868 205404 283932
rect 205468 283868 205469 283932
rect 205403 283867 205469 283868
rect 204408 255454 204728 255486
rect 204408 255218 204450 255454
rect 204686 255218 204728 255454
rect 204408 255134 204728 255218
rect 204408 254898 204450 255134
rect 204686 254898 204728 255134
rect 204408 254866 204728 254898
rect 203011 238644 203077 238645
rect 203011 238580 203012 238644
rect 203076 238580 203077 238644
rect 203011 238579 203077 238580
rect 203514 205174 204134 238182
rect 203514 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 204134 205174
rect 203514 204854 204134 204938
rect 203514 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 204134 204854
rect 203514 169174 204134 204618
rect 203514 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 204134 169174
rect 203514 168854 204134 168938
rect 203514 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 204134 168854
rect 203514 133174 204134 168618
rect 203514 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 204134 133174
rect 203514 132854 204134 132938
rect 203514 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 204134 132854
rect 203514 97174 204134 132618
rect 203514 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 204134 97174
rect 203514 96854 204134 96938
rect 203514 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 204134 96854
rect 200619 93668 200685 93669
rect 200619 93604 200620 93668
rect 200684 93604 200685 93668
rect 200619 93603 200685 93604
rect 199794 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 200414 93454
rect 199794 93134 200414 93218
rect 199794 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 200414 93134
rect 199794 57454 200414 92898
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 195099 14516 195165 14517
rect 195099 14452 195100 14516
rect 195164 14452 195165 14516
rect 195099 14451 195165 14452
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 61174 204134 96618
rect 205406 95165 205466 283867
rect 207982 239461 208042 327659
rect 207979 239460 208045 239461
rect 207979 239396 207980 239460
rect 208044 239396 208045 239460
rect 207979 239395 208045 239396
rect 207234 208894 207854 238182
rect 208902 237285 208962 367099
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 471454 218414 506898
rect 217794 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 218414 471454
rect 217794 471134 218414 471218
rect 217794 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 218414 471134
rect 217794 435454 218414 470898
rect 217794 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 218414 435454
rect 217794 435134 218414 435218
rect 217794 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 218414 435134
rect 217794 399454 218414 434898
rect 217794 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 218414 399454
rect 217794 399134 218414 399218
rect 217794 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 218414 399134
rect 217794 363454 218414 398898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 475174 222134 510618
rect 221514 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 222134 475174
rect 221514 474854 222134 474938
rect 221514 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 222134 474854
rect 221514 439174 222134 474618
rect 221514 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 222134 439174
rect 221514 438854 222134 438938
rect 221514 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 222134 438854
rect 221514 403174 222134 438618
rect 221514 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 222134 403174
rect 221514 402854 222134 402938
rect 221514 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 222134 402854
rect 221514 367174 222134 402618
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 218651 365804 218717 365805
rect 218651 365740 218652 365804
rect 218716 365740 218717 365804
rect 218651 365739 218717 365740
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 212579 334388 212645 334389
rect 212579 334324 212580 334388
rect 212644 334324 212645 334388
rect 212579 334323 212645 334324
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 286182 211574 320058
rect 210739 285836 210805 285837
rect 210739 285772 210740 285836
rect 210804 285772 210805 285836
rect 210739 285771 210805 285772
rect 208899 237284 208965 237285
rect 208899 237220 208900 237284
rect 208964 237220 208965 237284
rect 208899 237219 208965 237220
rect 207234 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 207854 208894
rect 207234 208574 207854 208658
rect 207234 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 207854 208574
rect 207234 172894 207854 208338
rect 210742 207909 210802 285771
rect 212395 283932 212461 283933
rect 212395 283868 212396 283932
rect 212460 283868 212461 283932
rect 212395 283867 212461 283868
rect 210954 212614 211574 238182
rect 210954 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 211574 212614
rect 210954 212294 211574 212378
rect 210954 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 211574 212294
rect 210739 207908 210805 207909
rect 210739 207844 210740 207908
rect 210804 207844 210805 207908
rect 210739 207843 210805 207844
rect 207234 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 207854 172894
rect 207234 172574 207854 172658
rect 207234 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 207854 172574
rect 207234 136894 207854 172338
rect 207234 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 207854 136894
rect 207234 136574 207854 136658
rect 207234 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 207854 136574
rect 207234 100894 207854 136338
rect 207234 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 207854 100894
rect 207234 100574 207854 100658
rect 207234 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 207854 100574
rect 205403 95164 205469 95165
rect 205403 95100 205404 95164
rect 205468 95100 205469 95164
rect 205403 95099 205469 95100
rect 203514 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 204134 61174
rect 203514 60854 204134 60938
rect 203514 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 204134 60854
rect 203514 25174 204134 60618
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 64894 207854 100338
rect 207234 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 207854 64894
rect 207234 64574 207854 64658
rect 207234 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 207854 64574
rect 207234 28894 207854 64338
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 176614 211574 212058
rect 210954 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 211574 176614
rect 210954 176294 211574 176378
rect 210954 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 211574 176294
rect 210954 140614 211574 176058
rect 210954 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 211574 140614
rect 210954 140294 211574 140378
rect 210954 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 211574 140294
rect 210954 104614 211574 140058
rect 210954 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 211574 104614
rect 210954 104294 211574 104378
rect 210954 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 211574 104294
rect 210954 68614 211574 104058
rect 212398 95029 212458 283867
rect 212582 238645 212642 334323
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 214051 297532 214117 297533
rect 214051 297468 214052 297532
rect 214116 297468 214117 297532
rect 214051 297467 214117 297468
rect 214054 238645 214114 297467
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 286182 218414 290898
rect 214419 283932 214485 283933
rect 214419 283868 214420 283932
rect 214484 283868 214485 283932
rect 214419 283867 214485 283868
rect 215891 283932 215957 283933
rect 215891 283868 215892 283932
rect 215956 283868 215957 283932
rect 215891 283867 215957 283868
rect 216627 283932 216693 283933
rect 216627 283868 216628 283932
rect 216692 283868 216693 283932
rect 216627 283867 216693 283868
rect 212579 238644 212645 238645
rect 212579 238580 212580 238644
rect 212644 238580 212645 238644
rect 212579 238579 212645 238580
rect 214051 238644 214117 238645
rect 214051 238580 214052 238644
rect 214116 238580 214117 238644
rect 214051 238579 214117 238580
rect 214422 211173 214482 283867
rect 215894 226405 215954 283867
rect 216630 230485 216690 283867
rect 218654 240141 218714 365739
rect 221514 331174 222134 366618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 478894 225854 514338
rect 225234 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 225854 478894
rect 225234 478574 225854 478658
rect 225234 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 225854 478574
rect 225234 442894 225854 478338
rect 225234 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 225854 442894
rect 225234 442574 225854 442658
rect 225234 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 225854 442574
rect 225234 406894 225854 442338
rect 225234 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 225854 406894
rect 225234 406574 225854 406658
rect 225234 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 225854 406574
rect 225234 370894 225854 406338
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 223619 347852 223685 347853
rect 223619 347788 223620 347852
rect 223684 347788 223685 347852
rect 223619 347787 223685 347788
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 286182 222134 294618
rect 223622 285701 223682 347787
rect 225234 334894 225854 370338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 482614 229574 518058
rect 228954 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 229574 482614
rect 228954 482294 229574 482378
rect 228954 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 229574 482294
rect 228954 446614 229574 482058
rect 228954 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 229574 446614
rect 228954 446294 229574 446378
rect 228954 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 229574 446294
rect 228954 410614 229574 446058
rect 228954 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 229574 410614
rect 228954 410294 229574 410378
rect 228954 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 229574 410294
rect 228954 374614 229574 410058
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228219 341052 228285 341053
rect 228219 340988 228220 341052
rect 228284 340988 228285 341052
rect 228219 340987 228285 340988
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 286182 225854 298338
rect 223619 285700 223685 285701
rect 223619 285636 223620 285700
rect 223684 285636 223685 285700
rect 223619 285635 223685 285636
rect 222699 284068 222765 284069
rect 222699 284004 222700 284068
rect 222764 284004 222765 284068
rect 222699 284003 222765 284004
rect 226931 284068 226997 284069
rect 226931 284004 226932 284068
rect 226996 284004 226997 284068
rect 226931 284003 226997 284004
rect 221227 283932 221293 283933
rect 221227 283868 221228 283932
rect 221292 283868 221293 283932
rect 221227 283867 221293 283868
rect 219768 273454 220088 273486
rect 219768 273218 219810 273454
rect 220046 273218 220088 273454
rect 219768 273134 220088 273218
rect 219768 272898 219810 273134
rect 220046 272898 220088 273134
rect 219768 272866 220088 272898
rect 218651 240140 218717 240141
rect 218651 240076 218652 240140
rect 218716 240076 218717 240140
rect 218651 240075 218717 240076
rect 216627 230484 216693 230485
rect 216627 230420 216628 230484
rect 216692 230420 216693 230484
rect 216627 230419 216693 230420
rect 215891 226404 215957 226405
rect 215891 226340 215892 226404
rect 215956 226340 215957 226404
rect 215891 226339 215957 226340
rect 216630 222869 216690 230419
rect 216627 222868 216693 222869
rect 216627 222804 216628 222868
rect 216692 222804 216693 222868
rect 216627 222803 216693 222804
rect 217794 219454 218414 238182
rect 217794 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 218414 219454
rect 217794 219134 218414 219218
rect 217794 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 218414 219134
rect 214419 211172 214485 211173
rect 214419 211108 214420 211172
rect 214484 211108 214485 211172
rect 214419 211107 214485 211108
rect 217794 183454 218414 218898
rect 221230 188597 221290 283867
rect 221514 223174 222134 238182
rect 221514 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 222134 223174
rect 221514 222854 222134 222938
rect 221514 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 222134 222854
rect 221227 188596 221293 188597
rect 221227 188532 221228 188596
rect 221292 188532 221293 188596
rect 221227 188531 221293 188532
rect 217794 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 218414 183454
rect 217794 183134 218414 183218
rect 217794 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 218414 183134
rect 217794 178000 218414 182898
rect 221514 187174 222134 222618
rect 222702 198253 222762 284003
rect 224723 283932 224789 283933
rect 224723 283868 224724 283932
rect 224788 283868 224789 283932
rect 224723 283867 224789 283868
rect 226195 283932 226261 283933
rect 226195 283868 226196 283932
rect 226260 283868 226261 283932
rect 226195 283867 226261 283868
rect 223619 225996 223685 225997
rect 223619 225932 223620 225996
rect 223684 225932 223685 225996
rect 223619 225931 223685 225932
rect 222699 198252 222765 198253
rect 222699 198188 222700 198252
rect 222764 198188 222765 198252
rect 222699 198187 222765 198188
rect 221514 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 222134 187174
rect 221514 186854 222134 186938
rect 221514 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 222134 186854
rect 221514 178000 222134 186618
rect 223622 175949 223682 225931
rect 224726 196757 224786 283867
rect 225234 226894 225854 238182
rect 225234 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 225854 226894
rect 225234 226574 225854 226658
rect 225234 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 225854 226574
rect 224723 196756 224789 196757
rect 224723 196692 224724 196756
rect 224788 196692 224789 196756
rect 224723 196691 224789 196692
rect 225234 190894 225854 226338
rect 225234 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 225854 190894
rect 225234 190574 225854 190658
rect 225234 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 225854 190574
rect 225234 178000 225854 190338
rect 226198 176629 226258 283867
rect 226934 183021 226994 284003
rect 228222 240141 228282 340987
rect 228954 338614 229574 374058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 453454 236414 488898
rect 235794 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 236414 453454
rect 235794 453134 236414 453218
rect 235794 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 236414 453134
rect 235794 417454 236414 452898
rect 235794 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 236414 417454
rect 235794 417134 236414 417218
rect 235794 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 236414 417134
rect 235794 381454 236414 416898
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 232451 354924 232517 354925
rect 232451 354860 232452 354924
rect 232516 354860 232517 354924
rect 232451 354859 232517 354860
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 286182 229574 302058
rect 230243 283932 230309 283933
rect 230243 283868 230244 283932
rect 230308 283868 230309 283932
rect 230243 283867 230309 283868
rect 231715 283932 231781 283933
rect 231715 283868 231716 283932
rect 231780 283868 231781 283932
rect 231715 283867 231781 283868
rect 228219 240140 228285 240141
rect 228219 240076 228220 240140
rect 228284 240076 228285 240140
rect 228219 240075 228285 240076
rect 228954 230614 229574 238182
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 230246 225181 230306 283867
rect 230243 225180 230309 225181
rect 230243 225116 230244 225180
rect 230308 225116 230309 225180
rect 230243 225115 230309 225116
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 226931 183020 226997 183021
rect 226931 182956 226932 183020
rect 226996 182956 226997 183020
rect 226931 182955 226997 182956
rect 228954 178000 229574 194058
rect 230611 181524 230677 181525
rect 230611 181460 230612 181524
rect 230676 181460 230677 181524
rect 230611 181459 230677 181460
rect 229875 180708 229941 180709
rect 229875 180644 229876 180708
rect 229940 180644 229941 180708
rect 229875 180643 229941 180644
rect 229139 176900 229205 176901
rect 229139 176836 229140 176900
rect 229204 176836 229205 176900
rect 229139 176835 229205 176836
rect 226195 176628 226261 176629
rect 226195 176564 226196 176628
rect 226260 176564 226261 176628
rect 226195 176563 226261 176564
rect 223619 175948 223685 175949
rect 223619 175884 223620 175948
rect 223684 175884 223685 175948
rect 223619 175883 223685 175884
rect 221207 165454 221527 165486
rect 221207 165218 221249 165454
rect 221485 165218 221527 165454
rect 221207 165134 221527 165218
rect 221207 164898 221249 165134
rect 221485 164898 221527 165134
rect 221207 164866 221527 164898
rect 224471 165454 224791 165486
rect 224471 165218 224513 165454
rect 224749 165218 224791 165454
rect 224471 165134 224791 165218
rect 224471 164898 224513 165134
rect 224749 164898 224791 165134
rect 224471 164866 224791 164898
rect 229142 149701 229202 176835
rect 229878 173909 229938 180643
rect 230427 177444 230493 177445
rect 230427 177380 230428 177444
rect 230492 177380 230493 177444
rect 230427 177379 230493 177380
rect 229875 173908 229941 173909
rect 229875 173844 229876 173908
rect 229940 173844 229941 173908
rect 229875 173843 229941 173844
rect 229139 149700 229205 149701
rect 229139 149636 229140 149700
rect 229204 149636 229205 149700
rect 229139 149635 229205 149636
rect 219575 147454 219895 147486
rect 219575 147218 219617 147454
rect 219853 147218 219895 147454
rect 219575 147134 219895 147218
rect 219575 146898 219617 147134
rect 219853 146898 219895 147134
rect 219575 146866 219895 146898
rect 222839 147454 223159 147486
rect 222839 147218 222881 147454
rect 223117 147218 223159 147454
rect 222839 147134 223159 147218
rect 222839 146898 222881 147134
rect 223117 146898 223159 147134
rect 222839 146866 223159 146898
rect 226103 147454 226423 147486
rect 226103 147218 226145 147454
rect 226381 147218 226423 147454
rect 226103 147134 226423 147218
rect 226103 146898 226145 147134
rect 226381 146898 226423 147134
rect 226103 146866 226423 146898
rect 230430 145349 230490 177379
rect 230614 176629 230674 181459
rect 231718 178397 231778 283867
rect 232454 238645 232514 354859
rect 233739 350572 233805 350573
rect 233739 350508 233740 350572
rect 233804 350508 233805 350572
rect 233739 350507 233805 350508
rect 233742 240141 233802 350507
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 457174 240134 492618
rect 239514 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 240134 457174
rect 239514 456854 240134 456938
rect 239514 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 240134 456854
rect 239514 421174 240134 456618
rect 239514 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 240134 421174
rect 239514 420854 240134 420938
rect 239514 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 240134 420854
rect 239514 385174 240134 420618
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 238523 318340 238589 318341
rect 238523 318276 238524 318340
rect 238588 318276 238589 318340
rect 238523 318275 238589 318276
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 286182 236414 308898
rect 236499 285700 236565 285701
rect 236499 285636 236500 285700
rect 236564 285636 236565 285700
rect 236499 285635 236565 285636
rect 236502 283933 236562 285635
rect 237419 284612 237485 284613
rect 237419 284548 237420 284612
rect 237484 284548 237485 284612
rect 237419 284547 237485 284548
rect 236499 283932 236565 283933
rect 236499 283868 236500 283932
rect 236564 283868 236565 283932
rect 236499 283867 236565 283868
rect 235128 255454 235448 255486
rect 235128 255218 235170 255454
rect 235406 255218 235448 255454
rect 235128 255134 235448 255218
rect 235128 254898 235170 255134
rect 235406 254898 235448 255134
rect 235128 254866 235448 254898
rect 233739 240140 233805 240141
rect 233739 240076 233740 240140
rect 233804 240076 233805 240140
rect 233739 240075 233805 240076
rect 232451 238644 232517 238645
rect 232451 238580 232452 238644
rect 232516 238580 232517 238644
rect 232451 238579 232517 238580
rect 235794 237454 236414 238182
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 231899 216748 231965 216749
rect 231899 216684 231900 216748
rect 231964 216684 231965 216748
rect 231899 216683 231965 216684
rect 231715 178396 231781 178397
rect 231715 178332 231716 178396
rect 231780 178332 231781 178396
rect 231715 178331 231781 178332
rect 230611 176628 230677 176629
rect 230611 176564 230612 176628
rect 230676 176564 230677 176628
rect 230611 176563 230677 176564
rect 231902 157453 231962 216683
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 233187 182068 233253 182069
rect 233187 182004 233188 182068
rect 233252 182004 233253 182068
rect 233187 182003 233253 182004
rect 232083 175948 232149 175949
rect 232083 175884 232084 175948
rect 232148 175884 232149 175948
rect 232083 175883 232149 175884
rect 232086 170917 232146 175883
rect 232083 170916 232149 170917
rect 232083 170852 232084 170916
rect 232148 170852 232149 170916
rect 232083 170851 232149 170852
rect 232635 157996 232701 157997
rect 232635 157932 232636 157996
rect 232700 157932 232701 157996
rect 232635 157931 232701 157932
rect 231899 157452 231965 157453
rect 231899 157388 231900 157452
rect 231964 157388 231965 157452
rect 231899 157387 231965 157388
rect 230979 152420 231045 152421
rect 230979 152356 230980 152420
rect 231044 152356 231045 152420
rect 230979 152355 231045 152356
rect 230427 145348 230493 145349
rect 230427 145284 230428 145348
rect 230492 145284 230493 145348
rect 230427 145283 230493 145284
rect 230982 131613 231042 152355
rect 231163 142764 231229 142765
rect 231163 142700 231164 142764
rect 231228 142700 231229 142764
rect 231163 142699 231229 142700
rect 230979 131612 231045 131613
rect 230979 131548 230980 131612
rect 231044 131548 231045 131612
rect 230979 131547 231045 131548
rect 221207 129454 221527 129486
rect 221207 129218 221249 129454
rect 221485 129218 221527 129454
rect 221207 129134 221527 129218
rect 221207 128898 221249 129134
rect 221485 128898 221527 129134
rect 221207 128866 221527 128898
rect 224471 129454 224791 129486
rect 224471 129218 224513 129454
rect 224749 129218 224791 129454
rect 224471 129134 224791 129218
rect 224471 128898 224513 129134
rect 224749 128898 224791 129134
rect 224471 128866 224791 128898
rect 230979 126580 231045 126581
rect 230979 126516 230980 126580
rect 231044 126516 231045 126580
rect 230979 126515 231045 126516
rect 230243 112164 230309 112165
rect 230243 112100 230244 112164
rect 230308 112100 230309 112164
rect 230243 112099 230309 112100
rect 219575 111454 219895 111486
rect 219575 111218 219617 111454
rect 219853 111218 219895 111454
rect 219575 111134 219895 111218
rect 219575 110898 219617 111134
rect 219853 110898 219895 111134
rect 219575 110866 219895 110898
rect 222839 111454 223159 111486
rect 222839 111218 222881 111454
rect 223117 111218 223159 111454
rect 222839 111134 223159 111218
rect 222839 110898 222881 111134
rect 223117 110898 223159 111134
rect 222839 110866 223159 110898
rect 226103 111454 226423 111486
rect 226103 111218 226145 111454
rect 226381 111218 226423 111454
rect 226103 111134 226423 111218
rect 226103 110898 226145 111134
rect 226381 110898 226423 111134
rect 226103 110866 226423 110898
rect 229139 96660 229205 96661
rect 229139 96596 229140 96660
rect 229204 96596 229205 96660
rect 229139 96595 229205 96596
rect 229142 96250 229202 96595
rect 228958 96190 229202 96250
rect 223619 95980 223685 95981
rect 223619 95916 223620 95980
rect 223684 95916 223685 95980
rect 223619 95915 223685 95916
rect 212395 95028 212461 95029
rect 212395 94964 212396 95028
rect 212460 94964 212461 95028
rect 212395 94963 212461 94964
rect 210954 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 211574 68614
rect 210954 68294 211574 68378
rect 210954 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 211574 68294
rect 210954 32614 211574 68058
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 75454 218414 94000
rect 217794 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 218414 75454
rect 217794 75134 218414 75218
rect 217794 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 218414 75134
rect 217794 39454 218414 74898
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 79174 222134 94000
rect 221514 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 222134 79174
rect 221514 78854 222134 78938
rect 221514 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 222134 78854
rect 221514 43174 222134 78618
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 223622 7717 223682 95915
rect 228958 95570 229018 96190
rect 228774 95510 229018 95570
rect 225234 82894 225854 94000
rect 228774 89730 228834 95510
rect 230246 95301 230306 112099
rect 230243 95300 230309 95301
rect 230243 95236 230244 95300
rect 230308 95236 230309 95300
rect 230243 95235 230309 95236
rect 225234 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 225854 82894
rect 225234 82574 225854 82658
rect 225234 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 225854 82574
rect 225234 46894 225854 82338
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 227670 89670 228834 89730
rect 227670 24173 227730 89670
rect 228954 86614 229574 94000
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 228954 50614 229574 86058
rect 230982 51781 231042 126515
rect 231166 123589 231226 142699
rect 232638 142085 232698 157931
rect 233003 151196 233069 151197
rect 233003 151132 233004 151196
rect 233068 151132 233069 151196
rect 233003 151131 233069 151132
rect 233006 142493 233066 151131
rect 233003 142492 233069 142493
rect 233003 142428 233004 142492
rect 233068 142428 233069 142492
rect 233003 142427 233069 142428
rect 232635 142084 232701 142085
rect 232635 142020 232636 142084
rect 232700 142020 232701 142084
rect 232635 142019 232701 142020
rect 232451 141132 232517 141133
rect 232451 141068 232452 141132
rect 232516 141068 232517 141132
rect 232451 141067 232517 141068
rect 231163 123588 231229 123589
rect 231163 123524 231164 123588
rect 231228 123524 231229 123588
rect 231163 123523 231229 123524
rect 232454 98021 232514 141067
rect 233190 139229 233250 182003
rect 234659 175812 234725 175813
rect 234659 175748 234660 175812
rect 234724 175748 234725 175812
rect 234659 175747 234725 175748
rect 233739 159084 233805 159085
rect 233739 159020 233740 159084
rect 233804 159020 233805 159084
rect 233739 159019 233805 159020
rect 233187 139228 233253 139229
rect 233187 139164 233188 139228
rect 233252 139164 233253 139228
rect 233187 139163 233253 139164
rect 233742 118421 233802 159019
rect 234662 137869 234722 175747
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 236502 165205 236562 283867
rect 237422 168061 237482 284547
rect 238526 240141 238586 318275
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 286182 240134 312618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 460894 243854 496338
rect 243234 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 243854 460894
rect 243234 460574 243854 460658
rect 243234 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 243854 460574
rect 243234 424894 243854 460338
rect 243234 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 243854 424894
rect 243234 424574 243854 424658
rect 243234 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 243854 424574
rect 243234 388894 243854 424338
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 464614 247574 500058
rect 246954 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 247574 464614
rect 246954 464294 247574 464378
rect 246954 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 247574 464294
rect 246954 428614 247574 464058
rect 246954 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 247574 428614
rect 246954 428294 247574 428378
rect 246954 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 247574 428294
rect 246954 392614 247574 428058
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 244227 375460 244293 375461
rect 244227 375396 244228 375460
rect 244292 375396 244293 375460
rect 244227 375395 244293 375396
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 286182 243854 316338
rect 244043 299708 244109 299709
rect 244043 299644 244044 299708
rect 244108 299644 244109 299708
rect 244043 299643 244109 299644
rect 240363 283932 240429 283933
rect 240363 283868 240364 283932
rect 240428 283868 240429 283932
rect 240363 283867 240429 283868
rect 238523 240140 238589 240141
rect 238523 240076 238524 240140
rect 238588 240076 238589 240140
rect 238523 240075 238589 240076
rect 238891 238780 238957 238781
rect 238891 238716 238892 238780
rect 238956 238716 238957 238780
rect 238891 238715 238957 238716
rect 237603 183156 237669 183157
rect 237603 183092 237604 183156
rect 237668 183092 237669 183156
rect 237603 183091 237669 183092
rect 237419 168060 237485 168061
rect 237419 167996 237420 168060
rect 237484 167996 237485 168060
rect 237419 167995 237485 167996
rect 236499 165204 236565 165205
rect 236499 165140 236500 165204
rect 236564 165140 236565 165204
rect 236499 165139 236565 165140
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 234659 137868 234725 137869
rect 234659 137804 234660 137868
rect 234724 137804 234725 137868
rect 234659 137803 234725 137804
rect 235794 129454 236414 164898
rect 237606 138821 237666 183091
rect 238894 153781 238954 238715
rect 239514 205174 240134 238182
rect 240366 234021 240426 283867
rect 244046 271010 244106 299643
rect 244230 275637 244290 375395
rect 246954 356614 247574 392058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 253794 471454 254414 506898
rect 253794 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 254414 471454
rect 253794 471134 254414 471218
rect 253794 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 254414 471134
rect 253794 435454 254414 470898
rect 253794 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 254414 435454
rect 253794 435134 254414 435218
rect 253794 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 254414 435134
rect 253794 399454 254414 434898
rect 253794 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 254414 399454
rect 253794 399134 254414 399218
rect 253794 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 254414 399134
rect 253794 363454 254414 398898
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 248459 360228 248525 360229
rect 248459 360164 248460 360228
rect 248524 360164 248525 360228
rect 248459 360163 248525 360164
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246251 304196 246317 304197
rect 246251 304132 246252 304196
rect 246316 304132 246317 304196
rect 246251 304131 246317 304132
rect 244411 282436 244477 282437
rect 244411 282372 244412 282436
rect 244476 282372 244477 282436
rect 244411 282371 244477 282372
rect 244227 275636 244293 275637
rect 244227 275572 244228 275636
rect 244292 275572 244293 275636
rect 244227 275571 244293 275572
rect 244046 270950 244290 271010
rect 244046 269109 244106 270950
rect 244230 270605 244290 270950
rect 244227 270604 244293 270605
rect 244227 270540 244228 270604
rect 244292 270540 244293 270604
rect 244227 270539 244293 270540
rect 244043 269108 244109 269109
rect 244043 269044 244044 269108
rect 244108 269044 244109 269108
rect 244043 269043 244109 269044
rect 244043 250612 244109 250613
rect 244043 250548 244044 250612
rect 244108 250548 244109 250612
rect 244043 250547 244109 250548
rect 242019 237556 242085 237557
rect 242019 237492 242020 237556
rect 242084 237492 242085 237556
rect 242019 237491 242085 237492
rect 240363 234020 240429 234021
rect 240363 233956 240364 234020
rect 240428 233956 240429 234020
rect 240363 233955 240429 233956
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 169174 240134 204618
rect 240363 199476 240429 199477
rect 240363 199412 240364 199476
rect 240428 199412 240429 199476
rect 240363 199411 240429 199412
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 238891 153780 238957 153781
rect 238891 153716 238892 153780
rect 238956 153716 238957 153780
rect 238891 153715 238957 153716
rect 237971 139772 238037 139773
rect 237971 139708 237972 139772
rect 238036 139708 238037 139772
rect 237971 139707 238037 139708
rect 237603 138820 237669 138821
rect 237603 138756 237604 138820
rect 237668 138756 237669 138820
rect 237603 138755 237669 138756
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 233739 118420 233805 118421
rect 233739 118356 233740 118420
rect 233804 118356 233805 118420
rect 233739 118355 233805 118356
rect 232451 98020 232517 98021
rect 232451 97956 232452 98020
rect 232516 97956 232517 98020
rect 232451 97955 232517 97956
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 230979 51780 231045 51781
rect 230979 51716 230980 51780
rect 231044 51716 231045 51780
rect 230979 51715 231045 51716
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 227667 24172 227733 24173
rect 227667 24108 227668 24172
rect 227732 24108 227733 24172
rect 227667 24107 227733 24108
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 223619 7716 223685 7717
rect 223619 7652 223620 7716
rect 223684 7652 223685 7716
rect 223619 7651 223685 7652
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 21454 236414 56898
rect 237974 25533 238034 139707
rect 238155 138412 238221 138413
rect 238155 138348 238156 138412
rect 238220 138348 238221 138412
rect 238155 138347 238221 138348
rect 238158 98837 238218 138347
rect 239514 133174 240134 168618
rect 240366 166973 240426 199411
rect 240731 186420 240797 186421
rect 240731 186356 240732 186420
rect 240796 186356 240797 186420
rect 240731 186355 240797 186356
rect 240363 166972 240429 166973
rect 240363 166908 240364 166972
rect 240428 166908 240429 166972
rect 240363 166907 240429 166908
rect 240734 144669 240794 186355
rect 242022 151197 242082 237491
rect 243234 208894 243854 238182
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 242939 188460 243005 188461
rect 242939 188396 242940 188460
rect 243004 188396 243005 188460
rect 242939 188395 243005 188396
rect 242019 151196 242085 151197
rect 242019 151132 242020 151196
rect 242084 151132 242085 151196
rect 242019 151131 242085 151132
rect 242019 148068 242085 148069
rect 242019 148004 242020 148068
rect 242084 148004 242085 148068
rect 242019 148003 242085 148004
rect 240731 144668 240797 144669
rect 240731 144604 240732 144668
rect 240796 144604 240797 144668
rect 240731 144603 240797 144604
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 238155 98836 238221 98837
rect 238155 98772 238156 98836
rect 238220 98772 238221 98836
rect 238155 98771 238221 98772
rect 239514 97174 240134 132618
rect 240731 119100 240797 119101
rect 240731 119036 240732 119100
rect 240796 119036 240797 119100
rect 240731 119035 240797 119036
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 237971 25532 238037 25533
rect 237971 25468 237972 25532
rect 238036 25468 238037 25532
rect 237971 25467 238037 25468
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 25174 240134 60618
rect 240734 39405 240794 119035
rect 242022 106181 242082 148003
rect 242942 136373 243002 188395
rect 243234 172894 243854 208338
rect 244046 205189 244106 250547
rect 244414 229110 244474 282371
rect 246254 273325 246314 304131
rect 246954 284614 247574 320058
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 246251 273324 246317 273325
rect 246251 273260 246252 273324
rect 246316 273260 246317 273324
rect 246251 273259 246317 273260
rect 246954 248614 247574 284058
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 245699 247348 245765 247349
rect 245699 247284 245700 247348
rect 245764 247284 245765 247348
rect 245699 247283 245765 247284
rect 245702 230349 245762 247283
rect 245883 240276 245949 240277
rect 245883 240212 245884 240276
rect 245948 240212 245949 240276
rect 245883 240211 245949 240212
rect 245699 230348 245765 230349
rect 245699 230284 245700 230348
rect 245764 230284 245765 230348
rect 245699 230283 245765 230284
rect 244230 229050 244474 229110
rect 244230 224773 244290 229050
rect 245886 227629 245946 240211
rect 245883 227628 245949 227629
rect 245883 227564 245884 227628
rect 245948 227564 245949 227628
rect 245883 227563 245949 227564
rect 244227 224772 244293 224773
rect 244227 224708 244228 224772
rect 244292 224708 244293 224772
rect 244227 224707 244293 224708
rect 244043 205188 244109 205189
rect 244043 205124 244044 205188
rect 244108 205124 244109 205188
rect 244043 205123 244109 205124
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 244230 160717 244290 224707
rect 246954 212614 247574 248058
rect 248462 242997 248522 360163
rect 252507 358868 252573 358869
rect 252507 358804 252508 358868
rect 252572 358804 252573 358868
rect 252507 358803 252573 358804
rect 249747 288692 249813 288693
rect 249747 288628 249748 288692
rect 249812 288628 249813 288692
rect 249747 288627 249813 288628
rect 248459 242996 248525 242997
rect 248459 242932 248460 242996
rect 248524 242932 248525 242996
rect 248459 242931 248525 242932
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246251 185740 246317 185741
rect 246251 185676 246252 185740
rect 246316 185676 246317 185740
rect 246251 185675 246317 185676
rect 244227 160716 244293 160717
rect 244227 160652 244228 160716
rect 244292 160652 244293 160716
rect 244227 160651 244293 160652
rect 244779 151876 244845 151877
rect 244779 151812 244780 151876
rect 244844 151812 244845 151876
rect 244779 151811 244845 151812
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 242939 136372 243005 136373
rect 242939 136308 242940 136372
rect 243004 136308 243005 136372
rect 242939 136307 243005 136308
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 242019 106180 242085 106181
rect 242019 106116 242020 106180
rect 242084 106116 242085 106180
rect 242019 106115 242085 106116
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 244782 96525 244842 151811
rect 244779 96524 244845 96525
rect 244779 96460 244780 96524
rect 244844 96460 244845 96524
rect 244779 96459 244845 96460
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 240731 39404 240797 39405
rect 240731 39340 240732 39404
rect 240796 39340 240797 39404
rect 240731 39339 240797 39340
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 246254 3501 246314 185675
rect 246954 176614 247574 212058
rect 249011 191180 249077 191181
rect 249011 191116 249012 191180
rect 249076 191116 249077 191180
rect 249011 191115 249077 191116
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 246251 3500 246317 3501
rect 246251 3436 246252 3500
rect 246316 3436 246317 3500
rect 246251 3435 246317 3436
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 249014 3501 249074 191115
rect 249750 151877 249810 288627
rect 251219 278900 251285 278901
rect 251219 278836 251220 278900
rect 251284 278836 251285 278900
rect 251219 278835 251285 278836
rect 251222 223141 251282 278835
rect 252510 235925 252570 358803
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 252507 235924 252573 235925
rect 252507 235860 252508 235924
rect 252572 235860 252573 235924
rect 252507 235859 252573 235860
rect 251219 223140 251285 223141
rect 251219 223076 251220 223140
rect 251284 223076 251285 223140
rect 251219 223075 251285 223076
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 251771 203556 251837 203557
rect 251771 203492 251772 203556
rect 251836 203492 251837 203556
rect 251771 203491 251837 203492
rect 249747 151876 249813 151877
rect 249747 151812 249748 151876
rect 249812 151812 249813 151876
rect 249747 151811 249813 151812
rect 250483 143988 250549 143989
rect 250483 143924 250484 143988
rect 250548 143924 250549 143988
rect 250483 143923 250549 143924
rect 250299 119236 250365 119237
rect 250299 119172 250300 119236
rect 250364 119172 250365 119236
rect 250299 119171 250365 119172
rect 250302 7581 250362 119171
rect 250486 111077 250546 143923
rect 250483 111076 250549 111077
rect 250483 111012 250484 111076
rect 250548 111012 250549 111076
rect 250483 111011 250549 111012
rect 250299 7580 250365 7581
rect 250299 7516 250300 7580
rect 250364 7516 250365 7580
rect 250299 7515 250365 7516
rect 251774 3637 251834 203491
rect 252507 199612 252573 199613
rect 252507 199548 252508 199612
rect 252572 199548 252573 199612
rect 252507 199547 252573 199548
rect 252510 140181 252570 199547
rect 253794 183454 254414 218898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 257514 475174 258134 510618
rect 257514 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 258134 475174
rect 257514 474854 258134 474938
rect 257514 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 258134 474854
rect 257514 439174 258134 474618
rect 257514 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 258134 439174
rect 257514 438854 258134 438938
rect 257514 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 258134 438854
rect 257514 403174 258134 438618
rect 257514 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 258134 403174
rect 257514 402854 258134 402938
rect 257514 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 258134 402854
rect 257514 367174 258134 402618
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 255819 192540 255885 192541
rect 255819 192476 255820 192540
rect 255884 192476 255885 192540
rect 255819 192475 255885 192476
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 252507 140180 252573 140181
rect 252507 140116 252508 140180
rect 252572 140116 252573 140180
rect 252507 140115 252573 140116
rect 253059 128756 253125 128757
rect 253059 128692 253060 128756
rect 253124 128692 253125 128756
rect 253059 128691 253125 128692
rect 253062 62797 253122 128691
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253059 62796 253125 62797
rect 253059 62732 253060 62796
rect 253124 62732 253125 62796
rect 253059 62731 253125 62732
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 251771 3636 251837 3637
rect 251771 3572 251772 3636
rect 251836 3572 251837 3636
rect 251771 3571 251837 3572
rect 249011 3500 249077 3501
rect 249011 3436 249012 3500
rect 249076 3436 249077 3500
rect 249011 3435 249077 3436
rect 253794 3454 254414 38898
rect 255822 3637 255882 192475
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 261234 478894 261854 514338
rect 261234 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 261854 478894
rect 261234 478574 261854 478658
rect 261234 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 261854 478574
rect 261234 442894 261854 478338
rect 261234 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 261854 442894
rect 261234 442574 261854 442658
rect 261234 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 261854 442574
rect 261234 406894 261854 442338
rect 261234 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 261854 406894
rect 261234 406574 261854 406658
rect 261234 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 261854 406574
rect 261234 370894 261854 406338
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 260051 134604 260117 134605
rect 260051 134540 260052 134604
rect 260116 134540 260117 134604
rect 260051 134539 260117 134540
rect 258579 127124 258645 127125
rect 258579 127060 258580 127124
rect 258644 127060 258645 127124
rect 258579 127059 258645 127060
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 258582 66877 258642 127059
rect 260054 102781 260114 134539
rect 261234 118894 261854 154338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 264954 482614 265574 518058
rect 264954 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 265574 482614
rect 264954 482294 265574 482378
rect 264954 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 265574 482294
rect 264954 446614 265574 482058
rect 264954 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 265574 446614
rect 264954 446294 265574 446378
rect 264954 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 265574 446294
rect 264954 410614 265574 446058
rect 264954 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 265574 410614
rect 264954 410294 265574 410378
rect 264954 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 265574 410294
rect 264954 374614 265574 410058
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271794 453454 272414 488898
rect 271794 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 272414 453454
rect 271794 453134 272414 453218
rect 271794 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 272414 453134
rect 271794 417454 272414 452898
rect 271794 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 272414 417454
rect 271794 417134 272414 417218
rect 271794 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 272414 417134
rect 271794 381454 272414 416898
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 457174 276134 492618
rect 275514 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 276134 457174
rect 275514 456854 276134 456938
rect 275514 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 276134 456854
rect 275514 421174 276134 456618
rect 275514 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 276134 421174
rect 275514 420854 276134 420938
rect 275514 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 276134 420854
rect 275514 385174 276134 420618
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 274587 272236 274653 272237
rect 274587 272172 274588 272236
rect 274652 272172 274653 272236
rect 274587 272171 274653 272172
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 178000 272414 200898
rect 274590 179077 274650 272171
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 274587 179076 274653 179077
rect 274587 179012 274588 179076
rect 274652 179012 274653 179076
rect 274587 179011 274653 179012
rect 275514 178000 276134 204618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 279234 460894 279854 496338
rect 279234 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 279854 460894
rect 279234 460574 279854 460658
rect 279234 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 279854 460574
rect 279234 424894 279854 460338
rect 279234 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 279854 424894
rect 279234 424574 279854 424658
rect 279234 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 279854 424574
rect 279234 388894 279854 424338
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 464614 283574 500058
rect 282954 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 283574 464614
rect 282954 464294 283574 464378
rect 282954 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 283574 464294
rect 282954 428614 283574 464058
rect 282954 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 283574 428614
rect 282954 428294 283574 428378
rect 282954 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 283574 428294
rect 282954 392614 283574 428058
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 289794 471454 290414 506898
rect 289794 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 290414 471454
rect 289794 471134 290414 471218
rect 289794 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 290414 471134
rect 289794 435454 290414 470898
rect 289794 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 290414 435454
rect 289794 435134 290414 435218
rect 289794 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 290414 435134
rect 289794 399454 290414 434898
rect 289794 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 290414 399454
rect 289794 399134 290414 399218
rect 289794 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 290414 399134
rect 289794 363454 290414 398898
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 475174 294134 510618
rect 293514 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 294134 475174
rect 293514 474854 294134 474938
rect 293514 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 294134 474854
rect 293514 439174 294134 474618
rect 293514 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 294134 439174
rect 293514 438854 294134 438938
rect 293514 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 294134 438854
rect 293514 403174 294134 438618
rect 293514 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 294134 403174
rect 293514 402854 294134 402938
rect 293514 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 294134 402854
rect 293514 367174 294134 402618
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 291147 339556 291213 339557
rect 291147 339492 291148 339556
rect 291212 339492 291213 339556
rect 291147 339491 291213 339492
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 285627 288556 285693 288557
rect 285627 288492 285628 288556
rect 285692 288492 285693 288556
rect 285627 288491 285693 288492
rect 284339 287604 284405 287605
rect 284339 287540 284340 287604
rect 284404 287540 284405 287604
rect 284339 287539 284405 287540
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 280291 219468 280357 219469
rect 280291 219404 280292 219468
rect 280356 219404 280357 219468
rect 280291 219403 280357 219404
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 278819 178668 278885 178669
rect 278819 178604 278820 178668
rect 278884 178604 278885 178668
rect 278819 178603 278885 178604
rect 278822 167650 278882 178603
rect 279234 178000 279854 208338
rect 280294 190470 280354 219403
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 280475 192676 280541 192677
rect 280475 192612 280476 192676
rect 280540 192612 280541 192676
rect 280475 192611 280541 192612
rect 280110 190410 280354 190470
rect 279371 177036 279437 177037
rect 279371 176972 279372 177036
rect 279436 176972 279437 177036
rect 279371 176971 279437 176972
rect 279374 173773 279434 176971
rect 279371 173772 279437 173773
rect 279371 173708 279372 173772
rect 279436 173708 279437 173772
rect 279371 173707 279437 173708
rect 279371 167652 279437 167653
rect 279371 167650 279372 167652
rect 278822 167590 279372 167650
rect 279371 167588 279372 167590
rect 279436 167588 279437 167652
rect 279371 167587 279437 167588
rect 272207 165454 272527 165486
rect 272207 165218 272249 165454
rect 272485 165218 272527 165454
rect 272207 165134 272527 165218
rect 272207 164898 272249 165134
rect 272485 164898 272527 165134
rect 272207 164866 272527 164898
rect 275471 165454 275791 165486
rect 275471 165218 275513 165454
rect 275749 165218 275791 165454
rect 275471 165134 275791 165218
rect 275471 164898 275513 165134
rect 275749 164898 275791 165134
rect 275471 164866 275791 164898
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 262811 131068 262877 131069
rect 262811 131004 262812 131068
rect 262876 131004 262877 131068
rect 262811 131003 262877 131004
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 260051 102780 260117 102781
rect 260051 102716 260052 102780
rect 260116 102716 260117 102780
rect 260051 102715 260117 102716
rect 260051 99788 260117 99789
rect 260051 99724 260052 99788
rect 260116 99724 260117 99788
rect 260051 99723 260117 99724
rect 258579 66876 258645 66877
rect 258579 66812 258580 66876
rect 258644 66812 258645 66876
rect 258579 66811 258645 66812
rect 260054 55861 260114 99723
rect 261234 82894 261854 118338
rect 262075 114612 262141 114613
rect 262075 114548 262076 114612
rect 262140 114548 262141 114612
rect 262075 114547 262141 114548
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 260051 55860 260117 55861
rect 260051 55796 260052 55860
rect 260116 55796 260117 55860
rect 260051 55795 260117 55796
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 255819 3636 255885 3637
rect 255819 3572 255820 3636
rect 255884 3572 255885 3636
rect 255819 3571 255885 3572
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 262078 21317 262138 114547
rect 262814 72589 262874 131003
rect 264099 127940 264165 127941
rect 264099 127876 264100 127940
rect 264164 127876 264165 127940
rect 264099 127875 264165 127876
rect 262995 100468 263061 100469
rect 262995 100404 262996 100468
rect 263060 100404 263061 100468
rect 262995 100403 263061 100404
rect 262998 98837 263058 100403
rect 263179 99244 263245 99245
rect 263179 99180 263180 99244
rect 263244 99180 263245 99244
rect 263179 99179 263245 99180
rect 262995 98836 263061 98837
rect 262995 98772 262996 98836
rect 263060 98772 263061 98836
rect 262995 98771 263061 98772
rect 263182 96389 263242 99179
rect 263179 96388 263245 96389
rect 263179 96324 263180 96388
rect 263244 96324 263245 96388
rect 263179 96323 263245 96324
rect 262811 72588 262877 72589
rect 262811 72524 262812 72588
rect 262876 72524 262877 72588
rect 262811 72523 262877 72524
rect 264102 39269 264162 127875
rect 264954 122614 265574 158058
rect 270575 147454 270895 147486
rect 270575 147218 270617 147454
rect 270853 147218 270895 147454
rect 270575 147134 270895 147218
rect 270575 146898 270617 147134
rect 270853 146898 270895 147134
rect 270575 146866 270895 146898
rect 273839 147454 274159 147486
rect 273839 147218 273881 147454
rect 274117 147218 274159 147454
rect 273839 147134 274159 147218
rect 273839 146898 273881 147134
rect 274117 146898 274159 147134
rect 273839 146866 274159 146898
rect 277103 147454 277423 147486
rect 277103 147218 277145 147454
rect 277381 147218 277423 147454
rect 277103 147134 277423 147218
rect 277103 146898 277145 147134
rect 277381 146898 277423 147134
rect 277103 146866 277423 146898
rect 272207 129454 272527 129486
rect 266859 129300 266925 129301
rect 266859 129236 266860 129300
rect 266924 129236 266925 129300
rect 266859 129235 266925 129236
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264099 39268 264165 39269
rect 264099 39204 264100 39268
rect 264164 39204 264165 39268
rect 264099 39203 264165 39204
rect 262075 21316 262141 21317
rect 262075 21252 262076 21316
rect 262140 21252 262141 21316
rect 262075 21251 262141 21252
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 14614 265574 50058
rect 266862 48925 266922 129235
rect 272207 129218 272249 129454
rect 272485 129218 272527 129454
rect 272207 129134 272527 129218
rect 272207 128898 272249 129134
rect 272485 128898 272527 129134
rect 272207 128866 272527 128898
rect 275471 129454 275791 129486
rect 275471 129218 275513 129454
rect 275749 129218 275791 129454
rect 275471 129134 275791 129218
rect 275471 128898 275513 129134
rect 275749 128898 275791 129134
rect 275471 128866 275791 128898
rect 267779 128484 267845 128485
rect 267779 128420 267780 128484
rect 267844 128420 267845 128484
rect 267779 128419 267845 128420
rect 266859 48924 266925 48925
rect 266859 48860 266860 48924
rect 266924 48860 266925 48924
rect 266859 48859 266925 48860
rect 267782 26893 267842 128419
rect 280110 126853 280170 190410
rect 280478 180810 280538 192611
rect 281579 181524 281645 181525
rect 281579 181460 281580 181524
rect 281644 181460 281645 181524
rect 281579 181459 281645 181460
rect 280294 180750 280538 180810
rect 280294 151830 280354 180750
rect 281582 170917 281642 181459
rect 282954 176614 283574 212058
rect 283787 194036 283853 194037
rect 283787 193972 283788 194036
rect 283852 193972 283853 194036
rect 283787 193971 283853 193972
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 281579 170916 281645 170917
rect 281579 170852 281580 170916
rect 281644 170852 281645 170916
rect 281579 170851 281645 170852
rect 280294 151770 280538 151830
rect 280107 126852 280173 126853
rect 280107 126788 280108 126852
rect 280172 126788 280173 126852
rect 280107 126787 280173 126788
rect 280478 122850 280538 151770
rect 280294 122790 280538 122850
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 280294 120733 280354 122790
rect 280291 120732 280357 120733
rect 280291 120668 280292 120732
rect 280356 120668 280357 120732
rect 280291 120667 280357 120668
rect 270575 111454 270895 111486
rect 270575 111218 270617 111454
rect 270853 111218 270895 111454
rect 270575 111134 270895 111218
rect 270575 110898 270617 111134
rect 270853 110898 270895 111134
rect 270575 110866 270895 110898
rect 273839 111454 274159 111486
rect 273839 111218 273881 111454
rect 274117 111218 274159 111454
rect 273839 111134 274159 111218
rect 273839 110898 273881 111134
rect 274117 110898 274159 111134
rect 273839 110866 274159 110898
rect 277103 111454 277423 111486
rect 277103 111218 277145 111454
rect 277381 111218 277423 111454
rect 277103 111134 277423 111218
rect 277103 110898 277145 111134
rect 277381 110898 277423 111134
rect 277103 110866 277423 110898
rect 282954 104614 283574 140058
rect 283790 135149 283850 193971
rect 283787 135148 283853 135149
rect 283787 135084 283788 135148
rect 283852 135084 283853 135148
rect 283787 135083 283853 135084
rect 284342 111621 284402 287539
rect 284523 183020 284589 183021
rect 284523 182956 284524 183020
rect 284588 182956 284589 183020
rect 284523 182955 284589 182956
rect 284526 167925 284586 182955
rect 284523 167924 284589 167925
rect 284523 167860 284524 167924
rect 284588 167860 284589 167924
rect 284523 167859 284589 167860
rect 284339 111620 284405 111621
rect 284339 111556 284340 111620
rect 284404 111556 284405 111620
rect 284339 111555 284405 111556
rect 285630 106997 285690 288491
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 288387 200836 288453 200837
rect 288387 200772 288388 200836
rect 288452 200772 288453 200836
rect 288387 200771 288453 200772
rect 287099 193900 287165 193901
rect 287099 193836 287100 193900
rect 287164 193836 287165 193900
rect 287099 193835 287165 193836
rect 285811 182884 285877 182885
rect 285811 182820 285812 182884
rect 285876 182820 285877 182884
rect 285811 182819 285877 182820
rect 285627 106996 285693 106997
rect 285627 106932 285628 106996
rect 285692 106932 285693 106996
rect 285627 106931 285693 106932
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 268515 97612 268581 97613
rect 268515 97548 268516 97612
rect 268580 97548 268581 97612
rect 268515 97547 268581 97548
rect 268518 94893 268578 97547
rect 268515 94892 268581 94893
rect 268515 94828 268516 94892
rect 268580 94828 268581 94892
rect 268515 94827 268581 94828
rect 271794 93454 272414 94000
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 267779 26892 267845 26893
rect 267779 26828 267780 26892
rect 267844 26828 267845 26892
rect 267779 26827 267845 26828
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 61174 276134 94000
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 64894 279854 94000
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 285814 3501 285874 182819
rect 287102 3501 287162 193835
rect 287283 177444 287349 177445
rect 287283 177380 287284 177444
rect 287348 177380 287349 177444
rect 287283 177379 287349 177380
rect 287286 149157 287346 177379
rect 287283 149156 287349 149157
rect 287283 149092 287284 149156
rect 287348 149092 287349 149156
rect 287283 149091 287349 149092
rect 288390 3501 288450 200771
rect 288571 184244 288637 184245
rect 288571 184180 288572 184244
rect 288636 184180 288637 184244
rect 288571 184179 288637 184180
rect 288574 104957 288634 184179
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 288571 104956 288637 104957
rect 288571 104892 288572 104956
rect 288636 104892 288637 104956
rect 288571 104891 288637 104892
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 285811 3500 285877 3501
rect 285811 3436 285812 3500
rect 285876 3436 285877 3500
rect 285811 3435 285877 3436
rect 287099 3500 287165 3501
rect 287099 3436 287100 3500
rect 287164 3436 287165 3500
rect 287099 3435 287165 3436
rect 288387 3500 288453 3501
rect 288387 3436 288388 3500
rect 288452 3436 288453 3500
rect 288387 3435 288453 3436
rect 289794 3454 290414 38898
rect 291150 3501 291210 339491
rect 293514 331174 294134 366618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 478894 297854 514338
rect 297234 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 297854 478894
rect 297234 478574 297854 478658
rect 297234 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 297854 478574
rect 297234 442894 297854 478338
rect 297234 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 297854 442894
rect 297234 442574 297854 442658
rect 297234 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 297854 442574
rect 297234 406894 297854 442338
rect 297234 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 297854 406894
rect 297234 406574 297854 406658
rect 297234 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 297854 406574
rect 297234 370894 297854 406338
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 295931 334116 295997 334117
rect 295931 334052 295932 334116
rect 295996 334052 295997 334116
rect 295931 334051 295997 334052
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 291331 185740 291397 185741
rect 291331 185676 291332 185740
rect 291396 185676 291397 185740
rect 291331 185675 291397 185676
rect 291334 156093 291394 185675
rect 291331 156092 291397 156093
rect 291331 156028 291332 156092
rect 291396 156028 291397 156092
rect 291331 156027 291397 156028
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 291147 3500 291213 3501
rect 291147 3436 291148 3500
rect 291212 3436 291213 3500
rect 291147 3435 291213 3436
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 -2266 294134 6618
rect 295934 4045 295994 334051
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 482614 301574 518058
rect 300954 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 301574 482614
rect 300954 482294 301574 482378
rect 300954 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 301574 482294
rect 300954 446614 301574 482058
rect 300954 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 301574 446614
rect 300954 446294 301574 446378
rect 300954 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 301574 446294
rect 300954 410614 301574 446058
rect 300954 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 301574 410614
rect 300954 410294 301574 410378
rect 300954 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 301574 410294
rect 300954 374614 301574 410058
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 453454 308414 488898
rect 307794 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 308414 453454
rect 307794 453134 308414 453218
rect 307794 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 308414 453134
rect 307794 417454 308414 452898
rect 307794 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 308414 417454
rect 307794 417134 308414 417218
rect 307794 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 308414 417134
rect 307794 381454 308414 416898
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 302739 309228 302805 309229
rect 302739 309164 302740 309228
rect 302804 309164 302805 309228
rect 302739 309163 302805 309164
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 299611 214572 299677 214573
rect 299611 214508 299612 214572
rect 299676 214508 299677 214572
rect 299611 214507 299677 214508
rect 298139 206276 298205 206277
rect 298139 206212 298140 206276
rect 298204 206212 298205 206276
rect 298139 206211 298205 206212
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 295931 4044 295997 4045
rect 295931 3980 295932 4044
rect 295996 3980 295997 4044
rect 295931 3979 295997 3980
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 -4186 297854 10338
rect 298142 3909 298202 206211
rect 298139 3908 298205 3909
rect 298139 3844 298140 3908
rect 298204 3844 298205 3908
rect 298139 3843 298205 3844
rect 299614 3501 299674 214507
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 299611 3500 299677 3501
rect 299611 3436 299612 3500
rect 299676 3436 299677 3500
rect 299611 3435 299677 3436
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 302742 4861 302802 309163
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 302739 4860 302805 4861
rect 302739 4796 302740 4860
rect 302804 4796 302805 4860
rect 302739 4795 302805 4796
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 457174 312134 492618
rect 311514 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 312134 457174
rect 311514 456854 312134 456938
rect 311514 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 312134 456854
rect 311514 421174 312134 456618
rect 311514 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 312134 421174
rect 311514 420854 312134 420938
rect 311514 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 312134 420854
rect 311514 385174 312134 420618
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 315234 460894 315854 496338
rect 315234 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 315854 460894
rect 315234 460574 315854 460658
rect 315234 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 315854 460574
rect 315234 424894 315854 460338
rect 315234 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 315854 424894
rect 315234 424574 315854 424658
rect 315234 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 315854 424574
rect 315234 388894 315854 424338
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318954 464614 319574 500058
rect 318954 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 319574 464614
rect 318954 464294 319574 464378
rect 318954 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 319574 464294
rect 318954 428614 319574 464058
rect 318954 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 319574 428614
rect 318954 428294 319574 428378
rect 318954 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 319574 428294
rect 318954 392614 319574 428058
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 325794 471454 326414 506898
rect 325794 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 326414 471454
rect 325794 471134 326414 471218
rect 325794 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 326414 471134
rect 325794 435454 326414 470898
rect 325794 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 326414 435454
rect 325794 435134 326414 435218
rect 325794 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 326414 435134
rect 325794 399454 326414 434898
rect 325794 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 326414 399454
rect 325794 399134 326414 399218
rect 325794 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 326414 399134
rect 325794 363454 326414 398898
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 475174 330134 510618
rect 329514 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 330134 475174
rect 329514 474854 330134 474938
rect 329514 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 330134 474854
rect 329514 439174 330134 474618
rect 329514 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 330134 439174
rect 329514 438854 330134 438938
rect 329514 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 330134 438854
rect 329514 403174 330134 438618
rect 329514 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 330134 403174
rect 329514 402854 330134 402938
rect 329514 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 330134 402854
rect 329514 367174 330134 402618
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 478894 333854 514338
rect 333234 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 333854 478894
rect 333234 478574 333854 478658
rect 333234 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 333854 478574
rect 333234 442894 333854 478338
rect 333234 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 333854 442894
rect 333234 442574 333854 442658
rect 333234 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 333854 442574
rect 333234 406894 333854 442338
rect 333234 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 333854 406894
rect 333234 406574 333854 406658
rect 333234 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 333854 406574
rect 333234 370894 333854 406338
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 482614 337574 518058
rect 336954 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 337574 482614
rect 336954 482294 337574 482378
rect 336954 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 337574 482294
rect 336954 446614 337574 482058
rect 336954 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 337574 446614
rect 336954 446294 337574 446378
rect 336954 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 337574 446294
rect 336954 410614 337574 446058
rect 336954 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 337574 410614
rect 336954 410294 337574 410378
rect 336954 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 337574 410294
rect 336954 374614 337574 410058
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 343794 453454 344414 488898
rect 343794 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 344414 453454
rect 343794 453134 344414 453218
rect 343794 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 344414 453134
rect 343794 417454 344414 452898
rect 343794 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 344414 417454
rect 343794 417134 344414 417218
rect 343794 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 344414 417134
rect 343794 381454 344414 416898
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 457174 348134 492618
rect 347514 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 348134 457174
rect 347514 456854 348134 456938
rect 347514 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 348134 456854
rect 347514 421174 348134 456618
rect 347514 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 348134 421174
rect 347514 420854 348134 420938
rect 347514 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 348134 420854
rect 347514 385174 348134 420618
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 351234 460894 351854 496338
rect 351234 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 351854 460894
rect 351234 460574 351854 460658
rect 351234 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 351854 460574
rect 351234 424894 351854 460338
rect 351234 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 351854 424894
rect 351234 424574 351854 424658
rect 351234 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 351854 424574
rect 351234 388894 351854 424338
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 464614 355574 500058
rect 354954 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 355574 464614
rect 354954 464294 355574 464378
rect 354954 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 355574 464294
rect 354954 428614 355574 464058
rect 354954 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 355574 428614
rect 354954 428294 355574 428378
rect 354954 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 355574 428294
rect 354954 392614 355574 428058
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 59546 456938 59782 457174
rect 59866 456938 60102 457174
rect 59546 456618 59782 456854
rect 59866 456618 60102 456854
rect 59546 420938 59782 421174
rect 59866 420938 60102 421174
rect 59546 420618 59782 420854
rect 59866 420618 60102 420854
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 59546 204938 59782 205174
rect 59866 204938 60102 205174
rect 59546 204618 59782 204854
rect 59866 204618 60102 204854
rect 59546 168938 59782 169174
rect 59866 168938 60102 169174
rect 59546 168618 59782 168854
rect 59866 168618 60102 168854
rect 59546 132938 59782 133174
rect 59866 132938 60102 133174
rect 59546 132618 59782 132854
rect 59866 132618 60102 132854
rect 59546 96938 59782 97174
rect 59866 96938 60102 97174
rect 59546 96618 59782 96854
rect 59866 96618 60102 96854
rect 59546 60938 59782 61174
rect 59866 60938 60102 61174
rect 59546 60618 59782 60854
rect 59866 60618 60102 60854
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 72721 579218 72957 579454
rect 72721 578898 72957 579134
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 63266 460658 63502 460894
rect 63586 460658 63822 460894
rect 63266 460338 63502 460574
rect 63586 460338 63822 460574
rect 63266 424658 63502 424894
rect 63586 424658 63822 424894
rect 63266 424338 63502 424574
rect 63586 424338 63822 424574
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 75686 561218 75922 561454
rect 75686 560898 75922 561134
rect 72721 543218 72957 543454
rect 72721 542898 72957 543134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 78651 579218 78887 579454
rect 78651 578898 78887 579134
rect 84582 579218 84818 579454
rect 84582 578898 84818 579134
rect 81617 561218 81853 561454
rect 81617 560898 81853 561134
rect 78651 543218 78887 543454
rect 78651 542898 78887 543134
rect 84582 543218 84818 543454
rect 84582 542898 84818 543134
rect 66986 464378 67222 464614
rect 67306 464378 67542 464614
rect 66986 464058 67222 464294
rect 67306 464058 67542 464294
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 63266 208658 63502 208894
rect 63586 208658 63822 208894
rect 63266 208338 63502 208574
rect 63586 208338 63822 208574
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 73826 471218 74062 471454
rect 74146 471218 74382 471454
rect 73826 470898 74062 471134
rect 74146 470898 74382 471134
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 77546 474938 77782 475174
rect 77866 474938 78102 475174
rect 77546 474618 77782 474854
rect 77866 474618 78102 474854
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 81266 478658 81502 478894
rect 81586 478658 81822 478894
rect 81266 478338 81502 478574
rect 81586 478338 81822 478574
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 84986 482378 85222 482614
rect 85306 482378 85542 482614
rect 84986 482058 85222 482294
rect 85306 482058 85542 482294
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 73020 435218 73256 435454
rect 73020 434898 73256 435134
rect 88380 417218 88616 417454
rect 88380 416898 88616 417134
rect 73020 399218 73256 399454
rect 73020 398898 73256 399134
rect 63266 172658 63502 172894
rect 63586 172658 63822 172894
rect 63266 172338 63502 172574
rect 63586 172338 63822 172574
rect 63266 136658 63502 136894
rect 63586 136658 63822 136894
rect 63266 136338 63502 136574
rect 63586 136338 63822 136574
rect 63266 100658 63502 100894
rect 63586 100658 63822 100894
rect 63266 100338 63502 100574
rect 63586 100338 63822 100574
rect 63266 64658 63502 64894
rect 63586 64658 63822 64894
rect 63266 64338 63502 64574
rect 63586 64338 63822 64574
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 66986 212378 67222 212614
rect 67306 212378 67542 212614
rect 66986 212058 67222 212294
rect 67306 212058 67542 212294
rect 66986 68378 67222 68614
rect 67306 68378 67542 68614
rect 66986 68058 67222 68294
rect 67306 68058 67542 68294
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 91826 453218 92062 453454
rect 92146 453218 92382 453454
rect 91826 452898 92062 453134
rect 92146 452898 92382 453134
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 95546 456938 95782 457174
rect 95866 456938 96102 457174
rect 95546 456618 95782 456854
rect 95866 456618 96102 456854
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 99266 460658 99502 460894
rect 99586 460658 99822 460894
rect 99266 460338 99502 460574
rect 99586 460338 99822 460574
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 109826 471218 110062 471454
rect 110146 471218 110382 471454
rect 109826 470898 110062 471134
rect 110146 470898 110382 471134
rect 102986 464378 103222 464614
rect 103306 464378 103542 464614
rect 102986 464058 103222 464294
rect 103306 464058 103542 464294
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 103740 435218 103976 435454
rect 103740 434898 103976 435134
rect 103740 399218 103976 399454
rect 103740 398898 103976 399134
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 113546 474938 113782 475174
rect 113866 474938 114102 475174
rect 113546 474618 113782 474854
rect 113866 474618 114102 474854
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 117266 478658 117502 478894
rect 117586 478658 117822 478894
rect 117266 478338 117502 478574
rect 117586 478338 117822 478574
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 120986 482378 121222 482614
rect 121306 482378 121542 482614
rect 120986 482058 121222 482294
rect 121306 482058 121542 482294
rect 119100 417218 119336 417454
rect 119100 416898 119336 417134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 127826 453218 128062 453454
rect 128146 453218 128382 453454
rect 127826 452898 128062 453134
rect 128146 452898 128382 453134
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 127826 417218 128062 417454
rect 128146 417218 128382 417454
rect 127826 416898 128062 417134
rect 128146 416898 128382 417134
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 131546 456938 131782 457174
rect 131866 456938 132102 457174
rect 131546 456618 131782 456854
rect 131866 456618 132102 456854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 135266 460658 135502 460894
rect 135586 460658 135822 460894
rect 135266 460338 135502 460574
rect 135586 460338 135822 460574
rect 131546 420938 131782 421174
rect 131866 420938 132102 421174
rect 131546 420618 131782 420854
rect 131866 420618 132102 420854
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 73020 291218 73256 291454
rect 73020 290898 73256 291134
rect 73020 255218 73256 255454
rect 73020 254898 73256 255134
rect 73826 219218 74062 219454
rect 74146 219218 74382 219454
rect 73826 218898 74062 219134
rect 74146 218898 74382 219134
rect 73826 183218 74062 183454
rect 74146 183218 74382 183454
rect 73826 182898 74062 183134
rect 74146 182898 74382 183134
rect 77546 222938 77782 223174
rect 77866 222938 78102 223174
rect 77546 222618 77782 222854
rect 77866 222618 78102 222854
rect 77546 186938 77782 187174
rect 77866 186938 78102 187174
rect 77546 186618 77782 186854
rect 77866 186618 78102 186854
rect 81266 226658 81502 226894
rect 81586 226658 81822 226894
rect 81266 226338 81502 226574
rect 81586 226338 81822 226574
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 81266 190658 81502 190894
rect 81586 190658 81822 190894
rect 81266 190338 81502 190574
rect 81586 190338 81822 190574
rect 88380 309218 88616 309454
rect 88380 308898 88616 309134
rect 119100 309218 119336 309454
rect 119100 308898 119336 309134
rect 103740 291218 103976 291454
rect 103740 290898 103976 291134
rect 88380 273218 88616 273454
rect 88380 272898 88616 273134
rect 119100 273218 119336 273454
rect 119100 272898 119336 273134
rect 103740 255218 103976 255454
rect 103740 254898 103976 255134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 84986 194378 85222 194614
rect 85306 194378 85542 194614
rect 84986 194058 85222 194294
rect 85306 194058 85542 194294
rect 91826 201218 92062 201454
rect 92146 201218 92382 201454
rect 91826 200898 92062 201134
rect 92146 200898 92382 201134
rect 95546 204938 95782 205174
rect 95866 204938 96102 205174
rect 95546 204618 95782 204854
rect 95866 204618 96102 204854
rect 99266 208658 99502 208894
rect 99586 208658 99822 208894
rect 99266 208338 99502 208574
rect 99586 208338 99822 208574
rect 102986 212378 103222 212614
rect 103306 212378 103542 212614
rect 102986 212058 103222 212294
rect 103306 212058 103542 212294
rect 109826 219218 110062 219454
rect 110146 219218 110382 219454
rect 109826 218898 110062 219134
rect 110146 218898 110382 219134
rect 109826 183218 110062 183454
rect 110146 183218 110382 183454
rect 109826 182898 110062 183134
rect 110146 182898 110382 183134
rect 113546 222938 113782 223174
rect 113866 222938 114102 223174
rect 113546 222618 113782 222854
rect 113866 222618 114102 222854
rect 113546 186938 113782 187174
rect 113866 186938 114102 187174
rect 113546 186618 113782 186854
rect 113866 186618 114102 186854
rect 117266 226658 117502 226894
rect 117586 226658 117822 226894
rect 117266 226338 117502 226574
rect 117586 226338 117822 226574
rect 117266 190658 117502 190894
rect 117586 190658 117822 190894
rect 117266 190338 117502 190574
rect 117586 190338 117822 190574
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 120986 194378 121222 194614
rect 121306 194378 121542 194614
rect 120986 194058 121222 194294
rect 121306 194058 121542 194294
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 127826 201218 128062 201454
rect 128146 201218 128382 201454
rect 127826 200898 128062 201134
rect 128146 200898 128382 201134
rect 135266 424658 135502 424894
rect 135586 424658 135822 424894
rect 135266 424338 135502 424574
rect 135586 424338 135822 424574
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 138986 464378 139222 464614
rect 139306 464378 139542 464614
rect 138986 464058 139222 464294
rect 139306 464058 139542 464294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 145826 471218 146062 471454
rect 146146 471218 146382 471454
rect 145826 470898 146062 471134
rect 146146 470898 146382 471134
rect 138986 428378 139222 428614
rect 139306 428378 139542 428614
rect 138986 428058 139222 428294
rect 139306 428058 139542 428294
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 134460 291218 134696 291454
rect 134460 290898 134696 291134
rect 134460 255218 134696 255454
rect 134460 254898 134696 255134
rect 131546 204938 131782 205174
rect 131866 204938 132102 205174
rect 131546 204618 131782 204854
rect 131866 204618 132102 204854
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 135266 208658 135502 208894
rect 135586 208658 135822 208894
rect 135266 208338 135502 208574
rect 135586 208338 135822 208574
rect 145826 435218 146062 435454
rect 146146 435218 146382 435454
rect 145826 434898 146062 435134
rect 146146 434898 146382 435134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 149546 474938 149782 475174
rect 149866 474938 150102 475174
rect 149546 474618 149782 474854
rect 149866 474618 150102 474854
rect 149546 438938 149782 439174
rect 149866 438938 150102 439174
rect 149546 438618 149782 438854
rect 149866 438618 150102 438854
rect 145826 399218 146062 399454
rect 146146 399218 146382 399454
rect 145826 398898 146062 399134
rect 146146 398898 146382 399134
rect 149546 402938 149782 403174
rect 149866 402938 150102 403174
rect 149546 402618 149782 402854
rect 149866 402618 150102 402854
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 138986 212378 139222 212614
rect 139306 212378 139542 212614
rect 138986 212058 139222 212294
rect 139306 212058 139542 212294
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 153266 478658 153502 478894
rect 153586 478658 153822 478894
rect 153266 478338 153502 478574
rect 153586 478338 153822 478574
rect 153266 442658 153502 442894
rect 153586 442658 153822 442894
rect 153266 442338 153502 442574
rect 153586 442338 153822 442574
rect 153266 406658 153502 406894
rect 153586 406658 153822 406894
rect 153266 406338 153502 406574
rect 153586 406338 153822 406574
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149820 309218 150056 309454
rect 149820 308898 150056 309134
rect 149820 273218 150056 273454
rect 149820 272898 150056 273134
rect 145826 219218 146062 219454
rect 146146 219218 146382 219454
rect 145826 218898 146062 219134
rect 146146 218898 146382 219134
rect 145826 183218 146062 183454
rect 146146 183218 146382 183454
rect 145826 182898 146062 183134
rect 146146 182898 146382 183134
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 156986 482378 157222 482614
rect 157306 482378 157542 482614
rect 156986 482058 157222 482294
rect 157306 482058 157542 482294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 163826 453218 164062 453454
rect 164146 453218 164382 453454
rect 163826 452898 164062 453134
rect 164146 452898 164382 453134
rect 156986 446378 157222 446614
rect 157306 446378 157542 446614
rect 156986 446058 157222 446294
rect 157306 446058 157542 446294
rect 156986 410378 157222 410614
rect 157306 410378 157542 410614
rect 156986 410058 157222 410294
rect 157306 410058 157542 410294
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 163826 417218 164062 417454
rect 164146 417218 164382 417454
rect 163826 416898 164062 417134
rect 164146 416898 164382 417134
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 167546 456938 167782 457174
rect 167866 456938 168102 457174
rect 167546 456618 167782 456854
rect 167866 456618 168102 456854
rect 167546 420938 167782 421174
rect 167866 420938 168102 421174
rect 167546 420618 167782 420854
rect 167866 420618 168102 420854
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 153266 226658 153502 226894
rect 153586 226658 153822 226894
rect 153266 226338 153502 226574
rect 153586 226338 153822 226574
rect 149546 222938 149782 223174
rect 149866 222938 150102 223174
rect 149546 222618 149782 222854
rect 149866 222618 150102 222854
rect 149546 186938 149782 187174
rect 149866 186938 150102 187174
rect 149546 186618 149782 186854
rect 149866 186618 150102 186854
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 153266 190658 153502 190894
rect 153586 190658 153822 190894
rect 153266 190338 153502 190574
rect 153586 190338 153822 190574
rect 156986 194378 157222 194614
rect 157306 194378 157542 194614
rect 156986 194058 157222 194294
rect 157306 194058 157542 194294
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 163826 201218 164062 201454
rect 164146 201218 164382 201454
rect 163826 200898 164062 201134
rect 164146 200898 164382 201134
rect 69128 165218 69364 165454
rect 69128 164898 69364 165134
rect 164192 165218 164428 165454
rect 164192 164898 164428 165134
rect 69808 147218 70044 147454
rect 69808 146898 70044 147134
rect 163512 147218 163748 147454
rect 163512 146898 163748 147134
rect 69128 129218 69364 129454
rect 69128 128898 69364 129134
rect 164192 129218 164428 129454
rect 164192 128898 164428 129134
rect 69808 111218 70044 111454
rect 69808 110898 70044 111134
rect 163512 111218 163748 111454
rect 163512 110898 163748 111134
rect 73826 75218 74062 75454
rect 74146 75218 74382 75454
rect 73826 74898 74062 75134
rect 74146 74898 74382 75134
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 78938 77782 79174
rect 77866 78938 78102 79174
rect 77546 78618 77782 78854
rect 77866 78618 78102 78854
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 82658 81502 82894
rect 81586 82658 81822 82894
rect 81266 82338 81502 82574
rect 81586 82338 81822 82574
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 86378 85222 86614
rect 85306 86378 85542 86614
rect 84986 86058 85222 86294
rect 85306 86058 85542 86294
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 60938 95782 61174
rect 95866 60938 96102 61174
rect 95546 60618 95782 60854
rect 95866 60618 96102 60854
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 64658 99502 64894
rect 99586 64658 99822 64894
rect 99266 64338 99502 64574
rect 99586 64338 99822 64574
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 68378 103222 68614
rect 103306 68378 103542 68614
rect 102986 68058 103222 68294
rect 103306 68058 103542 68294
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 75218 110062 75454
rect 110146 75218 110382 75454
rect 109826 74898 110062 75134
rect 110146 74898 110382 75134
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 78938 113782 79174
rect 113866 78938 114102 79174
rect 113546 78618 113782 78854
rect 113866 78618 114102 78854
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 82658 117502 82894
rect 117586 82658 117822 82894
rect 117266 82338 117502 82574
rect 117586 82338 117822 82574
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 86378 121222 86614
rect 121306 86378 121542 86614
rect 120986 86058 121222 86294
rect 121306 86058 121542 86294
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 60938 131782 61174
rect 131866 60938 132102 61174
rect 131546 60618 131782 60854
rect 131866 60618 132102 60854
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 64658 135502 64894
rect 135586 64658 135822 64894
rect 135266 64338 135502 64574
rect 135586 64338 135822 64574
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 68378 139222 68614
rect 139306 68378 139542 68614
rect 138986 68058 139222 68294
rect 139306 68058 139542 68294
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 75218 146062 75454
rect 146146 75218 146382 75454
rect 145826 74898 146062 75134
rect 146146 74898 146382 75134
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 78938 149782 79174
rect 149866 78938 150102 79174
rect 149546 78618 149782 78854
rect 149866 78618 150102 78854
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 82658 153502 82894
rect 153586 82658 153822 82894
rect 153266 82338 153502 82574
rect 153586 82338 153822 82574
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 86378 157222 86614
rect 157306 86378 157542 86614
rect 156986 86058 157222 86294
rect 157306 86058 157542 86294
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 167546 204938 167782 205174
rect 167866 204938 168102 205174
rect 167546 204618 167782 204854
rect 167866 204618 168102 204854
rect 167546 168938 167782 169174
rect 167866 168938 168102 169174
rect 167546 168618 167782 168854
rect 167866 168618 168102 168854
rect 167546 132938 167782 133174
rect 167866 132938 168102 133174
rect 167546 132618 167782 132854
rect 167866 132618 168102 132854
rect 167546 96938 167782 97174
rect 167866 96938 168102 97174
rect 167546 96618 167782 96854
rect 167866 96618 168102 96854
rect 167546 60938 167782 61174
rect 167866 60938 168102 61174
rect 167546 60618 167782 60854
rect 167866 60618 168102 60854
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 171266 460658 171502 460894
rect 171586 460658 171822 460894
rect 171266 460338 171502 460574
rect 171586 460338 171822 460574
rect 171266 424658 171502 424894
rect 171586 424658 171822 424894
rect 171266 424338 171502 424574
rect 171586 424338 171822 424574
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 174986 464378 175222 464614
rect 175306 464378 175542 464614
rect 174986 464058 175222 464294
rect 175306 464058 175542 464294
rect 174986 428378 175222 428614
rect 175306 428378 175542 428614
rect 174986 428058 175222 428294
rect 175306 428058 175542 428294
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 181826 471218 182062 471454
rect 182146 471218 182382 471454
rect 181826 470898 182062 471134
rect 182146 470898 182382 471134
rect 181826 435218 182062 435454
rect 182146 435218 182382 435454
rect 181826 434898 182062 435134
rect 182146 434898 182382 435134
rect 181826 399218 182062 399454
rect 182146 399218 182382 399454
rect 181826 398898 182062 399134
rect 182146 398898 182382 399134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 185546 474938 185782 475174
rect 185866 474938 186102 475174
rect 185546 474618 185782 474854
rect 185866 474618 186102 474854
rect 185546 438938 185782 439174
rect 185866 438938 186102 439174
rect 185546 438618 185782 438854
rect 185866 438618 186102 438854
rect 185546 402938 185782 403174
rect 185866 402938 186102 403174
rect 185546 402618 185782 402854
rect 185866 402618 186102 402854
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 171266 208658 171502 208894
rect 171586 208658 171822 208894
rect 171266 208338 171502 208574
rect 171586 208338 171822 208574
rect 171266 172658 171502 172894
rect 171586 172658 171822 172894
rect 171266 172338 171502 172574
rect 171586 172338 171822 172574
rect 171266 136658 171502 136894
rect 171586 136658 171822 136894
rect 171266 136338 171502 136574
rect 171586 136338 171822 136574
rect 171266 100658 171502 100894
rect 171586 100658 171822 100894
rect 171266 100338 171502 100574
rect 171586 100338 171822 100574
rect 171266 64658 171502 64894
rect 171586 64658 171822 64894
rect 171266 64338 171502 64574
rect 171586 64338 171822 64574
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 174986 212378 175222 212614
rect 175306 212378 175542 212614
rect 174986 212058 175222 212294
rect 175306 212058 175542 212294
rect 174986 176378 175222 176614
rect 175306 176378 175542 176614
rect 174986 176058 175222 176294
rect 175306 176058 175542 176294
rect 174986 140378 175222 140614
rect 175306 140378 175542 140614
rect 174986 140058 175222 140294
rect 175306 140058 175542 140294
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 189266 478658 189502 478894
rect 189586 478658 189822 478894
rect 189266 478338 189502 478574
rect 189586 478338 189822 478574
rect 189266 442658 189502 442894
rect 189586 442658 189822 442894
rect 189266 442338 189502 442574
rect 189586 442338 189822 442574
rect 189266 406658 189502 406894
rect 189586 406658 189822 406894
rect 189266 406338 189502 406574
rect 189586 406338 189822 406574
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 181826 219218 182062 219454
rect 182146 219218 182382 219454
rect 181826 218898 182062 219134
rect 182146 218898 182382 219134
rect 181826 183218 182062 183454
rect 182146 183218 182382 183454
rect 181826 182898 182062 183134
rect 182146 182898 182382 183134
rect 181826 147218 182062 147454
rect 182146 147218 182382 147454
rect 181826 146898 182062 147134
rect 182146 146898 182382 147134
rect 174986 104378 175222 104614
rect 175306 104378 175542 104614
rect 174986 104058 175222 104294
rect 175306 104058 175542 104294
rect 174986 68378 175222 68614
rect 175306 68378 175542 68614
rect 174986 68058 175222 68294
rect 175306 68058 175542 68294
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 111218 182062 111454
rect 182146 111218 182382 111454
rect 181826 110898 182062 111134
rect 182146 110898 182382 111134
rect 181826 75218 182062 75454
rect 182146 75218 182382 75454
rect 181826 74898 182062 75134
rect 182146 74898 182382 75134
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 185546 222938 185782 223174
rect 185866 222938 186102 223174
rect 185546 222618 185782 222854
rect 185866 222618 186102 222854
rect 185546 186938 185782 187174
rect 185866 186938 186102 187174
rect 185546 186618 185782 186854
rect 185866 186618 186102 186854
rect 185546 150938 185782 151174
rect 185866 150938 186102 151174
rect 185546 150618 185782 150854
rect 185866 150618 186102 150854
rect 185546 114938 185782 115174
rect 185866 114938 186102 115174
rect 185546 114618 185782 114854
rect 185866 114618 186102 114854
rect 185546 78938 185782 79174
rect 185866 78938 186102 79174
rect 185546 78618 185782 78854
rect 185866 78618 186102 78854
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 192986 482378 193222 482614
rect 193306 482378 193542 482614
rect 192986 482058 193222 482294
rect 193306 482058 193542 482294
rect 192986 446378 193222 446614
rect 193306 446378 193542 446614
rect 192986 446058 193222 446294
rect 193306 446058 193542 446294
rect 192986 410378 193222 410614
rect 193306 410378 193542 410614
rect 192986 410058 193222 410294
rect 193306 410058 193542 410294
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 189266 226658 189502 226894
rect 189586 226658 189822 226894
rect 189266 226338 189502 226574
rect 189586 226338 189822 226574
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 189266 190658 189502 190894
rect 189586 190658 189822 190894
rect 189266 190338 189502 190574
rect 189586 190338 189822 190574
rect 189266 154658 189502 154894
rect 189586 154658 189822 154894
rect 189266 154338 189502 154574
rect 189586 154338 189822 154574
rect 189266 118658 189502 118894
rect 189586 118658 189822 118894
rect 189266 118338 189502 118574
rect 189586 118338 189822 118574
rect 189266 82658 189502 82894
rect 189586 82658 189822 82894
rect 189266 82338 189502 82574
rect 189586 82338 189822 82574
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 194378 193222 194614
rect 193306 194378 193542 194614
rect 192986 194058 193222 194294
rect 193306 194058 193542 194294
rect 192986 158378 193222 158614
rect 193306 158378 193542 158614
rect 192986 158058 193222 158294
rect 193306 158058 193542 158294
rect 192986 122378 193222 122614
rect 193306 122378 193542 122614
rect 192986 122058 193222 122294
rect 193306 122058 193542 122294
rect 192986 86378 193222 86614
rect 193306 86378 193542 86614
rect 192986 86058 193222 86294
rect 193306 86058 193542 86294
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 199826 201218 200062 201454
rect 200146 201218 200382 201454
rect 199826 200898 200062 201134
rect 200146 200898 200382 201134
rect 199826 165218 200062 165454
rect 200146 165218 200382 165454
rect 199826 164898 200062 165134
rect 200146 164898 200382 165134
rect 199826 129218 200062 129454
rect 200146 129218 200382 129454
rect 199826 128898 200062 129134
rect 200146 128898 200382 129134
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 204450 255218 204686 255454
rect 204450 254898 204686 255134
rect 203546 204938 203782 205174
rect 203866 204938 204102 205174
rect 203546 204618 203782 204854
rect 203866 204618 204102 204854
rect 203546 168938 203782 169174
rect 203866 168938 204102 169174
rect 203546 168618 203782 168854
rect 203866 168618 204102 168854
rect 203546 132938 203782 133174
rect 203866 132938 204102 133174
rect 203546 132618 203782 132854
rect 203866 132618 204102 132854
rect 203546 96938 203782 97174
rect 203866 96938 204102 97174
rect 203546 96618 203782 96854
rect 203866 96618 204102 96854
rect 199826 93218 200062 93454
rect 200146 93218 200382 93454
rect 199826 92898 200062 93134
rect 200146 92898 200382 93134
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 217826 471218 218062 471454
rect 218146 471218 218382 471454
rect 217826 470898 218062 471134
rect 218146 470898 218382 471134
rect 217826 435218 218062 435454
rect 218146 435218 218382 435454
rect 217826 434898 218062 435134
rect 218146 434898 218382 435134
rect 217826 399218 218062 399454
rect 218146 399218 218382 399454
rect 217826 398898 218062 399134
rect 218146 398898 218382 399134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 221546 474938 221782 475174
rect 221866 474938 222102 475174
rect 221546 474618 221782 474854
rect 221866 474618 222102 474854
rect 221546 438938 221782 439174
rect 221866 438938 222102 439174
rect 221546 438618 221782 438854
rect 221866 438618 222102 438854
rect 221546 402938 221782 403174
rect 221866 402938 222102 403174
rect 221546 402618 221782 402854
rect 221866 402618 222102 402854
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 207266 208658 207502 208894
rect 207586 208658 207822 208894
rect 207266 208338 207502 208574
rect 207586 208338 207822 208574
rect 210986 212378 211222 212614
rect 211306 212378 211542 212614
rect 210986 212058 211222 212294
rect 211306 212058 211542 212294
rect 207266 172658 207502 172894
rect 207586 172658 207822 172894
rect 207266 172338 207502 172574
rect 207586 172338 207822 172574
rect 207266 136658 207502 136894
rect 207586 136658 207822 136894
rect 207266 136338 207502 136574
rect 207586 136338 207822 136574
rect 207266 100658 207502 100894
rect 207586 100658 207822 100894
rect 207266 100338 207502 100574
rect 207586 100338 207822 100574
rect 203546 60938 203782 61174
rect 203866 60938 204102 61174
rect 203546 60618 203782 60854
rect 203866 60618 204102 60854
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 64658 207502 64894
rect 207586 64658 207822 64894
rect 207266 64338 207502 64574
rect 207586 64338 207822 64574
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 176378 211222 176614
rect 211306 176378 211542 176614
rect 210986 176058 211222 176294
rect 211306 176058 211542 176294
rect 210986 140378 211222 140614
rect 211306 140378 211542 140614
rect 210986 140058 211222 140294
rect 211306 140058 211542 140294
rect 210986 104378 211222 104614
rect 211306 104378 211542 104614
rect 210986 104058 211222 104294
rect 211306 104058 211542 104294
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 225266 478658 225502 478894
rect 225586 478658 225822 478894
rect 225266 478338 225502 478574
rect 225586 478338 225822 478574
rect 225266 442658 225502 442894
rect 225586 442658 225822 442894
rect 225266 442338 225502 442574
rect 225586 442338 225822 442574
rect 225266 406658 225502 406894
rect 225586 406658 225822 406894
rect 225266 406338 225502 406574
rect 225586 406338 225822 406574
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 228986 482378 229222 482614
rect 229306 482378 229542 482614
rect 228986 482058 229222 482294
rect 229306 482058 229542 482294
rect 228986 446378 229222 446614
rect 229306 446378 229542 446614
rect 228986 446058 229222 446294
rect 229306 446058 229542 446294
rect 228986 410378 229222 410614
rect 229306 410378 229542 410614
rect 228986 410058 229222 410294
rect 229306 410058 229542 410294
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 219810 273218 220046 273454
rect 219810 272898 220046 273134
rect 217826 219218 218062 219454
rect 218146 219218 218382 219454
rect 217826 218898 218062 219134
rect 218146 218898 218382 219134
rect 221546 222938 221782 223174
rect 221866 222938 222102 223174
rect 221546 222618 221782 222854
rect 221866 222618 222102 222854
rect 217826 183218 218062 183454
rect 218146 183218 218382 183454
rect 217826 182898 218062 183134
rect 218146 182898 218382 183134
rect 221546 186938 221782 187174
rect 221866 186938 222102 187174
rect 221546 186618 221782 186854
rect 221866 186618 222102 186854
rect 225266 226658 225502 226894
rect 225586 226658 225822 226894
rect 225266 226338 225502 226574
rect 225586 226338 225822 226574
rect 225266 190658 225502 190894
rect 225586 190658 225822 190894
rect 225266 190338 225502 190574
rect 225586 190338 225822 190574
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 235826 453218 236062 453454
rect 236146 453218 236382 453454
rect 235826 452898 236062 453134
rect 236146 452898 236382 453134
rect 235826 417218 236062 417454
rect 236146 417218 236382 417454
rect 235826 416898 236062 417134
rect 236146 416898 236382 417134
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 221249 165218 221485 165454
rect 221249 164898 221485 165134
rect 224513 165218 224749 165454
rect 224513 164898 224749 165134
rect 219617 147218 219853 147454
rect 219617 146898 219853 147134
rect 222881 147218 223117 147454
rect 222881 146898 223117 147134
rect 226145 147218 226381 147454
rect 226145 146898 226381 147134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 239546 456938 239782 457174
rect 239866 456938 240102 457174
rect 239546 456618 239782 456854
rect 239866 456618 240102 456854
rect 239546 420938 239782 421174
rect 239866 420938 240102 421174
rect 239546 420618 239782 420854
rect 239866 420618 240102 420854
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235170 255218 235406 255454
rect 235170 254898 235406 255134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 221249 129218 221485 129454
rect 221249 128898 221485 129134
rect 224513 129218 224749 129454
rect 224513 128898 224749 129134
rect 219617 111218 219853 111454
rect 219617 110898 219853 111134
rect 222881 111218 223117 111454
rect 222881 110898 223117 111134
rect 226145 111218 226381 111454
rect 226145 110898 226381 111134
rect 210986 68378 211222 68614
rect 211306 68378 211542 68614
rect 210986 68058 211222 68294
rect 211306 68058 211542 68294
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 75218 218062 75454
rect 218146 75218 218382 75454
rect 217826 74898 218062 75134
rect 218146 74898 218382 75134
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 78938 221782 79174
rect 221866 78938 222102 79174
rect 221546 78618 221782 78854
rect 221866 78618 222102 78854
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 225266 82658 225502 82894
rect 225586 82658 225822 82894
rect 225266 82338 225502 82574
rect 225586 82338 225822 82574
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 243266 460658 243502 460894
rect 243586 460658 243822 460894
rect 243266 460338 243502 460574
rect 243586 460338 243822 460574
rect 243266 424658 243502 424894
rect 243586 424658 243822 424894
rect 243266 424338 243502 424574
rect 243586 424338 243822 424574
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 246986 464378 247222 464614
rect 247306 464378 247542 464614
rect 246986 464058 247222 464294
rect 247306 464058 247542 464294
rect 246986 428378 247222 428614
rect 247306 428378 247542 428614
rect 246986 428058 247222 428294
rect 247306 428058 247542 428294
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 253826 471218 254062 471454
rect 254146 471218 254382 471454
rect 253826 470898 254062 471134
rect 254146 470898 254382 471134
rect 253826 435218 254062 435454
rect 254146 435218 254382 435454
rect 253826 434898 254062 435134
rect 254146 434898 254382 435134
rect 253826 399218 254062 399454
rect 254146 399218 254382 399454
rect 253826 398898 254062 399134
rect 254146 398898 254382 399134
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 257546 474938 257782 475174
rect 257866 474938 258102 475174
rect 257546 474618 257782 474854
rect 257866 474618 258102 474854
rect 257546 438938 257782 439174
rect 257866 438938 258102 439174
rect 257546 438618 257782 438854
rect 257866 438618 258102 438854
rect 257546 402938 257782 403174
rect 257866 402938 258102 403174
rect 257546 402618 257782 402854
rect 257866 402618 258102 402854
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 261266 478658 261502 478894
rect 261586 478658 261822 478894
rect 261266 478338 261502 478574
rect 261586 478338 261822 478574
rect 261266 442658 261502 442894
rect 261586 442658 261822 442894
rect 261266 442338 261502 442574
rect 261586 442338 261822 442574
rect 261266 406658 261502 406894
rect 261586 406658 261822 406894
rect 261266 406338 261502 406574
rect 261586 406338 261822 406574
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 264986 482378 265222 482614
rect 265306 482378 265542 482614
rect 264986 482058 265222 482294
rect 265306 482058 265542 482294
rect 264986 446378 265222 446614
rect 265306 446378 265542 446614
rect 264986 446058 265222 446294
rect 265306 446058 265542 446294
rect 264986 410378 265222 410614
rect 265306 410378 265542 410614
rect 264986 410058 265222 410294
rect 265306 410058 265542 410294
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 271826 453218 272062 453454
rect 272146 453218 272382 453454
rect 271826 452898 272062 453134
rect 272146 452898 272382 453134
rect 271826 417218 272062 417454
rect 272146 417218 272382 417454
rect 271826 416898 272062 417134
rect 272146 416898 272382 417134
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 275546 456938 275782 457174
rect 275866 456938 276102 457174
rect 275546 456618 275782 456854
rect 275866 456618 276102 456854
rect 275546 420938 275782 421174
rect 275866 420938 276102 421174
rect 275546 420618 275782 420854
rect 275866 420618 276102 420854
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 279266 460658 279502 460894
rect 279586 460658 279822 460894
rect 279266 460338 279502 460574
rect 279586 460338 279822 460574
rect 279266 424658 279502 424894
rect 279586 424658 279822 424894
rect 279266 424338 279502 424574
rect 279586 424338 279822 424574
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 282986 464378 283222 464614
rect 283306 464378 283542 464614
rect 282986 464058 283222 464294
rect 283306 464058 283542 464294
rect 282986 428378 283222 428614
rect 283306 428378 283542 428614
rect 282986 428058 283222 428294
rect 283306 428058 283542 428294
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 289826 471218 290062 471454
rect 290146 471218 290382 471454
rect 289826 470898 290062 471134
rect 290146 470898 290382 471134
rect 289826 435218 290062 435454
rect 290146 435218 290382 435454
rect 289826 434898 290062 435134
rect 290146 434898 290382 435134
rect 289826 399218 290062 399454
rect 290146 399218 290382 399454
rect 289826 398898 290062 399134
rect 290146 398898 290382 399134
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 293546 474938 293782 475174
rect 293866 474938 294102 475174
rect 293546 474618 293782 474854
rect 293866 474618 294102 474854
rect 293546 438938 293782 439174
rect 293866 438938 294102 439174
rect 293546 438618 293782 438854
rect 293866 438618 294102 438854
rect 293546 402938 293782 403174
rect 293866 402938 294102 403174
rect 293546 402618 293782 402854
rect 293866 402618 294102 402854
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 272249 165218 272485 165454
rect 272249 164898 272485 165134
rect 275513 165218 275749 165454
rect 275513 164898 275749 165134
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 270617 147218 270853 147454
rect 270617 146898 270853 147134
rect 273881 147218 274117 147454
rect 273881 146898 274117 147134
rect 277145 147218 277381 147454
rect 277145 146898 277381 147134
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 272249 129218 272485 129454
rect 272249 128898 272485 129134
rect 275513 129218 275749 129454
rect 275513 128898 275749 129134
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 270617 111218 270853 111454
rect 270617 110898 270853 111134
rect 273881 111218 274117 111454
rect 273881 110898 274117 111134
rect 277145 111218 277381 111454
rect 277145 110898 277381 111134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 297266 478658 297502 478894
rect 297586 478658 297822 478894
rect 297266 478338 297502 478574
rect 297586 478338 297822 478574
rect 297266 442658 297502 442894
rect 297586 442658 297822 442894
rect 297266 442338 297502 442574
rect 297586 442338 297822 442574
rect 297266 406658 297502 406894
rect 297586 406658 297822 406894
rect 297266 406338 297502 406574
rect 297586 406338 297822 406574
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 300986 482378 301222 482614
rect 301306 482378 301542 482614
rect 300986 482058 301222 482294
rect 301306 482058 301542 482294
rect 300986 446378 301222 446614
rect 301306 446378 301542 446614
rect 300986 446058 301222 446294
rect 301306 446058 301542 446294
rect 300986 410378 301222 410614
rect 301306 410378 301542 410614
rect 300986 410058 301222 410294
rect 301306 410058 301542 410294
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 307826 453218 308062 453454
rect 308146 453218 308382 453454
rect 307826 452898 308062 453134
rect 308146 452898 308382 453134
rect 307826 417218 308062 417454
rect 308146 417218 308382 417454
rect 307826 416898 308062 417134
rect 308146 416898 308382 417134
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 311546 456938 311782 457174
rect 311866 456938 312102 457174
rect 311546 456618 311782 456854
rect 311866 456618 312102 456854
rect 311546 420938 311782 421174
rect 311866 420938 312102 421174
rect 311546 420618 311782 420854
rect 311866 420618 312102 420854
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 315266 460658 315502 460894
rect 315586 460658 315822 460894
rect 315266 460338 315502 460574
rect 315586 460338 315822 460574
rect 315266 424658 315502 424894
rect 315586 424658 315822 424894
rect 315266 424338 315502 424574
rect 315586 424338 315822 424574
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 318986 464378 319222 464614
rect 319306 464378 319542 464614
rect 318986 464058 319222 464294
rect 319306 464058 319542 464294
rect 318986 428378 319222 428614
rect 319306 428378 319542 428614
rect 318986 428058 319222 428294
rect 319306 428058 319542 428294
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 325826 471218 326062 471454
rect 326146 471218 326382 471454
rect 325826 470898 326062 471134
rect 326146 470898 326382 471134
rect 325826 435218 326062 435454
rect 326146 435218 326382 435454
rect 325826 434898 326062 435134
rect 326146 434898 326382 435134
rect 325826 399218 326062 399454
rect 326146 399218 326382 399454
rect 325826 398898 326062 399134
rect 326146 398898 326382 399134
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 329546 474938 329782 475174
rect 329866 474938 330102 475174
rect 329546 474618 329782 474854
rect 329866 474618 330102 474854
rect 329546 438938 329782 439174
rect 329866 438938 330102 439174
rect 329546 438618 329782 438854
rect 329866 438618 330102 438854
rect 329546 402938 329782 403174
rect 329866 402938 330102 403174
rect 329546 402618 329782 402854
rect 329866 402618 330102 402854
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 333266 478658 333502 478894
rect 333586 478658 333822 478894
rect 333266 478338 333502 478574
rect 333586 478338 333822 478574
rect 333266 442658 333502 442894
rect 333586 442658 333822 442894
rect 333266 442338 333502 442574
rect 333586 442338 333822 442574
rect 333266 406658 333502 406894
rect 333586 406658 333822 406894
rect 333266 406338 333502 406574
rect 333586 406338 333822 406574
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 336986 482378 337222 482614
rect 337306 482378 337542 482614
rect 336986 482058 337222 482294
rect 337306 482058 337542 482294
rect 336986 446378 337222 446614
rect 337306 446378 337542 446614
rect 336986 446058 337222 446294
rect 337306 446058 337542 446294
rect 336986 410378 337222 410614
rect 337306 410378 337542 410614
rect 336986 410058 337222 410294
rect 337306 410058 337542 410294
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 343826 453218 344062 453454
rect 344146 453218 344382 453454
rect 343826 452898 344062 453134
rect 344146 452898 344382 453134
rect 343826 417218 344062 417454
rect 344146 417218 344382 417454
rect 343826 416898 344062 417134
rect 344146 416898 344382 417134
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 347546 456938 347782 457174
rect 347866 456938 348102 457174
rect 347546 456618 347782 456854
rect 347866 456618 348102 456854
rect 347546 420938 347782 421174
rect 347866 420938 348102 421174
rect 347546 420618 347782 420854
rect 347866 420618 348102 420854
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 351266 460658 351502 460894
rect 351586 460658 351822 460894
rect 351266 460338 351502 460574
rect 351586 460338 351822 460574
rect 351266 424658 351502 424894
rect 351586 424658 351822 424894
rect 351266 424338 351502 424574
rect 351586 424338 351822 424574
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 354986 464378 355222 464614
rect 355306 464378 355542 464614
rect 354986 464058 355222 464294
rect 355306 464058 355542 464294
rect 354986 428378 355222 428614
rect 355306 428378 355542 428614
rect 354986 428058 355222 428294
rect 355306 428058 355542 428294
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 72721 579454
rect 72957 579218 78651 579454
rect 78887 579218 84582 579454
rect 84818 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 72721 579134
rect 72957 578898 78651 579134
rect 78887 578898 84582 579134
rect 84818 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 75686 561454
rect 75922 561218 81617 561454
rect 81853 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 75686 561134
rect 75922 560898 81617 561134
rect 81853 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 72721 543454
rect 72957 543218 78651 543454
rect 78887 543218 84582 543454
rect 84818 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 72721 543134
rect 72957 542898 78651 543134
rect 78887 542898 84582 543134
rect 84818 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 84986 482614
rect 85222 482378 85306 482614
rect 85542 482378 120986 482614
rect 121222 482378 121306 482614
rect 121542 482378 156986 482614
rect 157222 482378 157306 482614
rect 157542 482378 192986 482614
rect 193222 482378 193306 482614
rect 193542 482378 228986 482614
rect 229222 482378 229306 482614
rect 229542 482378 264986 482614
rect 265222 482378 265306 482614
rect 265542 482378 300986 482614
rect 301222 482378 301306 482614
rect 301542 482378 336986 482614
rect 337222 482378 337306 482614
rect 337542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 84986 482294
rect 85222 482058 85306 482294
rect 85542 482058 120986 482294
rect 121222 482058 121306 482294
rect 121542 482058 156986 482294
rect 157222 482058 157306 482294
rect 157542 482058 192986 482294
rect 193222 482058 193306 482294
rect 193542 482058 228986 482294
rect 229222 482058 229306 482294
rect 229542 482058 264986 482294
rect 265222 482058 265306 482294
rect 265542 482058 300986 482294
rect 301222 482058 301306 482294
rect 301542 482058 336986 482294
rect 337222 482058 337306 482294
rect 337542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 81266 478894
rect 81502 478658 81586 478894
rect 81822 478658 117266 478894
rect 117502 478658 117586 478894
rect 117822 478658 153266 478894
rect 153502 478658 153586 478894
rect 153822 478658 189266 478894
rect 189502 478658 189586 478894
rect 189822 478658 225266 478894
rect 225502 478658 225586 478894
rect 225822 478658 261266 478894
rect 261502 478658 261586 478894
rect 261822 478658 297266 478894
rect 297502 478658 297586 478894
rect 297822 478658 333266 478894
rect 333502 478658 333586 478894
rect 333822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 81266 478574
rect 81502 478338 81586 478574
rect 81822 478338 117266 478574
rect 117502 478338 117586 478574
rect 117822 478338 153266 478574
rect 153502 478338 153586 478574
rect 153822 478338 189266 478574
rect 189502 478338 189586 478574
rect 189822 478338 225266 478574
rect 225502 478338 225586 478574
rect 225822 478338 261266 478574
rect 261502 478338 261586 478574
rect 261822 478338 297266 478574
rect 297502 478338 297586 478574
rect 297822 478338 333266 478574
rect 333502 478338 333586 478574
rect 333822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 77546 475174
rect 77782 474938 77866 475174
rect 78102 474938 113546 475174
rect 113782 474938 113866 475174
rect 114102 474938 149546 475174
rect 149782 474938 149866 475174
rect 150102 474938 185546 475174
rect 185782 474938 185866 475174
rect 186102 474938 221546 475174
rect 221782 474938 221866 475174
rect 222102 474938 257546 475174
rect 257782 474938 257866 475174
rect 258102 474938 293546 475174
rect 293782 474938 293866 475174
rect 294102 474938 329546 475174
rect 329782 474938 329866 475174
rect 330102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 77546 474854
rect 77782 474618 77866 474854
rect 78102 474618 113546 474854
rect 113782 474618 113866 474854
rect 114102 474618 149546 474854
rect 149782 474618 149866 474854
rect 150102 474618 185546 474854
rect 185782 474618 185866 474854
rect 186102 474618 221546 474854
rect 221782 474618 221866 474854
rect 222102 474618 257546 474854
rect 257782 474618 257866 474854
rect 258102 474618 293546 474854
rect 293782 474618 293866 474854
rect 294102 474618 329546 474854
rect 329782 474618 329866 474854
rect 330102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 73826 471454
rect 74062 471218 74146 471454
rect 74382 471218 109826 471454
rect 110062 471218 110146 471454
rect 110382 471218 145826 471454
rect 146062 471218 146146 471454
rect 146382 471218 181826 471454
rect 182062 471218 182146 471454
rect 182382 471218 217826 471454
rect 218062 471218 218146 471454
rect 218382 471218 253826 471454
rect 254062 471218 254146 471454
rect 254382 471218 289826 471454
rect 290062 471218 290146 471454
rect 290382 471218 325826 471454
rect 326062 471218 326146 471454
rect 326382 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 73826 471134
rect 74062 470898 74146 471134
rect 74382 470898 109826 471134
rect 110062 470898 110146 471134
rect 110382 470898 145826 471134
rect 146062 470898 146146 471134
rect 146382 470898 181826 471134
rect 182062 470898 182146 471134
rect 182382 470898 217826 471134
rect 218062 470898 218146 471134
rect 218382 470898 253826 471134
rect 254062 470898 254146 471134
rect 254382 470898 289826 471134
rect 290062 470898 290146 471134
rect 290382 470898 325826 471134
rect 326062 470898 326146 471134
rect 326382 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 66986 464614
rect 67222 464378 67306 464614
rect 67542 464378 102986 464614
rect 103222 464378 103306 464614
rect 103542 464378 138986 464614
rect 139222 464378 139306 464614
rect 139542 464378 174986 464614
rect 175222 464378 175306 464614
rect 175542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 246986 464614
rect 247222 464378 247306 464614
rect 247542 464378 282986 464614
rect 283222 464378 283306 464614
rect 283542 464378 318986 464614
rect 319222 464378 319306 464614
rect 319542 464378 354986 464614
rect 355222 464378 355306 464614
rect 355542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 66986 464294
rect 67222 464058 67306 464294
rect 67542 464058 102986 464294
rect 103222 464058 103306 464294
rect 103542 464058 138986 464294
rect 139222 464058 139306 464294
rect 139542 464058 174986 464294
rect 175222 464058 175306 464294
rect 175542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 246986 464294
rect 247222 464058 247306 464294
rect 247542 464058 282986 464294
rect 283222 464058 283306 464294
rect 283542 464058 318986 464294
rect 319222 464058 319306 464294
rect 319542 464058 354986 464294
rect 355222 464058 355306 464294
rect 355542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 63266 460894
rect 63502 460658 63586 460894
rect 63822 460658 99266 460894
rect 99502 460658 99586 460894
rect 99822 460658 135266 460894
rect 135502 460658 135586 460894
rect 135822 460658 171266 460894
rect 171502 460658 171586 460894
rect 171822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 243266 460894
rect 243502 460658 243586 460894
rect 243822 460658 279266 460894
rect 279502 460658 279586 460894
rect 279822 460658 315266 460894
rect 315502 460658 315586 460894
rect 315822 460658 351266 460894
rect 351502 460658 351586 460894
rect 351822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 63266 460574
rect 63502 460338 63586 460574
rect 63822 460338 99266 460574
rect 99502 460338 99586 460574
rect 99822 460338 135266 460574
rect 135502 460338 135586 460574
rect 135822 460338 171266 460574
rect 171502 460338 171586 460574
rect 171822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 243266 460574
rect 243502 460338 243586 460574
rect 243822 460338 279266 460574
rect 279502 460338 279586 460574
rect 279822 460338 315266 460574
rect 315502 460338 315586 460574
rect 315822 460338 351266 460574
rect 351502 460338 351586 460574
rect 351822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 59546 457174
rect 59782 456938 59866 457174
rect 60102 456938 95546 457174
rect 95782 456938 95866 457174
rect 96102 456938 131546 457174
rect 131782 456938 131866 457174
rect 132102 456938 167546 457174
rect 167782 456938 167866 457174
rect 168102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 239546 457174
rect 239782 456938 239866 457174
rect 240102 456938 275546 457174
rect 275782 456938 275866 457174
rect 276102 456938 311546 457174
rect 311782 456938 311866 457174
rect 312102 456938 347546 457174
rect 347782 456938 347866 457174
rect 348102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 59546 456854
rect 59782 456618 59866 456854
rect 60102 456618 95546 456854
rect 95782 456618 95866 456854
rect 96102 456618 131546 456854
rect 131782 456618 131866 456854
rect 132102 456618 167546 456854
rect 167782 456618 167866 456854
rect 168102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 239546 456854
rect 239782 456618 239866 456854
rect 240102 456618 275546 456854
rect 275782 456618 275866 456854
rect 276102 456618 311546 456854
rect 311782 456618 311866 456854
rect 312102 456618 347546 456854
rect 347782 456618 347866 456854
rect 348102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 91826 453454
rect 92062 453218 92146 453454
rect 92382 453218 127826 453454
rect 128062 453218 128146 453454
rect 128382 453218 163826 453454
rect 164062 453218 164146 453454
rect 164382 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 235826 453454
rect 236062 453218 236146 453454
rect 236382 453218 271826 453454
rect 272062 453218 272146 453454
rect 272382 453218 307826 453454
rect 308062 453218 308146 453454
rect 308382 453218 343826 453454
rect 344062 453218 344146 453454
rect 344382 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 91826 453134
rect 92062 452898 92146 453134
rect 92382 452898 127826 453134
rect 128062 452898 128146 453134
rect 128382 452898 163826 453134
rect 164062 452898 164146 453134
rect 164382 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 235826 453134
rect 236062 452898 236146 453134
rect 236382 452898 271826 453134
rect 272062 452898 272146 453134
rect 272382 452898 307826 453134
rect 308062 452898 308146 453134
rect 308382 452898 343826 453134
rect 344062 452898 344146 453134
rect 344382 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 156986 446614
rect 157222 446378 157306 446614
rect 157542 446378 192986 446614
rect 193222 446378 193306 446614
rect 193542 446378 228986 446614
rect 229222 446378 229306 446614
rect 229542 446378 264986 446614
rect 265222 446378 265306 446614
rect 265542 446378 300986 446614
rect 301222 446378 301306 446614
rect 301542 446378 336986 446614
rect 337222 446378 337306 446614
rect 337542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 156986 446294
rect 157222 446058 157306 446294
rect 157542 446058 192986 446294
rect 193222 446058 193306 446294
rect 193542 446058 228986 446294
rect 229222 446058 229306 446294
rect 229542 446058 264986 446294
rect 265222 446058 265306 446294
rect 265542 446058 300986 446294
rect 301222 446058 301306 446294
rect 301542 446058 336986 446294
rect 337222 446058 337306 446294
rect 337542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 153266 442894
rect 153502 442658 153586 442894
rect 153822 442658 189266 442894
rect 189502 442658 189586 442894
rect 189822 442658 225266 442894
rect 225502 442658 225586 442894
rect 225822 442658 261266 442894
rect 261502 442658 261586 442894
rect 261822 442658 297266 442894
rect 297502 442658 297586 442894
rect 297822 442658 333266 442894
rect 333502 442658 333586 442894
rect 333822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 153266 442574
rect 153502 442338 153586 442574
rect 153822 442338 189266 442574
rect 189502 442338 189586 442574
rect 189822 442338 225266 442574
rect 225502 442338 225586 442574
rect 225822 442338 261266 442574
rect 261502 442338 261586 442574
rect 261822 442338 297266 442574
rect 297502 442338 297586 442574
rect 297822 442338 333266 442574
rect 333502 442338 333586 442574
rect 333822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 149546 439174
rect 149782 438938 149866 439174
rect 150102 438938 185546 439174
rect 185782 438938 185866 439174
rect 186102 438938 221546 439174
rect 221782 438938 221866 439174
rect 222102 438938 257546 439174
rect 257782 438938 257866 439174
rect 258102 438938 293546 439174
rect 293782 438938 293866 439174
rect 294102 438938 329546 439174
rect 329782 438938 329866 439174
rect 330102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 149546 438854
rect 149782 438618 149866 438854
rect 150102 438618 185546 438854
rect 185782 438618 185866 438854
rect 186102 438618 221546 438854
rect 221782 438618 221866 438854
rect 222102 438618 257546 438854
rect 257782 438618 257866 438854
rect 258102 438618 293546 438854
rect 293782 438618 293866 438854
rect 294102 438618 329546 438854
rect 329782 438618 329866 438854
rect 330102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 73020 435454
rect 73256 435218 103740 435454
rect 103976 435218 145826 435454
rect 146062 435218 146146 435454
rect 146382 435218 181826 435454
rect 182062 435218 182146 435454
rect 182382 435218 217826 435454
rect 218062 435218 218146 435454
rect 218382 435218 253826 435454
rect 254062 435218 254146 435454
rect 254382 435218 289826 435454
rect 290062 435218 290146 435454
rect 290382 435218 325826 435454
rect 326062 435218 326146 435454
rect 326382 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 73020 435134
rect 73256 434898 103740 435134
rect 103976 434898 145826 435134
rect 146062 434898 146146 435134
rect 146382 434898 181826 435134
rect 182062 434898 182146 435134
rect 182382 434898 217826 435134
rect 218062 434898 218146 435134
rect 218382 434898 253826 435134
rect 254062 434898 254146 435134
rect 254382 434898 289826 435134
rect 290062 434898 290146 435134
rect 290382 434898 325826 435134
rect 326062 434898 326146 435134
rect 326382 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 138986 428614
rect 139222 428378 139306 428614
rect 139542 428378 174986 428614
rect 175222 428378 175306 428614
rect 175542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 246986 428614
rect 247222 428378 247306 428614
rect 247542 428378 282986 428614
rect 283222 428378 283306 428614
rect 283542 428378 318986 428614
rect 319222 428378 319306 428614
rect 319542 428378 354986 428614
rect 355222 428378 355306 428614
rect 355542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 138986 428294
rect 139222 428058 139306 428294
rect 139542 428058 174986 428294
rect 175222 428058 175306 428294
rect 175542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 246986 428294
rect 247222 428058 247306 428294
rect 247542 428058 282986 428294
rect 283222 428058 283306 428294
rect 283542 428058 318986 428294
rect 319222 428058 319306 428294
rect 319542 428058 354986 428294
rect 355222 428058 355306 428294
rect 355542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 63266 424894
rect 63502 424658 63586 424894
rect 63822 424658 135266 424894
rect 135502 424658 135586 424894
rect 135822 424658 171266 424894
rect 171502 424658 171586 424894
rect 171822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 243266 424894
rect 243502 424658 243586 424894
rect 243822 424658 279266 424894
rect 279502 424658 279586 424894
rect 279822 424658 315266 424894
rect 315502 424658 315586 424894
rect 315822 424658 351266 424894
rect 351502 424658 351586 424894
rect 351822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 63266 424574
rect 63502 424338 63586 424574
rect 63822 424338 135266 424574
rect 135502 424338 135586 424574
rect 135822 424338 171266 424574
rect 171502 424338 171586 424574
rect 171822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 243266 424574
rect 243502 424338 243586 424574
rect 243822 424338 279266 424574
rect 279502 424338 279586 424574
rect 279822 424338 315266 424574
rect 315502 424338 315586 424574
rect 315822 424338 351266 424574
rect 351502 424338 351586 424574
rect 351822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 59546 421174
rect 59782 420938 59866 421174
rect 60102 420938 131546 421174
rect 131782 420938 131866 421174
rect 132102 420938 167546 421174
rect 167782 420938 167866 421174
rect 168102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 239546 421174
rect 239782 420938 239866 421174
rect 240102 420938 275546 421174
rect 275782 420938 275866 421174
rect 276102 420938 311546 421174
rect 311782 420938 311866 421174
rect 312102 420938 347546 421174
rect 347782 420938 347866 421174
rect 348102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 59546 420854
rect 59782 420618 59866 420854
rect 60102 420618 131546 420854
rect 131782 420618 131866 420854
rect 132102 420618 167546 420854
rect 167782 420618 167866 420854
rect 168102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 239546 420854
rect 239782 420618 239866 420854
rect 240102 420618 275546 420854
rect 275782 420618 275866 420854
rect 276102 420618 311546 420854
rect 311782 420618 311866 420854
rect 312102 420618 347546 420854
rect 347782 420618 347866 420854
rect 348102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 88380 417454
rect 88616 417218 119100 417454
rect 119336 417218 127826 417454
rect 128062 417218 128146 417454
rect 128382 417218 163826 417454
rect 164062 417218 164146 417454
rect 164382 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 235826 417454
rect 236062 417218 236146 417454
rect 236382 417218 271826 417454
rect 272062 417218 272146 417454
rect 272382 417218 307826 417454
rect 308062 417218 308146 417454
rect 308382 417218 343826 417454
rect 344062 417218 344146 417454
rect 344382 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 88380 417134
rect 88616 416898 119100 417134
rect 119336 416898 127826 417134
rect 128062 416898 128146 417134
rect 128382 416898 163826 417134
rect 164062 416898 164146 417134
rect 164382 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 235826 417134
rect 236062 416898 236146 417134
rect 236382 416898 271826 417134
rect 272062 416898 272146 417134
rect 272382 416898 307826 417134
rect 308062 416898 308146 417134
rect 308382 416898 343826 417134
rect 344062 416898 344146 417134
rect 344382 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 156986 410614
rect 157222 410378 157306 410614
rect 157542 410378 192986 410614
rect 193222 410378 193306 410614
rect 193542 410378 228986 410614
rect 229222 410378 229306 410614
rect 229542 410378 264986 410614
rect 265222 410378 265306 410614
rect 265542 410378 300986 410614
rect 301222 410378 301306 410614
rect 301542 410378 336986 410614
rect 337222 410378 337306 410614
rect 337542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 156986 410294
rect 157222 410058 157306 410294
rect 157542 410058 192986 410294
rect 193222 410058 193306 410294
rect 193542 410058 228986 410294
rect 229222 410058 229306 410294
rect 229542 410058 264986 410294
rect 265222 410058 265306 410294
rect 265542 410058 300986 410294
rect 301222 410058 301306 410294
rect 301542 410058 336986 410294
rect 337222 410058 337306 410294
rect 337542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 153266 406894
rect 153502 406658 153586 406894
rect 153822 406658 189266 406894
rect 189502 406658 189586 406894
rect 189822 406658 225266 406894
rect 225502 406658 225586 406894
rect 225822 406658 261266 406894
rect 261502 406658 261586 406894
rect 261822 406658 297266 406894
rect 297502 406658 297586 406894
rect 297822 406658 333266 406894
rect 333502 406658 333586 406894
rect 333822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 153266 406574
rect 153502 406338 153586 406574
rect 153822 406338 189266 406574
rect 189502 406338 189586 406574
rect 189822 406338 225266 406574
rect 225502 406338 225586 406574
rect 225822 406338 261266 406574
rect 261502 406338 261586 406574
rect 261822 406338 297266 406574
rect 297502 406338 297586 406574
rect 297822 406338 333266 406574
rect 333502 406338 333586 406574
rect 333822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 149546 403174
rect 149782 402938 149866 403174
rect 150102 402938 185546 403174
rect 185782 402938 185866 403174
rect 186102 402938 221546 403174
rect 221782 402938 221866 403174
rect 222102 402938 257546 403174
rect 257782 402938 257866 403174
rect 258102 402938 293546 403174
rect 293782 402938 293866 403174
rect 294102 402938 329546 403174
rect 329782 402938 329866 403174
rect 330102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 149546 402854
rect 149782 402618 149866 402854
rect 150102 402618 185546 402854
rect 185782 402618 185866 402854
rect 186102 402618 221546 402854
rect 221782 402618 221866 402854
rect 222102 402618 257546 402854
rect 257782 402618 257866 402854
rect 258102 402618 293546 402854
rect 293782 402618 293866 402854
rect 294102 402618 329546 402854
rect 329782 402618 329866 402854
rect 330102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 73020 399454
rect 73256 399218 103740 399454
rect 103976 399218 145826 399454
rect 146062 399218 146146 399454
rect 146382 399218 181826 399454
rect 182062 399218 182146 399454
rect 182382 399218 217826 399454
rect 218062 399218 218146 399454
rect 218382 399218 253826 399454
rect 254062 399218 254146 399454
rect 254382 399218 289826 399454
rect 290062 399218 290146 399454
rect 290382 399218 325826 399454
rect 326062 399218 326146 399454
rect 326382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 73020 399134
rect 73256 398898 103740 399134
rect 103976 398898 145826 399134
rect 146062 398898 146146 399134
rect 146382 398898 181826 399134
rect 182062 398898 182146 399134
rect 182382 398898 217826 399134
rect 218062 398898 218146 399134
rect 218382 398898 253826 399134
rect 254062 398898 254146 399134
rect 254382 398898 289826 399134
rect 290062 398898 290146 399134
rect 290382 398898 325826 399134
rect 326062 398898 326146 399134
rect 326382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 88380 309454
rect 88616 309218 119100 309454
rect 119336 309218 149820 309454
rect 150056 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 88380 309134
rect 88616 308898 119100 309134
rect 119336 308898 149820 309134
rect 150056 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73020 291454
rect 73256 291218 103740 291454
rect 103976 291218 134460 291454
rect 134696 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73020 291134
rect 73256 290898 103740 291134
rect 103976 290898 134460 291134
rect 134696 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 88380 273454
rect 88616 273218 119100 273454
rect 119336 273218 149820 273454
rect 150056 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 219810 273454
rect 220046 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 88380 273134
rect 88616 272898 119100 273134
rect 119336 272898 149820 273134
rect 150056 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 219810 273134
rect 220046 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73020 255454
rect 73256 255218 103740 255454
rect 103976 255218 134460 255454
rect 134696 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 204450 255454
rect 204686 255218 235170 255454
rect 235406 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73020 255134
rect 73256 254898 103740 255134
rect 103976 254898 134460 255134
rect 134696 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 204450 255134
rect 204686 254898 235170 255134
rect 235406 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 81266 226894
rect 81502 226658 81586 226894
rect 81822 226658 117266 226894
rect 117502 226658 117586 226894
rect 117822 226658 153266 226894
rect 153502 226658 153586 226894
rect 153822 226658 189266 226894
rect 189502 226658 189586 226894
rect 189822 226658 225266 226894
rect 225502 226658 225586 226894
rect 225822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 81266 226574
rect 81502 226338 81586 226574
rect 81822 226338 117266 226574
rect 117502 226338 117586 226574
rect 117822 226338 153266 226574
rect 153502 226338 153586 226574
rect 153822 226338 189266 226574
rect 189502 226338 189586 226574
rect 189822 226338 225266 226574
rect 225502 226338 225586 226574
rect 225822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 77546 223174
rect 77782 222938 77866 223174
rect 78102 222938 113546 223174
rect 113782 222938 113866 223174
rect 114102 222938 149546 223174
rect 149782 222938 149866 223174
rect 150102 222938 185546 223174
rect 185782 222938 185866 223174
rect 186102 222938 221546 223174
rect 221782 222938 221866 223174
rect 222102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 77546 222854
rect 77782 222618 77866 222854
rect 78102 222618 113546 222854
rect 113782 222618 113866 222854
rect 114102 222618 149546 222854
rect 149782 222618 149866 222854
rect 150102 222618 185546 222854
rect 185782 222618 185866 222854
rect 186102 222618 221546 222854
rect 221782 222618 221866 222854
rect 222102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 73826 219454
rect 74062 219218 74146 219454
rect 74382 219218 109826 219454
rect 110062 219218 110146 219454
rect 110382 219218 145826 219454
rect 146062 219218 146146 219454
rect 146382 219218 181826 219454
rect 182062 219218 182146 219454
rect 182382 219218 217826 219454
rect 218062 219218 218146 219454
rect 218382 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 73826 219134
rect 74062 218898 74146 219134
rect 74382 218898 109826 219134
rect 110062 218898 110146 219134
rect 110382 218898 145826 219134
rect 146062 218898 146146 219134
rect 146382 218898 181826 219134
rect 182062 218898 182146 219134
rect 182382 218898 217826 219134
rect 218062 218898 218146 219134
rect 218382 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 66986 212614
rect 67222 212378 67306 212614
rect 67542 212378 102986 212614
rect 103222 212378 103306 212614
rect 103542 212378 138986 212614
rect 139222 212378 139306 212614
rect 139542 212378 174986 212614
rect 175222 212378 175306 212614
rect 175542 212378 210986 212614
rect 211222 212378 211306 212614
rect 211542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 66986 212294
rect 67222 212058 67306 212294
rect 67542 212058 102986 212294
rect 103222 212058 103306 212294
rect 103542 212058 138986 212294
rect 139222 212058 139306 212294
rect 139542 212058 174986 212294
rect 175222 212058 175306 212294
rect 175542 212058 210986 212294
rect 211222 212058 211306 212294
rect 211542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 63266 208894
rect 63502 208658 63586 208894
rect 63822 208658 99266 208894
rect 99502 208658 99586 208894
rect 99822 208658 135266 208894
rect 135502 208658 135586 208894
rect 135822 208658 171266 208894
rect 171502 208658 171586 208894
rect 171822 208658 207266 208894
rect 207502 208658 207586 208894
rect 207822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 63266 208574
rect 63502 208338 63586 208574
rect 63822 208338 99266 208574
rect 99502 208338 99586 208574
rect 99822 208338 135266 208574
rect 135502 208338 135586 208574
rect 135822 208338 171266 208574
rect 171502 208338 171586 208574
rect 171822 208338 207266 208574
rect 207502 208338 207586 208574
rect 207822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 59546 205174
rect 59782 204938 59866 205174
rect 60102 204938 95546 205174
rect 95782 204938 95866 205174
rect 96102 204938 131546 205174
rect 131782 204938 131866 205174
rect 132102 204938 167546 205174
rect 167782 204938 167866 205174
rect 168102 204938 203546 205174
rect 203782 204938 203866 205174
rect 204102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 59546 204854
rect 59782 204618 59866 204854
rect 60102 204618 95546 204854
rect 95782 204618 95866 204854
rect 96102 204618 131546 204854
rect 131782 204618 131866 204854
rect 132102 204618 167546 204854
rect 167782 204618 167866 204854
rect 168102 204618 203546 204854
rect 203782 204618 203866 204854
rect 204102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 91826 201454
rect 92062 201218 92146 201454
rect 92382 201218 127826 201454
rect 128062 201218 128146 201454
rect 128382 201218 163826 201454
rect 164062 201218 164146 201454
rect 164382 201218 199826 201454
rect 200062 201218 200146 201454
rect 200382 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 91826 201134
rect 92062 200898 92146 201134
rect 92382 200898 127826 201134
rect 128062 200898 128146 201134
rect 128382 200898 163826 201134
rect 164062 200898 164146 201134
rect 164382 200898 199826 201134
rect 200062 200898 200146 201134
rect 200382 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 84986 194614
rect 85222 194378 85306 194614
rect 85542 194378 120986 194614
rect 121222 194378 121306 194614
rect 121542 194378 156986 194614
rect 157222 194378 157306 194614
rect 157542 194378 192986 194614
rect 193222 194378 193306 194614
rect 193542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 84986 194294
rect 85222 194058 85306 194294
rect 85542 194058 120986 194294
rect 121222 194058 121306 194294
rect 121542 194058 156986 194294
rect 157222 194058 157306 194294
rect 157542 194058 192986 194294
rect 193222 194058 193306 194294
rect 193542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 81266 190894
rect 81502 190658 81586 190894
rect 81822 190658 117266 190894
rect 117502 190658 117586 190894
rect 117822 190658 153266 190894
rect 153502 190658 153586 190894
rect 153822 190658 189266 190894
rect 189502 190658 189586 190894
rect 189822 190658 225266 190894
rect 225502 190658 225586 190894
rect 225822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 81266 190574
rect 81502 190338 81586 190574
rect 81822 190338 117266 190574
rect 117502 190338 117586 190574
rect 117822 190338 153266 190574
rect 153502 190338 153586 190574
rect 153822 190338 189266 190574
rect 189502 190338 189586 190574
rect 189822 190338 225266 190574
rect 225502 190338 225586 190574
rect 225822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 77546 187174
rect 77782 186938 77866 187174
rect 78102 186938 113546 187174
rect 113782 186938 113866 187174
rect 114102 186938 149546 187174
rect 149782 186938 149866 187174
rect 150102 186938 185546 187174
rect 185782 186938 185866 187174
rect 186102 186938 221546 187174
rect 221782 186938 221866 187174
rect 222102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 77546 186854
rect 77782 186618 77866 186854
rect 78102 186618 113546 186854
rect 113782 186618 113866 186854
rect 114102 186618 149546 186854
rect 149782 186618 149866 186854
rect 150102 186618 185546 186854
rect 185782 186618 185866 186854
rect 186102 186618 221546 186854
rect 221782 186618 221866 186854
rect 222102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 73826 183454
rect 74062 183218 74146 183454
rect 74382 183218 109826 183454
rect 110062 183218 110146 183454
rect 110382 183218 145826 183454
rect 146062 183218 146146 183454
rect 146382 183218 181826 183454
rect 182062 183218 182146 183454
rect 182382 183218 217826 183454
rect 218062 183218 218146 183454
rect 218382 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 73826 183134
rect 74062 182898 74146 183134
rect 74382 182898 109826 183134
rect 110062 182898 110146 183134
rect 110382 182898 145826 183134
rect 146062 182898 146146 183134
rect 146382 182898 181826 183134
rect 182062 182898 182146 183134
rect 182382 182898 217826 183134
rect 218062 182898 218146 183134
rect 218382 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 174986 176614
rect 175222 176378 175306 176614
rect 175542 176378 210986 176614
rect 211222 176378 211306 176614
rect 211542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 174986 176294
rect 175222 176058 175306 176294
rect 175542 176058 210986 176294
rect 211222 176058 211306 176294
rect 211542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 63266 172894
rect 63502 172658 63586 172894
rect 63822 172658 171266 172894
rect 171502 172658 171586 172894
rect 171822 172658 207266 172894
rect 207502 172658 207586 172894
rect 207822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 63266 172574
rect 63502 172338 63586 172574
rect 63822 172338 171266 172574
rect 171502 172338 171586 172574
rect 171822 172338 207266 172574
rect 207502 172338 207586 172574
rect 207822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 59546 169174
rect 59782 168938 59866 169174
rect 60102 168938 167546 169174
rect 167782 168938 167866 169174
rect 168102 168938 203546 169174
rect 203782 168938 203866 169174
rect 204102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 59546 168854
rect 59782 168618 59866 168854
rect 60102 168618 167546 168854
rect 167782 168618 167866 168854
rect 168102 168618 203546 168854
rect 203782 168618 203866 168854
rect 204102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 69128 165454
rect 69364 165218 164192 165454
rect 164428 165218 199826 165454
rect 200062 165218 200146 165454
rect 200382 165218 221249 165454
rect 221485 165218 224513 165454
rect 224749 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 272249 165454
rect 272485 165218 275513 165454
rect 275749 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 69128 165134
rect 69364 164898 164192 165134
rect 164428 164898 199826 165134
rect 200062 164898 200146 165134
rect 200382 164898 221249 165134
rect 221485 164898 224513 165134
rect 224749 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 272249 165134
rect 272485 164898 275513 165134
rect 275749 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 192986 158614
rect 193222 158378 193306 158614
rect 193542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 192986 158294
rect 193222 158058 193306 158294
rect 193542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 189266 154894
rect 189502 154658 189586 154894
rect 189822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 189266 154574
rect 189502 154338 189586 154574
rect 189822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 185546 151174
rect 185782 150938 185866 151174
rect 186102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 185546 150854
rect 185782 150618 185866 150854
rect 186102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 69808 147454
rect 70044 147218 163512 147454
rect 163748 147218 181826 147454
rect 182062 147218 182146 147454
rect 182382 147218 219617 147454
rect 219853 147218 222881 147454
rect 223117 147218 226145 147454
rect 226381 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 270617 147454
rect 270853 147218 273881 147454
rect 274117 147218 277145 147454
rect 277381 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 69808 147134
rect 70044 146898 163512 147134
rect 163748 146898 181826 147134
rect 182062 146898 182146 147134
rect 182382 146898 219617 147134
rect 219853 146898 222881 147134
rect 223117 146898 226145 147134
rect 226381 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 270617 147134
rect 270853 146898 273881 147134
rect 274117 146898 277145 147134
rect 277381 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 174986 140614
rect 175222 140378 175306 140614
rect 175542 140378 210986 140614
rect 211222 140378 211306 140614
rect 211542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 174986 140294
rect 175222 140058 175306 140294
rect 175542 140058 210986 140294
rect 211222 140058 211306 140294
rect 211542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 63266 136894
rect 63502 136658 63586 136894
rect 63822 136658 171266 136894
rect 171502 136658 171586 136894
rect 171822 136658 207266 136894
rect 207502 136658 207586 136894
rect 207822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 63266 136574
rect 63502 136338 63586 136574
rect 63822 136338 171266 136574
rect 171502 136338 171586 136574
rect 171822 136338 207266 136574
rect 207502 136338 207586 136574
rect 207822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 59546 133174
rect 59782 132938 59866 133174
rect 60102 132938 167546 133174
rect 167782 132938 167866 133174
rect 168102 132938 203546 133174
rect 203782 132938 203866 133174
rect 204102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 59546 132854
rect 59782 132618 59866 132854
rect 60102 132618 167546 132854
rect 167782 132618 167866 132854
rect 168102 132618 203546 132854
rect 203782 132618 203866 132854
rect 204102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 69128 129454
rect 69364 129218 164192 129454
rect 164428 129218 199826 129454
rect 200062 129218 200146 129454
rect 200382 129218 221249 129454
rect 221485 129218 224513 129454
rect 224749 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 272249 129454
rect 272485 129218 275513 129454
rect 275749 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 69128 129134
rect 69364 128898 164192 129134
rect 164428 128898 199826 129134
rect 200062 128898 200146 129134
rect 200382 128898 221249 129134
rect 221485 128898 224513 129134
rect 224749 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 272249 129134
rect 272485 128898 275513 129134
rect 275749 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 192986 122614
rect 193222 122378 193306 122614
rect 193542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 192986 122294
rect 193222 122058 193306 122294
rect 193542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 189266 118894
rect 189502 118658 189586 118894
rect 189822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 189266 118574
rect 189502 118338 189586 118574
rect 189822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 185546 115174
rect 185782 114938 185866 115174
rect 186102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 185546 114854
rect 185782 114618 185866 114854
rect 186102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 69808 111454
rect 70044 111218 163512 111454
rect 163748 111218 181826 111454
rect 182062 111218 182146 111454
rect 182382 111218 219617 111454
rect 219853 111218 222881 111454
rect 223117 111218 226145 111454
rect 226381 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 270617 111454
rect 270853 111218 273881 111454
rect 274117 111218 277145 111454
rect 277381 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 69808 111134
rect 70044 110898 163512 111134
rect 163748 110898 181826 111134
rect 182062 110898 182146 111134
rect 182382 110898 219617 111134
rect 219853 110898 222881 111134
rect 223117 110898 226145 111134
rect 226381 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 270617 111134
rect 270853 110898 273881 111134
rect 274117 110898 277145 111134
rect 277381 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 174986 104614
rect 175222 104378 175306 104614
rect 175542 104378 210986 104614
rect 211222 104378 211306 104614
rect 211542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 174986 104294
rect 175222 104058 175306 104294
rect 175542 104058 210986 104294
rect 211222 104058 211306 104294
rect 211542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 63266 100894
rect 63502 100658 63586 100894
rect 63822 100658 171266 100894
rect 171502 100658 171586 100894
rect 171822 100658 207266 100894
rect 207502 100658 207586 100894
rect 207822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 63266 100574
rect 63502 100338 63586 100574
rect 63822 100338 171266 100574
rect 171502 100338 171586 100574
rect 171822 100338 207266 100574
rect 207502 100338 207586 100574
rect 207822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 59546 97174
rect 59782 96938 59866 97174
rect 60102 96938 167546 97174
rect 167782 96938 167866 97174
rect 168102 96938 203546 97174
rect 203782 96938 203866 97174
rect 204102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 59546 96854
rect 59782 96618 59866 96854
rect 60102 96618 167546 96854
rect 167782 96618 167866 96854
rect 168102 96618 203546 96854
rect 203782 96618 203866 96854
rect 204102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 199826 93454
rect 200062 93218 200146 93454
rect 200382 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 199826 93134
rect 200062 92898 200146 93134
rect 200382 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 84986 86614
rect 85222 86378 85306 86614
rect 85542 86378 120986 86614
rect 121222 86378 121306 86614
rect 121542 86378 156986 86614
rect 157222 86378 157306 86614
rect 157542 86378 192986 86614
rect 193222 86378 193306 86614
rect 193542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 84986 86294
rect 85222 86058 85306 86294
rect 85542 86058 120986 86294
rect 121222 86058 121306 86294
rect 121542 86058 156986 86294
rect 157222 86058 157306 86294
rect 157542 86058 192986 86294
rect 193222 86058 193306 86294
rect 193542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 81266 82894
rect 81502 82658 81586 82894
rect 81822 82658 117266 82894
rect 117502 82658 117586 82894
rect 117822 82658 153266 82894
rect 153502 82658 153586 82894
rect 153822 82658 189266 82894
rect 189502 82658 189586 82894
rect 189822 82658 225266 82894
rect 225502 82658 225586 82894
rect 225822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 81266 82574
rect 81502 82338 81586 82574
rect 81822 82338 117266 82574
rect 117502 82338 117586 82574
rect 117822 82338 153266 82574
rect 153502 82338 153586 82574
rect 153822 82338 189266 82574
rect 189502 82338 189586 82574
rect 189822 82338 225266 82574
rect 225502 82338 225586 82574
rect 225822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 77546 79174
rect 77782 78938 77866 79174
rect 78102 78938 113546 79174
rect 113782 78938 113866 79174
rect 114102 78938 149546 79174
rect 149782 78938 149866 79174
rect 150102 78938 185546 79174
rect 185782 78938 185866 79174
rect 186102 78938 221546 79174
rect 221782 78938 221866 79174
rect 222102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 77546 78854
rect 77782 78618 77866 78854
rect 78102 78618 113546 78854
rect 113782 78618 113866 78854
rect 114102 78618 149546 78854
rect 149782 78618 149866 78854
rect 150102 78618 185546 78854
rect 185782 78618 185866 78854
rect 186102 78618 221546 78854
rect 221782 78618 221866 78854
rect 222102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 73826 75454
rect 74062 75218 74146 75454
rect 74382 75218 109826 75454
rect 110062 75218 110146 75454
rect 110382 75218 145826 75454
rect 146062 75218 146146 75454
rect 146382 75218 181826 75454
rect 182062 75218 182146 75454
rect 182382 75218 217826 75454
rect 218062 75218 218146 75454
rect 218382 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 73826 75134
rect 74062 74898 74146 75134
rect 74382 74898 109826 75134
rect 110062 74898 110146 75134
rect 110382 74898 145826 75134
rect 146062 74898 146146 75134
rect 146382 74898 181826 75134
rect 182062 74898 182146 75134
rect 182382 74898 217826 75134
rect 218062 74898 218146 75134
rect 218382 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 66986 68614
rect 67222 68378 67306 68614
rect 67542 68378 102986 68614
rect 103222 68378 103306 68614
rect 103542 68378 138986 68614
rect 139222 68378 139306 68614
rect 139542 68378 174986 68614
rect 175222 68378 175306 68614
rect 175542 68378 210986 68614
rect 211222 68378 211306 68614
rect 211542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 66986 68294
rect 67222 68058 67306 68294
rect 67542 68058 102986 68294
rect 103222 68058 103306 68294
rect 103542 68058 138986 68294
rect 139222 68058 139306 68294
rect 139542 68058 174986 68294
rect 175222 68058 175306 68294
rect 175542 68058 210986 68294
rect 211222 68058 211306 68294
rect 211542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 63266 64894
rect 63502 64658 63586 64894
rect 63822 64658 99266 64894
rect 99502 64658 99586 64894
rect 99822 64658 135266 64894
rect 135502 64658 135586 64894
rect 135822 64658 171266 64894
rect 171502 64658 171586 64894
rect 171822 64658 207266 64894
rect 207502 64658 207586 64894
rect 207822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 63266 64574
rect 63502 64338 63586 64574
rect 63822 64338 99266 64574
rect 99502 64338 99586 64574
rect 99822 64338 135266 64574
rect 135502 64338 135586 64574
rect 135822 64338 171266 64574
rect 171502 64338 171586 64574
rect 171822 64338 207266 64574
rect 207502 64338 207586 64574
rect 207822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 59546 61174
rect 59782 60938 59866 61174
rect 60102 60938 95546 61174
rect 95782 60938 95866 61174
rect 96102 60938 131546 61174
rect 131782 60938 131866 61174
rect 132102 60938 167546 61174
rect 167782 60938 167866 61174
rect 168102 60938 203546 61174
rect 203782 60938 203866 61174
rect 204102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 59546 60854
rect 59782 60618 59866 60854
rect 60102 60618 95546 60854
rect 95782 60618 95866 60854
rect 96102 60618 131546 60854
rect 131782 60618 131866 60854
rect 132102 60618 167546 60854
rect 167782 60618 167866 60854
rect 168102 60618 203546 60854
rect 203782 60618 203866 60854
rect 204102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use wrapped_spell  wrapped_spell_1
timestamp 1640170089
transform 1 0 68770 0 1 241592
box 0 0 86000 86000
use wrapped_ppm_decoder  wrapped_ppm_decoder_3
timestamp 1640170089
transform 1 0 68770 0 1 539166
box 0 0 20000 50000
use wrapped_ppm_coder  wrapped_ppm_coder_2
timestamp 1640170089
transform 1 0 68770 0 1 390356
box 0 0 51907 54051
use wrapped_function_generator  wrapped_function_generator_0
timestamp 1640170089
transform 1 0 200200 0 1 240182
box 0 0 44000 44000
use wb_openram_wrapper  wb_openram_wrapper
timestamp 1640170089
transform 1 0 217000 0 1 96000
box 0 144 12000 79688
use wb_bridge_2way  wb_bridge_2way
timestamp 1640170089
transform 1 0 268000 0 1 96000
box 0 0 12000 79688
use sky130_sram_1kbyte_1rw1r_32x256_8  openram_1kB
timestamp 1640170089
transform 1 0 68800 0 1 95100
box 0 0 95956 79500
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 93100 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 94000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 178000 218414 238182 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 176600 74414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 176600 110414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 176600 146414 239592 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 329592 74414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 329592 110414 388356 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 446407 74414 537166 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 591166 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 446407 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 329592 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 286182 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 93100 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 94000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 178000 222134 238182 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 176600 78134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 176600 114134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 176600 150134 239592 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 329592 78134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 329592 114134 388356 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 446407 78134 537166 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 591166 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 446407 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 329592 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 286182 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 93100 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 94000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 178000 225854 238182 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 176600 81854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 176600 117854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 176600 153854 239592 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 329592 81854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 329592 117854 388356 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 446407 81854 537166 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 591166 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 446407 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 329592 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 286182 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 93100 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 94000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 178000 229574 238182 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 176600 85574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 176600 121574 239592 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 329592 85574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 329592 121574 388356 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 446407 85574 537166 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 591166 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 446407 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 176600 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 286182 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 93100 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 94000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 238182 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 238182 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 176600 99854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 176600 135854 239592 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 329592 99854 388356 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 446407 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 329592 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 286182 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 286182 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 178000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 93100 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 238182 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 176600 67574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 176600 103574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 176600 139574 239592 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 329592 67574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 329592 103574 388356 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 446407 67574 537166 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 591166 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 446407 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 329592 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 286182 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 93100 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 94000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 238182 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 238182 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 176600 92414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 176600 128414 239592 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 329592 92414 388356 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 446407 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 329592 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 176600 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 286182 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 286182 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 178000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 93100 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 94000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 238182 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 238182 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 176600 96134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 176600 132134 239592 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 329592 96134 388356 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 446407 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 329592 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 286182 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 286182 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 178000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
