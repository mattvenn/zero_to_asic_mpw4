VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_ppm_decoder
  CLASS BLOCK ;
  FOREIGN wrapped_ppm_decoder ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 250.000 ;
  PIN active
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 241.820 100.000 243.020 ;
    END
  END active
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 97.660 100.000 98.860 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.700 4.000 219.900 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.540 4.000 109.740 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.510 246.000 86.070 250.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.510 246.000 63.070 250.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.140 4.000 123.340 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.740 4.000 34.940 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.910 246.000 12.470 250.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.750 0.000 37.310 4.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.940 4.000 28.140 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 228.220 100.000 229.420 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 56.860 100.000 58.060 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.910 246.000 81.470 250.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.100 4.000 138.300 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.900 4.000 179.100 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 139.820 100.000 141.020 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.140 4.000 21.340 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.700 4.000 185.900 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.310 246.000 30.870 250.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 235.020 100.000 236.220 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 43.260 100.000 44.460 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 111.260 100.000 112.460 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.710 246.000 26.270 250.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.750 0.000 83.310 4.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 153.420 100.000 154.620 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.340 4.000 116.540 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 0.000 32.710 4.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.550 0.000 51.110 4.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 70.460 100.000 71.660 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 150.700 4.000 151.900 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.390 246.000 6.950 250.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 119.420 100.000 120.620 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 160.220 100.000 161.420 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.510 246.000 40.070 250.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 133.020 100.000 134.220 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.110 246.000 44.670 250.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.310 246.000 53.870 250.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.710 246.000 72.270 250.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.310 246.000 99.870 250.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 214.620 100.000 215.820 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.350 0.000 18.910 4.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.300 4.000 233.500 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.750 0.000 60.310 4.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.150 0.000 78.710 4.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 221.420 100.000 222.620 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 29.660 100.000 30.860 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 180.620 100.000 181.820 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.110 246.000 21.670 250.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 94.940 4.000 96.140 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 245.900 4.000 247.100 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.910 246.000 35.470 250.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 9.260 100.000 10.460 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.350 0.000 41.910 4.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 104.460 100.000 105.660 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.790 246.000 2.350 250.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 187.420 100.000 188.620 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.150 0.000 9.710 4.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 36.460 100.000 37.660 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 90.860 100.000 92.060 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.710 246.000 95.270 250.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.300 4.000 165.500 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 16.060 100.000 17.260 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.150 0.000 55.710 4.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.500 4.000 158.700 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 201.020 100.000 202.220 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.140 4.000 89.340 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 63.660 100.000 64.860 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.300 4.000 199.500 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.500 4.000 226.700 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.940 4.000 130.140 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.470 0.000 98.030 4.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.750 0.000 14.310 4.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.340 4.000 82.540 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 50.060 100.000 51.260 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 167.020 100.000 168.220 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 126.220 100.000 127.420 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 2.460 100.000 3.660 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.900 4.000 145.100 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 84.060 100.000 85.260 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 101.740 4.000 102.940 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.540 4.000 7.740 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 194.220 100.000 195.420 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 22.860 100.000 24.060 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 207.820 100.000 209.020 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.950 0.000 69.510 4.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.540 4.000 41.740 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.540 4.000 75.740 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT -0.050 0.000 0.510 4.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.350 0.000 87.910 4.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.900 4.000 213.100 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.510 246.000 17.070 250.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.910 246.000 58.470 250.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.340 4.000 14.540 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.950 0.000 23.510 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.550 0.000 5.110 4.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.310 246.000 76.870 250.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.710 246.000 49.270 250.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.350 0.000 64.910 4.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.110 246.000 90.670 250.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 77.260 100.000 78.460 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.500 4.000 192.700 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 67.740 4.000 68.940 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.550 0.000 28.110 4.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.950 0.000 46.510 4.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.940 4.000 62.140 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 173.820 100.000 175.020 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.550 0.000 74.110 4.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.340 4.000 48.540 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.110 246.000 67.670 250.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.100 4.000 206.300 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.100 4.000 240.300 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.870 0.000 93.430 4.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.140 4.000 55.340 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.100 4.000 172.300 ;
    END
  END io_out[9]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 19.545 10.640 21.145 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.195 10.640 50.795 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 78.850 10.640 80.450 236.880 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 34.370 10.640 35.970 236.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 64.025 10.640 65.625 236.880 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 96.000 146.620 100.000 147.820 ;
    END
  END wb_clk_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 95.075 236.725 ;
      LAYER met1 ;
        RECT 0.070 10.640 99.750 236.880 ;
      LAYER met2 ;
        RECT 0.100 245.720 1.510 246.005 ;
        RECT 2.630 245.720 6.110 246.005 ;
        RECT 7.230 245.720 11.630 246.005 ;
        RECT 12.750 245.720 16.230 246.005 ;
        RECT 17.350 245.720 20.830 246.005 ;
        RECT 21.950 245.720 25.430 246.005 ;
        RECT 26.550 245.720 30.030 246.005 ;
        RECT 31.150 245.720 34.630 246.005 ;
        RECT 35.750 245.720 39.230 246.005 ;
        RECT 40.350 245.720 43.830 246.005 ;
        RECT 44.950 245.720 48.430 246.005 ;
        RECT 49.550 245.720 53.030 246.005 ;
        RECT 54.150 245.720 57.630 246.005 ;
        RECT 58.750 245.720 62.230 246.005 ;
        RECT 63.350 245.720 66.830 246.005 ;
        RECT 67.950 245.720 71.430 246.005 ;
        RECT 72.550 245.720 76.030 246.005 ;
        RECT 77.150 245.720 80.630 246.005 ;
        RECT 81.750 245.720 85.230 246.005 ;
        RECT 86.350 245.720 89.830 246.005 ;
        RECT 90.950 245.720 94.430 246.005 ;
        RECT 95.550 245.720 99.030 246.005 ;
        RECT 0.100 4.280 99.720 245.720 ;
        RECT 0.790 2.875 4.270 4.280 ;
        RECT 5.390 2.875 8.870 4.280 ;
        RECT 9.990 2.875 13.470 4.280 ;
        RECT 14.590 2.875 18.070 4.280 ;
        RECT 19.190 2.875 22.670 4.280 ;
        RECT 23.790 2.875 27.270 4.280 ;
        RECT 28.390 2.875 31.870 4.280 ;
        RECT 32.990 2.875 36.470 4.280 ;
        RECT 37.590 2.875 41.070 4.280 ;
        RECT 42.190 2.875 45.670 4.280 ;
        RECT 46.790 2.875 50.270 4.280 ;
        RECT 51.390 2.875 54.870 4.280 ;
        RECT 55.990 2.875 59.470 4.280 ;
        RECT 60.590 2.875 64.070 4.280 ;
        RECT 65.190 2.875 68.670 4.280 ;
        RECT 69.790 2.875 73.270 4.280 ;
        RECT 74.390 2.875 77.870 4.280 ;
        RECT 78.990 2.875 82.470 4.280 ;
        RECT 83.590 2.875 87.070 4.280 ;
        RECT 88.190 2.875 92.590 4.280 ;
        RECT 93.710 2.875 97.190 4.280 ;
        RECT 98.310 2.875 99.720 4.280 ;
      LAYER met3 ;
        RECT 4.400 245.500 96.000 246.650 ;
        RECT 4.000 243.420 96.000 245.500 ;
        RECT 4.000 241.420 95.600 243.420 ;
        RECT 4.000 240.700 96.000 241.420 ;
        RECT 4.400 238.700 96.000 240.700 ;
        RECT 4.000 236.620 96.000 238.700 ;
        RECT 4.000 234.620 95.600 236.620 ;
        RECT 4.000 233.900 96.000 234.620 ;
        RECT 4.400 231.900 96.000 233.900 ;
        RECT 4.000 229.820 96.000 231.900 ;
        RECT 4.000 227.820 95.600 229.820 ;
        RECT 4.000 227.100 96.000 227.820 ;
        RECT 4.400 225.100 96.000 227.100 ;
        RECT 4.000 223.020 96.000 225.100 ;
        RECT 4.000 221.020 95.600 223.020 ;
        RECT 4.000 220.300 96.000 221.020 ;
        RECT 4.400 218.300 96.000 220.300 ;
        RECT 4.000 216.220 96.000 218.300 ;
        RECT 4.000 214.220 95.600 216.220 ;
        RECT 4.000 213.500 96.000 214.220 ;
        RECT 4.400 211.500 96.000 213.500 ;
        RECT 4.000 209.420 96.000 211.500 ;
        RECT 4.000 207.420 95.600 209.420 ;
        RECT 4.000 206.700 96.000 207.420 ;
        RECT 4.400 204.700 96.000 206.700 ;
        RECT 4.000 202.620 96.000 204.700 ;
        RECT 4.000 200.620 95.600 202.620 ;
        RECT 4.000 199.900 96.000 200.620 ;
        RECT 4.400 197.900 96.000 199.900 ;
        RECT 4.000 195.820 96.000 197.900 ;
        RECT 4.000 193.820 95.600 195.820 ;
        RECT 4.000 193.100 96.000 193.820 ;
        RECT 4.400 191.100 96.000 193.100 ;
        RECT 4.000 189.020 96.000 191.100 ;
        RECT 4.000 187.020 95.600 189.020 ;
        RECT 4.000 186.300 96.000 187.020 ;
        RECT 4.400 184.300 96.000 186.300 ;
        RECT 4.000 182.220 96.000 184.300 ;
        RECT 4.000 180.220 95.600 182.220 ;
        RECT 4.000 179.500 96.000 180.220 ;
        RECT 4.400 177.500 96.000 179.500 ;
        RECT 4.000 175.420 96.000 177.500 ;
        RECT 4.000 173.420 95.600 175.420 ;
        RECT 4.000 172.700 96.000 173.420 ;
        RECT 4.400 170.700 96.000 172.700 ;
        RECT 4.000 168.620 96.000 170.700 ;
        RECT 4.000 166.620 95.600 168.620 ;
        RECT 4.000 165.900 96.000 166.620 ;
        RECT 4.400 163.900 96.000 165.900 ;
        RECT 4.000 161.820 96.000 163.900 ;
        RECT 4.000 159.820 95.600 161.820 ;
        RECT 4.000 159.100 96.000 159.820 ;
        RECT 4.400 157.100 96.000 159.100 ;
        RECT 4.000 155.020 96.000 157.100 ;
        RECT 4.000 153.020 95.600 155.020 ;
        RECT 4.000 152.300 96.000 153.020 ;
        RECT 4.400 150.300 96.000 152.300 ;
        RECT 4.000 148.220 96.000 150.300 ;
        RECT 4.000 146.220 95.600 148.220 ;
        RECT 4.000 145.500 96.000 146.220 ;
        RECT 4.400 143.500 96.000 145.500 ;
        RECT 4.000 141.420 96.000 143.500 ;
        RECT 4.000 139.420 95.600 141.420 ;
        RECT 4.000 138.700 96.000 139.420 ;
        RECT 4.400 136.700 96.000 138.700 ;
        RECT 4.000 134.620 96.000 136.700 ;
        RECT 4.000 132.620 95.600 134.620 ;
        RECT 4.000 130.540 96.000 132.620 ;
        RECT 4.400 128.540 96.000 130.540 ;
        RECT 4.000 127.820 96.000 128.540 ;
        RECT 4.000 125.820 95.600 127.820 ;
        RECT 4.000 123.740 96.000 125.820 ;
        RECT 4.400 121.740 96.000 123.740 ;
        RECT 4.000 121.020 96.000 121.740 ;
        RECT 4.000 119.020 95.600 121.020 ;
        RECT 4.000 116.940 96.000 119.020 ;
        RECT 4.400 114.940 96.000 116.940 ;
        RECT 4.000 112.860 96.000 114.940 ;
        RECT 4.000 110.860 95.600 112.860 ;
        RECT 4.000 110.140 96.000 110.860 ;
        RECT 4.400 108.140 96.000 110.140 ;
        RECT 4.000 106.060 96.000 108.140 ;
        RECT 4.000 104.060 95.600 106.060 ;
        RECT 4.000 103.340 96.000 104.060 ;
        RECT 4.400 101.340 96.000 103.340 ;
        RECT 4.000 99.260 96.000 101.340 ;
        RECT 4.000 97.260 95.600 99.260 ;
        RECT 4.000 96.540 96.000 97.260 ;
        RECT 4.400 94.540 96.000 96.540 ;
        RECT 4.000 92.460 96.000 94.540 ;
        RECT 4.000 90.460 95.600 92.460 ;
        RECT 4.000 89.740 96.000 90.460 ;
        RECT 4.400 87.740 96.000 89.740 ;
        RECT 4.000 85.660 96.000 87.740 ;
        RECT 4.000 83.660 95.600 85.660 ;
        RECT 4.000 82.940 96.000 83.660 ;
        RECT 4.400 80.940 96.000 82.940 ;
        RECT 4.000 78.860 96.000 80.940 ;
        RECT 4.000 76.860 95.600 78.860 ;
        RECT 4.000 76.140 96.000 76.860 ;
        RECT 4.400 74.140 96.000 76.140 ;
        RECT 4.000 72.060 96.000 74.140 ;
        RECT 4.000 70.060 95.600 72.060 ;
        RECT 4.000 69.340 96.000 70.060 ;
        RECT 4.400 67.340 96.000 69.340 ;
        RECT 4.000 65.260 96.000 67.340 ;
        RECT 4.000 63.260 95.600 65.260 ;
        RECT 4.000 62.540 96.000 63.260 ;
        RECT 4.400 60.540 96.000 62.540 ;
        RECT 4.000 58.460 96.000 60.540 ;
        RECT 4.000 56.460 95.600 58.460 ;
        RECT 4.000 55.740 96.000 56.460 ;
        RECT 4.400 53.740 96.000 55.740 ;
        RECT 4.000 51.660 96.000 53.740 ;
        RECT 4.000 49.660 95.600 51.660 ;
        RECT 4.000 48.940 96.000 49.660 ;
        RECT 4.400 46.940 96.000 48.940 ;
        RECT 4.000 44.860 96.000 46.940 ;
        RECT 4.000 42.860 95.600 44.860 ;
        RECT 4.000 42.140 96.000 42.860 ;
        RECT 4.400 40.140 96.000 42.140 ;
        RECT 4.000 38.060 96.000 40.140 ;
        RECT 4.000 36.060 95.600 38.060 ;
        RECT 4.000 35.340 96.000 36.060 ;
        RECT 4.400 33.340 96.000 35.340 ;
        RECT 4.000 31.260 96.000 33.340 ;
        RECT 4.000 29.260 95.600 31.260 ;
        RECT 4.000 28.540 96.000 29.260 ;
        RECT 4.400 26.540 96.000 28.540 ;
        RECT 4.000 24.460 96.000 26.540 ;
        RECT 4.000 22.460 95.600 24.460 ;
        RECT 4.000 21.740 96.000 22.460 ;
        RECT 4.400 19.740 96.000 21.740 ;
        RECT 4.000 17.660 96.000 19.740 ;
        RECT 4.000 15.660 95.600 17.660 ;
        RECT 4.000 14.940 96.000 15.660 ;
        RECT 4.400 12.940 96.000 14.940 ;
        RECT 4.000 10.860 96.000 12.940 ;
        RECT 4.000 8.860 95.600 10.860 ;
        RECT 4.000 8.140 96.000 8.860 ;
        RECT 4.400 6.140 96.000 8.140 ;
        RECT 4.000 4.060 96.000 6.140 ;
        RECT 4.000 2.895 95.600 4.060 ;
  END
END wrapped_ppm_decoder
END LIBRARY

